

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737;

  INV_X2 U373 ( .A(G953), .ZN(n725) );
  XOR2_X1 U374 ( .A(KEYINPUT73), .B(n559), .Z(n351) );
  XNOR2_X2 U375 ( .A(n368), .B(n390), .ZN(n532) );
  XNOR2_X1 U376 ( .A(n514), .B(n505), .ZN(n688) );
  XNOR2_X1 U377 ( .A(n720), .B(n500), .ZN(n514) );
  NOR2_X2 U378 ( .A1(n678), .A2(n530), .ZN(n524) );
  XNOR2_X2 U379 ( .A(n523), .B(n359), .ZN(n678) );
  NOR2_X1 U380 ( .A1(n351), .A2(n372), .ZN(n560) );
  NOR2_X1 U381 ( .A1(G902), .A2(n612), .ZN(n515) );
  XNOR2_X1 U382 ( .A(G113), .B(KEYINPUT3), .ZN(n457) );
  NAND2_X1 U383 ( .A1(n582), .A2(n424), .ZN(n594) );
  XNOR2_X1 U384 ( .A(n366), .B(KEYINPUT40), .ZN(n735) );
  NOR2_X1 U385 ( .A1(n631), .A2(n566), .ZN(n567) );
  XNOR2_X1 U386 ( .A(n411), .B(KEYINPUT116), .ZN(n566) );
  OR2_X1 U387 ( .A1(n565), .A2(n351), .ZN(n411) );
  XNOR2_X1 U388 ( .A(n369), .B(G134), .ZN(n498) );
  XNOR2_X1 U389 ( .A(n506), .B(G469), .ZN(n507) );
  XNOR2_X1 U390 ( .A(n457), .B(G119), .ZN(n383) );
  NAND2_X1 U391 ( .A1(n556), .A2(n406), .ZN(n654) );
  NAND2_X1 U392 ( .A1(n557), .A2(n427), .ZN(n425) );
  NAND2_X1 U393 ( .A1(G214), .A2(n463), .ZN(n652) );
  XNOR2_X1 U394 ( .A(n364), .B(n363), .ZN(n525) );
  XNOR2_X1 U395 ( .A(n490), .B(G475), .ZN(n363) );
  OR2_X1 U396 ( .A1(n692), .A2(G902), .ZN(n364) );
  INV_X1 U397 ( .A(G472), .ZN(n373) );
  NAND2_X1 U398 ( .A1(n604), .A2(n590), .ZN(n380) );
  XNOR2_X1 U399 ( .A(n408), .B(n407), .ZN(n537) );
  XNOR2_X1 U400 ( .A(KEYINPUT112), .B(G478), .ZN(n407) );
  NOR2_X1 U401 ( .A1(n702), .A2(G902), .ZN(n408) );
  INV_X1 U402 ( .A(n639), .ZN(n398) );
  NAND2_X1 U403 ( .A1(G234), .A2(G237), .ZN(n465) );
  INV_X1 U404 ( .A(KEYINPUT70), .ZN(n436) );
  AND2_X1 U405 ( .A1(n542), .A2(KEYINPUT70), .ZN(n528) );
  INV_X1 U406 ( .A(KEYINPUT2), .ZN(n423) );
  AND2_X1 U407 ( .A1(n642), .A2(n581), .ZN(n424) );
  XNOR2_X1 U408 ( .A(n496), .B(KEYINPUT25), .ZN(n430) );
  OR2_X1 U409 ( .A1(n705), .A2(G902), .ZN(n431) );
  XNOR2_X1 U410 ( .A(n561), .B(KEYINPUT1), .ZN(n521) );
  XNOR2_X1 U411 ( .A(n362), .B(G104), .ZN(n483) );
  INV_X1 U412 ( .A(G122), .ZN(n362) );
  XNOR2_X1 U413 ( .A(G110), .B(KEYINPUT16), .ZN(n459) );
  INV_X1 U414 ( .A(KEYINPUT76), .ZN(n458) );
  XNOR2_X1 U415 ( .A(n422), .B(n421), .ZN(n420) );
  XNOR2_X1 U416 ( .A(G119), .B(G137), .ZN(n422) );
  XNOR2_X1 U417 ( .A(G110), .B(G128), .ZN(n421) );
  XNOR2_X1 U418 ( .A(n419), .B(n418), .ZN(n417) );
  XNOR2_X1 U419 ( .A(KEYINPUT23), .B(KEYINPUT100), .ZN(n419) );
  XNOR2_X1 U420 ( .A(KEYINPUT24), .B(KEYINPUT101), .ZN(n418) );
  XNOR2_X1 U421 ( .A(n381), .B(n713), .ZN(n604) );
  XNOR2_X1 U422 ( .A(n455), .B(n382), .ZN(n381) );
  XNOR2_X1 U423 ( .A(n500), .B(n451), .ZN(n455) );
  NAND2_X1 U424 ( .A1(n649), .A2(n406), .ZN(n651) );
  INV_X1 U425 ( .A(n678), .ZN(n370) );
  OR2_X1 U426 ( .A1(n553), .A2(n555), .ZN(n401) );
  XNOR2_X1 U427 ( .A(n464), .B(KEYINPUT19), .ZN(n394) );
  NOR2_X1 U428 ( .A1(n543), .A2(n545), .ZN(n518) );
  XNOR2_X1 U429 ( .A(n391), .B(KEYINPUT22), .ZN(n543) );
  NAND2_X1 U430 ( .A1(n533), .A2(n387), .ZN(n391) );
  NOR2_X1 U431 ( .A1(n650), .A2(n354), .ZN(n387) );
  INV_X1 U432 ( .A(n660), .ZN(n545) );
  XNOR2_X1 U433 ( .A(n514), .B(n412), .ZN(n612) );
  XNOR2_X1 U434 ( .A(n498), .B(n357), .ZN(n477) );
  INV_X1 U435 ( .A(KEYINPUT48), .ZN(n395) );
  INV_X1 U436 ( .A(KEYINPUT82), .ZN(n427) );
  XOR2_X1 U437 ( .A(G113), .B(G143), .Z(n441) );
  XOR2_X1 U438 ( .A(KEYINPUT106), .B(KEYINPUT12), .Z(n480) );
  XNOR2_X1 U439 ( .A(n483), .B(n361), .ZN(n485) );
  INV_X1 U440 ( .A(KEYINPUT107), .ZN(n361) );
  XNOR2_X1 U441 ( .A(n498), .B(n499), .ZN(n720) );
  XNOR2_X1 U442 ( .A(KEYINPUT69), .B(G101), .ZN(n440) );
  XNOR2_X1 U443 ( .A(n450), .B(n449), .ZN(n451) );
  INV_X1 U444 ( .A(G125), .ZN(n449) );
  INV_X1 U445 ( .A(G143), .ZN(n371) );
  XNOR2_X1 U446 ( .A(KEYINPUT97), .B(KEYINPUT96), .ZN(n452) );
  XOR2_X1 U447 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n453) );
  INV_X1 U448 ( .A(n617), .ZN(n433) );
  INV_X1 U449 ( .A(n429), .ZN(n406) );
  INV_X1 U450 ( .A(KEYINPUT78), .ZN(n390) );
  XNOR2_X1 U451 ( .A(G902), .B(KEYINPUT15), .ZN(n590) );
  NOR2_X1 U452 ( .A1(G902), .A2(G237), .ZN(n447) );
  NOR2_X1 U453 ( .A1(n660), .A2(n354), .ZN(n657) );
  NAND2_X1 U454 ( .A1(n525), .A2(n537), .ZN(n650) );
  NOR2_X1 U455 ( .A1(G953), .A2(G237), .ZN(n511) );
  XNOR2_X1 U456 ( .A(G116), .B(KEYINPUT5), .ZN(n509) );
  XOR2_X1 U457 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n510) );
  INV_X1 U458 ( .A(n594), .ZN(n723) );
  XOR2_X1 U459 ( .A(KEYINPUT111), .B(KEYINPUT110), .Z(n472) );
  XNOR2_X1 U460 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n471) );
  XNOR2_X1 U461 ( .A(G122), .B(KEYINPUT109), .ZN(n469) );
  XOR2_X1 U462 ( .A(G140), .B(G104), .Z(n502) );
  XNOR2_X1 U463 ( .A(G107), .B(G110), .ZN(n501) );
  XNOR2_X1 U464 ( .A(n589), .B(n588), .ZN(n646) );
  AND2_X1 U465 ( .A1(n377), .A2(n587), .ZN(n589) );
  XNOR2_X1 U466 ( .A(n409), .B(KEYINPUT41), .ZN(n677) );
  NOR2_X1 U467 ( .A1(n654), .A2(n410), .ZN(n409) );
  INV_X1 U468 ( .A(n652), .ZN(n410) );
  INV_X1 U469 ( .A(KEYINPUT0), .ZN(n378) );
  NAND2_X1 U470 ( .A1(n394), .A2(n355), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n385), .B(KEYINPUT30), .ZN(n553) );
  NAND2_X1 U472 ( .A1(n666), .A2(n652), .ZN(n385) );
  INV_X1 U473 ( .A(n525), .ZN(n538) );
  XNOR2_X1 U474 ( .A(n462), .B(n461), .ZN(n713) );
  XNOR2_X1 U475 ( .A(n383), .B(n470), .ZN(n462) );
  XNOR2_X1 U476 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U477 ( .A(n492), .B(n442), .ZN(n493) );
  XNOR2_X1 U478 ( .A(n420), .B(n417), .ZN(n492) );
  XNOR2_X1 U479 ( .A(n694), .B(n693), .ZN(n695) );
  NAND2_X1 U480 ( .A1(n656), .A2(n370), .ZN(n673) );
  XNOR2_X1 U481 ( .A(n365), .B(KEYINPUT42), .ZN(n737) );
  OR2_X1 U482 ( .A1(n677), .A2(n570), .ZN(n365) );
  NAND2_X1 U483 ( .A1(n376), .A2(n358), .ZN(n580) );
  NAND2_X1 U484 ( .A1(n367), .A2(n376), .ZN(n366) );
  NOR2_X1 U485 ( .A1(n375), .A2(n374), .ZN(n367) );
  NOR2_X1 U486 ( .A1(n585), .A2(n583), .ZN(n568) );
  INV_X1 U487 ( .A(KEYINPUT35), .ZN(n389) );
  XNOR2_X1 U488 ( .A(n439), .B(n438), .ZN(n734) );
  XNOR2_X1 U489 ( .A(n517), .B(KEYINPUT32), .ZN(n438) );
  NOR2_X2 U490 ( .A1(n570), .A2(n379), .ZN(n628) );
  XNOR2_X1 U491 ( .A(n520), .B(KEYINPUT115), .ZN(n733) );
  XNOR2_X1 U492 ( .A(n612), .B(n611), .ZN(n613) );
  INV_X1 U493 ( .A(n702), .ZN(n393) );
  XNOR2_X1 U494 ( .A(n689), .B(n690), .ZN(n388) );
  OR2_X1 U495 ( .A1(n552), .A2(n353), .ZN(n352) );
  OR2_X1 U496 ( .A1(n557), .A2(n427), .ZN(n353) );
  XNOR2_X1 U497 ( .A(n446), .B(KEYINPUT21), .ZN(n354) );
  XOR2_X1 U498 ( .A(n468), .B(KEYINPUT98), .Z(n355) );
  XNOR2_X1 U499 ( .A(n554), .B(KEYINPUT38), .ZN(n429) );
  NAND2_X1 U500 ( .A1(n356), .A2(n352), .ZN(n428) );
  AND2_X1 U501 ( .A1(n426), .A2(n425), .ZN(n356) );
  NAND2_X1 U502 ( .A1(G217), .A2(n491), .ZN(n357) );
  AND2_X1 U503 ( .A1(n384), .A2(n404), .ZN(n358) );
  XOR2_X1 U504 ( .A(n522), .B(KEYINPUT33), .Z(n359) );
  XNOR2_X1 U505 ( .A(KEYINPUT88), .B(KEYINPUT45), .ZN(n360) );
  INV_X1 U506 ( .A(n707), .ZN(n697) );
  NAND2_X1 U507 ( .A1(n735), .A2(n737), .ZN(n564) );
  NAND2_X1 U508 ( .A1(n521), .A2(n657), .ZN(n368) );
  XNOR2_X2 U509 ( .A(n508), .B(n507), .ZN(n561) );
  XNOR2_X1 U510 ( .A(n454), .B(n369), .ZN(n382) );
  XNOR2_X2 U511 ( .A(n456), .B(n371), .ZN(n369) );
  XNOR2_X1 U512 ( .A(n666), .B(KEYINPUT6), .ZN(n565) );
  NAND2_X1 U513 ( .A1(n531), .A2(n372), .ZN(n619) );
  INV_X1 U514 ( .A(n666), .ZN(n372) );
  XNOR2_X2 U515 ( .A(n515), .B(n373), .ZN(n666) );
  INV_X1 U516 ( .A(n384), .ZN(n374) );
  NAND2_X1 U517 ( .A1(n404), .A2(n627), .ZN(n375) );
  NAND2_X1 U518 ( .A1(n400), .A2(n428), .ZN(n376) );
  AND2_X1 U519 ( .A1(n597), .A2(n377), .ZN(n598) );
  NOR2_X1 U520 ( .A1(n377), .A2(KEYINPUT2), .ZN(n643) );
  NAND2_X1 U521 ( .A1(n377), .A2(n725), .ZN(n711) );
  XNOR2_X2 U522 ( .A(n414), .B(n360), .ZN(n377) );
  XNOR2_X1 U523 ( .A(n533), .B(KEYINPUT99), .ZN(n530) );
  XNOR2_X2 U524 ( .A(n413), .B(n378), .ZN(n533) );
  INV_X1 U525 ( .A(n394), .ZN(n379) );
  XNOR2_X2 U526 ( .A(n380), .B(n444), .ZN(n554) );
  XNOR2_X1 U527 ( .A(n513), .B(n383), .ZN(n412) );
  NAND2_X1 U528 ( .A1(n402), .A2(n555), .ZN(n384) );
  NOR2_X1 U529 ( .A1(n434), .A2(n432), .ZN(n416) );
  BUF_X1 U530 ( .A(n666), .Z(n386) );
  NOR2_X1 U531 ( .A1(n429), .A2(n401), .ZN(n400) );
  NOR2_X1 U532 ( .A1(n579), .A2(n398), .ZN(n397) );
  XNOR2_X1 U533 ( .A(n564), .B(n563), .ZN(n399) );
  NOR2_X2 U534 ( .A1(n733), .A2(n734), .ZN(n542) );
  XNOR2_X1 U535 ( .A(n396), .B(n395), .ZN(n582) );
  NAND2_X1 U536 ( .A1(n399), .A2(n397), .ZN(n396) );
  NOR2_X1 U537 ( .A1(n388), .A2(n707), .ZN(G54) );
  NAND2_X1 U538 ( .A1(n541), .A2(n433), .ZN(n432) );
  NAND2_X1 U539 ( .A1(n528), .A2(n732), .ZN(n437) );
  XNOR2_X2 U540 ( .A(n527), .B(n389), .ZN(n732) );
  NOR2_X2 U541 ( .A1(G902), .A2(n688), .ZN(n508) );
  NAND2_X1 U542 ( .A1(n532), .A2(n544), .ZN(n523) );
  NAND2_X1 U543 ( .A1(n554), .A2(n652), .ZN(n464) );
  AND2_X1 U544 ( .A1(n392), .A2(n697), .ZN(G63) );
  XNOR2_X1 U545 ( .A(n701), .B(n393), .ZN(n392) );
  NAND2_X1 U546 ( .A1(n403), .A2(n406), .ZN(n402) );
  INV_X1 U547 ( .A(n553), .ZN(n403) );
  NAND2_X1 U548 ( .A1(n405), .A2(n555), .ZN(n404) );
  INV_X1 U549 ( .A(n428), .ZN(n405) );
  NAND2_X1 U550 ( .A1(n416), .A2(n415), .ZN(n414) );
  XNOR2_X1 U551 ( .A(n437), .B(n529), .ZN(n415) );
  NOR2_X1 U552 ( .A1(n594), .A2(n423), .ZN(n587) );
  NAND2_X1 U553 ( .A1(n552), .A2(n427), .ZN(n426) );
  NOR2_X1 U554 ( .A1(n405), .A2(n553), .ZN(n573) );
  XNOR2_X2 U555 ( .A(n431), .B(n430), .ZN(n660) );
  NOR2_X1 U556 ( .A1(n732), .A2(n435), .ZN(n434) );
  NAND2_X1 U557 ( .A1(n542), .A2(n436), .ZN(n435) );
  NAND2_X1 U558 ( .A1(n518), .A2(n516), .ZN(n439) );
  XNOR2_X2 U559 ( .A(n722), .B(n440), .ZN(n500) );
  XNOR2_X2 U560 ( .A(n448), .B(G146), .ZN(n722) );
  INV_X2 U561 ( .A(KEYINPUT4), .ZN(n448) );
  XNOR2_X1 U562 ( .A(n497), .B(n441), .ZN(n486) );
  AND2_X1 U563 ( .A1(G221), .A2(n491), .ZN(n442) );
  AND2_X1 U564 ( .A1(n511), .A2(G210), .ZN(n443) );
  AND2_X1 U565 ( .A1(n463), .A2(G210), .ZN(n444) );
  INV_X1 U566 ( .A(KEYINPUT80), .ZN(n593) );
  XNOR2_X1 U567 ( .A(n512), .B(n443), .ZN(n513) );
  XNOR2_X1 U568 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U569 ( .A(n460), .B(n483), .ZN(n461) );
  XNOR2_X1 U570 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n478), .B(n477), .ZN(n702) );
  XOR2_X1 U572 ( .A(KEYINPUT95), .B(n607), .Z(n707) );
  NAND2_X1 U573 ( .A1(G234), .A2(n590), .ZN(n445) );
  XNOR2_X1 U574 ( .A(KEYINPUT20), .B(n445), .ZN(n495) );
  NAND2_X1 U575 ( .A1(n495), .A2(G221), .ZN(n446) );
  XNOR2_X1 U576 ( .A(n447), .B(KEYINPUT79), .ZN(n463) );
  NAND2_X1 U577 ( .A1(G224), .A2(n725), .ZN(n450) );
  XNOR2_X1 U578 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X2 U579 ( .A(G128), .B(KEYINPUT84), .ZN(n456) );
  XOR2_X1 U580 ( .A(G116), .B(G107), .Z(n470) );
  XNOR2_X1 U581 ( .A(KEYINPUT14), .B(n465), .ZN(n466) );
  NAND2_X1 U582 ( .A1(G952), .A2(n466), .ZN(n676) );
  NOR2_X1 U583 ( .A1(G953), .A2(n676), .ZN(n550) );
  NAND2_X1 U584 ( .A1(G902), .A2(n466), .ZN(n548) );
  OR2_X1 U585 ( .A1(n725), .A2(G898), .ZN(n715) );
  NOR2_X1 U586 ( .A1(n548), .A2(n715), .ZN(n467) );
  NOR2_X1 U587 ( .A1(n550), .A2(n467), .ZN(n468) );
  XNOR2_X1 U588 ( .A(n470), .B(n469), .ZN(n474) );
  XNOR2_X1 U589 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U590 ( .A(n474), .B(n473), .Z(n478) );
  NAND2_X1 U591 ( .A1(n725), .A2(G234), .ZN(n476) );
  XNOR2_X1 U592 ( .A(KEYINPUT8), .B(KEYINPUT71), .ZN(n475) );
  XNOR2_X1 U593 ( .A(n476), .B(n475), .ZN(n491) );
  XNOR2_X1 U594 ( .A(KEYINPUT11), .B(KEYINPUT105), .ZN(n479) );
  XNOR2_X1 U595 ( .A(n480), .B(n479), .ZN(n482) );
  XNOR2_X1 U596 ( .A(G125), .B(G140), .ZN(n481) );
  XNOR2_X1 U597 ( .A(n481), .B(KEYINPUT10), .ZN(n718) );
  XNOR2_X1 U598 ( .A(G146), .B(n718), .ZN(n494) );
  XNOR2_X1 U599 ( .A(n482), .B(n494), .ZN(n489) );
  NAND2_X1 U600 ( .A1(G214), .A2(n511), .ZN(n484) );
  XNOR2_X1 U601 ( .A(n485), .B(n484), .ZN(n487) );
  XOR2_X1 U602 ( .A(KEYINPUT72), .B(G131), .Z(n497) );
  XNOR2_X1 U603 ( .A(n489), .B(n488), .ZN(n692) );
  XNOR2_X1 U604 ( .A(KEYINPUT108), .B(KEYINPUT13), .ZN(n490) );
  XNOR2_X1 U605 ( .A(n494), .B(n493), .ZN(n705) );
  NAND2_X1 U606 ( .A1(G217), .A2(n495), .ZN(n496) );
  XOR2_X1 U607 ( .A(G137), .B(n497), .Z(n499) );
  XOR2_X1 U608 ( .A(n502), .B(n501), .Z(n504) );
  NAND2_X1 U609 ( .A1(G227), .A2(n725), .ZN(n503) );
  XNOR2_X1 U610 ( .A(KEYINPUT74), .B(KEYINPUT75), .ZN(n506) );
  BUF_X1 U611 ( .A(n521), .Z(n658) );
  XNOR2_X1 U612 ( .A(n510), .B(n509), .ZN(n512) );
  AND2_X1 U613 ( .A1(n565), .A2(n658), .ZN(n516) );
  XOR2_X1 U614 ( .A(KEYINPUT83), .B(KEYINPUT65), .Z(n517) );
  NOR2_X1 U615 ( .A1(n658), .A2(n386), .ZN(n519) );
  NAND2_X1 U616 ( .A1(n518), .A2(n519), .ZN(n520) );
  INV_X1 U617 ( .A(n565), .ZN(n544) );
  INV_X1 U618 ( .A(KEYINPUT93), .ZN(n522) );
  XNOR2_X1 U619 ( .A(n524), .B(KEYINPUT34), .ZN(n526) );
  NOR2_X1 U620 ( .A1(n537), .A2(n525), .ZN(n575) );
  NAND2_X1 U621 ( .A1(n526), .A2(n575), .ZN(n527) );
  INV_X1 U622 ( .A(KEYINPUT44), .ZN(n529) );
  NAND2_X1 U623 ( .A1(n657), .A2(n561), .ZN(n552) );
  NOR2_X1 U624 ( .A1(n530), .A2(n552), .ZN(n531) );
  XOR2_X1 U625 ( .A(KEYINPUT104), .B(KEYINPUT31), .Z(n535) );
  AND2_X1 U626 ( .A1(n386), .A2(n532), .ZN(n668) );
  NAND2_X1 U627 ( .A1(n668), .A2(n533), .ZN(n534) );
  XNOR2_X1 U628 ( .A(n535), .B(n534), .ZN(n635) );
  NAND2_X1 U629 ( .A1(n619), .A2(n635), .ZN(n539) );
  NAND2_X1 U630 ( .A1(n537), .A2(n538), .ZN(n536) );
  XNOR2_X1 U631 ( .A(KEYINPUT113), .B(n536), .ZN(n627) );
  INV_X1 U632 ( .A(n627), .ZN(n631) );
  NOR2_X1 U633 ( .A1(n538), .A2(n537), .ZN(n623) );
  INV_X1 U634 ( .A(n623), .ZN(n634) );
  NAND2_X1 U635 ( .A1(n631), .A2(n634), .ZN(n649) );
  NAND2_X1 U636 ( .A1(n539), .A2(n649), .ZN(n540) );
  XNOR2_X1 U637 ( .A(n540), .B(KEYINPUT114), .ZN(n541) );
  NOR2_X1 U638 ( .A1(n544), .A2(n543), .ZN(n546) );
  NAND2_X1 U639 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U640 ( .A1(n658), .A2(n547), .ZN(n617) );
  XOR2_X1 U641 ( .A(KEYINPUT90), .B(KEYINPUT39), .Z(n555) );
  OR2_X1 U642 ( .A1(n725), .A2(n548), .ZN(n549) );
  NOR2_X1 U643 ( .A1(G900), .A2(n549), .ZN(n551) );
  NOR2_X1 U644 ( .A1(n551), .A2(n550), .ZN(n557) );
  INV_X1 U645 ( .A(n650), .ZN(n556) );
  NOR2_X1 U646 ( .A1(n557), .A2(n354), .ZN(n558) );
  NAND2_X1 U647 ( .A1(n558), .A2(n660), .ZN(n559) );
  XNOR2_X1 U648 ( .A(n560), .B(KEYINPUT28), .ZN(n562) );
  NAND2_X1 U649 ( .A1(n562), .A2(n561), .ZN(n570) );
  XOR2_X1 U650 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n563) );
  INV_X1 U651 ( .A(n554), .ZN(n585) );
  NAND2_X1 U652 ( .A1(n567), .A2(n652), .ZN(n583) );
  XNOR2_X1 U653 ( .A(KEYINPUT36), .B(n568), .ZN(n569) );
  NAND2_X1 U654 ( .A1(n569), .A2(n658), .ZN(n639) );
  NAND2_X1 U655 ( .A1(n628), .A2(n649), .ZN(n572) );
  NOR2_X1 U656 ( .A1(n572), .A2(KEYINPUT77), .ZN(n571) );
  XNOR2_X1 U657 ( .A(n571), .B(KEYINPUT47), .ZN(n578) );
  NAND2_X1 U658 ( .A1(n572), .A2(KEYINPUT77), .ZN(n576) );
  AND2_X1 U659 ( .A1(n554), .A2(n573), .ZN(n574) );
  NAND2_X1 U660 ( .A1(n575), .A2(n574), .ZN(n626) );
  AND2_X1 U661 ( .A1(n576), .A2(n626), .ZN(n577) );
  NAND2_X1 U662 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U663 ( .A1(n580), .A2(n634), .ZN(n640) );
  INV_X1 U664 ( .A(n640), .ZN(n581) );
  OR2_X1 U665 ( .A1(n583), .A2(n658), .ZN(n584) );
  XNOR2_X1 U666 ( .A(n584), .B(KEYINPUT43), .ZN(n586) );
  NAND2_X1 U667 ( .A1(n586), .A2(n585), .ZN(n642) );
  INV_X1 U668 ( .A(KEYINPUT81), .ZN(n588) );
  INV_X1 U669 ( .A(n590), .ZN(n595) );
  XOR2_X1 U670 ( .A(KEYINPUT87), .B(n595), .Z(n591) );
  NAND2_X1 U671 ( .A1(n591), .A2(KEYINPUT2), .ZN(n592) );
  XNOR2_X1 U672 ( .A(n592), .B(KEYINPUT67), .ZN(n599) );
  XNOR2_X1 U673 ( .A(n594), .B(n593), .ZN(n596) );
  AND2_X1 U674 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U675 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X2 U676 ( .A1(n646), .A2(n600), .ZN(n691) );
  NAND2_X1 U677 ( .A1(n691), .A2(G210), .ZN(n606) );
  XOR2_X1 U678 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n602) );
  XNOR2_X1 U679 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n601) );
  XNOR2_X1 U680 ( .A(n602), .B(n601), .ZN(n603) );
  XOR2_X1 U681 ( .A(n604), .B(n603), .Z(n605) );
  XNOR2_X1 U682 ( .A(n606), .B(n605), .ZN(n608) );
  NOR2_X1 U683 ( .A1(G952), .A2(n725), .ZN(n607) );
  NAND2_X1 U684 ( .A1(n608), .A2(n697), .ZN(n610) );
  XNOR2_X1 U685 ( .A(KEYINPUT89), .B(KEYINPUT56), .ZN(n609) );
  XNOR2_X1 U686 ( .A(n610), .B(n609), .ZN(G51) );
  NAND2_X1 U687 ( .A1(n691), .A2(G472), .ZN(n614) );
  XOR2_X1 U688 ( .A(KEYINPUT62), .B(KEYINPUT94), .Z(n611) );
  XNOR2_X1 U689 ( .A(n614), .B(n613), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n615), .A2(n697), .ZN(n616) );
  XNOR2_X1 U691 ( .A(n616), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U692 ( .A(G101), .B(n617), .Z(G3) );
  NOR2_X1 U693 ( .A1(n631), .A2(n619), .ZN(n618) );
  XOR2_X1 U694 ( .A(G104), .B(n618), .Z(G6) );
  NOR2_X1 U695 ( .A1(n634), .A2(n619), .ZN(n621) );
  XNOR2_X1 U696 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n620) );
  XNOR2_X1 U697 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U698 ( .A(G107), .B(n622), .ZN(G9) );
  XOR2_X1 U699 ( .A(G128), .B(KEYINPUT29), .Z(n625) );
  NAND2_X1 U700 ( .A1(n628), .A2(n623), .ZN(n624) );
  XNOR2_X1 U701 ( .A(n625), .B(n624), .ZN(G30) );
  XNOR2_X1 U702 ( .A(G143), .B(n626), .ZN(G45) );
  XOR2_X1 U703 ( .A(G146), .B(KEYINPUT117), .Z(n630) );
  NAND2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U705 ( .A(n630), .B(n629), .ZN(G48) );
  NOR2_X1 U706 ( .A1(n635), .A2(n631), .ZN(n632) );
  XOR2_X1 U707 ( .A(KEYINPUT118), .B(n632), .Z(n633) );
  XNOR2_X1 U708 ( .A(G113), .B(n633), .ZN(G15) );
  NOR2_X1 U709 ( .A1(n635), .A2(n634), .ZN(n637) );
  XNOR2_X1 U710 ( .A(G116), .B(KEYINPUT119), .ZN(n636) );
  XNOR2_X1 U711 ( .A(n637), .B(n636), .ZN(G18) );
  XOR2_X1 U712 ( .A(G125), .B(KEYINPUT37), .Z(n638) );
  XNOR2_X1 U713 ( .A(n639), .B(n638), .ZN(G27) );
  XOR2_X1 U714 ( .A(G134), .B(n640), .Z(n641) );
  XNOR2_X1 U715 ( .A(KEYINPUT120), .B(n641), .ZN(G36) );
  XNOR2_X1 U716 ( .A(G140), .B(n642), .ZN(G42) );
  XNOR2_X1 U717 ( .A(n643), .B(KEYINPUT85), .ZN(n648) );
  NOR2_X1 U718 ( .A1(n723), .A2(KEYINPUT2), .ZN(n644) );
  XNOR2_X1 U719 ( .A(KEYINPUT86), .B(n644), .ZN(n645) );
  NOR2_X1 U720 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U721 ( .A1(n648), .A2(n647), .ZN(n682) );
  NAND2_X1 U722 ( .A1(n651), .A2(n650), .ZN(n653) );
  NAND2_X1 U723 ( .A1(n653), .A2(n652), .ZN(n655) );
  NAND2_X1 U724 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U725 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U726 ( .A(KEYINPUT50), .B(n659), .Z(n664) );
  NAND2_X1 U727 ( .A1(n354), .A2(n660), .ZN(n661) );
  XNOR2_X1 U728 ( .A(n661), .B(KEYINPUT49), .ZN(n662) );
  XNOR2_X1 U729 ( .A(KEYINPUT121), .B(n662), .ZN(n663) );
  NAND2_X1 U730 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U731 ( .A1(n386), .A2(n665), .ZN(n667) );
  NOR2_X1 U732 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U733 ( .A(KEYINPUT51), .B(n669), .ZN(n671) );
  INV_X1 U734 ( .A(n677), .ZN(n670) );
  NAND2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U736 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U737 ( .A(KEYINPUT52), .B(n674), .Z(n675) );
  NOR2_X1 U738 ( .A1(n676), .A2(n675), .ZN(n680) );
  NOR2_X1 U739 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U740 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U741 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U742 ( .A1(n683), .A2(G953), .ZN(n684) );
  XNOR2_X1 U743 ( .A(n684), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U744 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n686) );
  XNOR2_X1 U745 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n685) );
  XNOR2_X1 U746 ( .A(n686), .B(n685), .ZN(n687) );
  XOR2_X1 U747 ( .A(n688), .B(n687), .Z(n690) );
  BUF_X2 U748 ( .A(n691), .Z(n703) );
  NAND2_X1 U749 ( .A1(n703), .A2(G469), .ZN(n689) );
  NAND2_X1 U750 ( .A1(n691), .A2(G475), .ZN(n696) );
  XNOR2_X1 U751 ( .A(KEYINPUT59), .B(KEYINPUT124), .ZN(n694) );
  XNOR2_X1 U752 ( .A(n692), .B(KEYINPUT66), .ZN(n693) );
  XNOR2_X1 U753 ( .A(n696), .B(n695), .ZN(n698) );
  NAND2_X1 U754 ( .A1(n698), .A2(n697), .ZN(n700) );
  XOR2_X1 U755 ( .A(KEYINPUT68), .B(KEYINPUT60), .Z(n699) );
  XNOR2_X1 U756 ( .A(n700), .B(n699), .ZN(G60) );
  NAND2_X1 U757 ( .A1(G478), .A2(n703), .ZN(n701) );
  NAND2_X1 U758 ( .A1(G217), .A2(n703), .ZN(n704) );
  XNOR2_X1 U759 ( .A(n704), .B(n705), .ZN(n706) );
  NOR2_X1 U760 ( .A1(n707), .A2(n706), .ZN(G66) );
  XOR2_X1 U761 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n709) );
  NAND2_X1 U762 ( .A1(G224), .A2(G953), .ZN(n708) );
  XNOR2_X1 U763 ( .A(n709), .B(n708), .ZN(n710) );
  NAND2_X1 U764 ( .A1(n710), .A2(G898), .ZN(n712) );
  NAND2_X1 U765 ( .A1(n712), .A2(n711), .ZN(n717) );
  XNOR2_X1 U766 ( .A(n713), .B(G101), .ZN(n714) );
  NAND2_X1 U767 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U768 ( .A(n717), .B(n716), .Z(G69) );
  XOR2_X1 U769 ( .A(n718), .B(KEYINPUT126), .Z(n719) );
  XNOR2_X1 U770 ( .A(n720), .B(n719), .ZN(n721) );
  XOR2_X1 U771 ( .A(n722), .B(n721), .Z(n727) );
  INV_X1 U772 ( .A(n727), .ZN(n724) );
  XOR2_X1 U773 ( .A(n724), .B(n723), .Z(n726) );
  NAND2_X1 U774 ( .A1(n726), .A2(n725), .ZN(n731) );
  XOR2_X1 U775 ( .A(G227), .B(n727), .Z(n728) );
  NAND2_X1 U776 ( .A1(n728), .A2(G900), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n729), .A2(G953), .ZN(n730) );
  NAND2_X1 U778 ( .A1(n731), .A2(n730), .ZN(G72) );
  XNOR2_X1 U779 ( .A(G122), .B(n732), .ZN(G24) );
  XOR2_X1 U780 ( .A(n733), .B(G110), .Z(G12) );
  XOR2_X1 U781 ( .A(n734), .B(G119), .Z(G21) );
  XOR2_X1 U782 ( .A(n735), .B(G131), .Z(n736) );
  XNOR2_X1 U783 ( .A(KEYINPUT127), .B(n736), .ZN(G33) );
  XNOR2_X1 U784 ( .A(G137), .B(n737), .ZN(G39) );
endmodule

