//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  NAND3_X1  g001(.A1(new_n202), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n203));
  AND2_X1   g002(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(new_n206), .B2(G36gat), .ZN(new_n207));
  OR2_X1    g006(.A1(new_n207), .A2(KEYINPUT15), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(KEYINPUT15), .ZN(new_n209));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(new_n209), .B2(new_n210), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(KEYINPUT17), .ZN(new_n213));
  XNOR2_X1  g012(.A(G15gat), .B(G22gat), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n214), .A2(G1gat), .ZN(new_n215));
  AOI21_X1  g014(.A(G8gat), .B1(new_n215), .B2(KEYINPUT96), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT16), .ZN(new_n217));
  NOR3_X1   g016(.A1(new_n217), .A2(KEYINPUT95), .A3(G1gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT95), .B1(new_n217), .B2(G1gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n215), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n216), .B(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT97), .ZN(new_n223));
  INV_X1    g022(.A(new_n222), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n213), .A2(new_n223), .B1(new_n224), .B2(new_n212), .ZN(new_n225));
  NAND2_X1  g024(.A1(G229gat), .A2(G233gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(KEYINPUT18), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT98), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(new_n212), .B(new_n222), .Z(new_n230));
  XOR2_X1   g029(.A(new_n226), .B(KEYINPUT13), .Z(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n227), .A2(new_n228), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n229), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n225), .A2(new_n226), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT18), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n238), .A2(KEYINPUT99), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(KEYINPUT99), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G113gat), .B(G141gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(G197gat), .ZN(new_n243));
  XOR2_X1   g042(.A(KEYINPUT11), .B(G169gat), .Z(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n245), .B(KEYINPUT12), .Z(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n235), .A2(new_n241), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n247), .B1(new_n235), .B2(new_n238), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT31), .B(G50gat), .ZN(new_n252));
  XOR2_X1   g051(.A(new_n252), .B(G106gat), .Z(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G141gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G148gat), .ZN(new_n256));
  INV_X1    g055(.A(G148gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G141gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n256), .A2(new_n258), .A3(KEYINPUT82), .ZN(new_n259));
  XNOR2_X1  g058(.A(G155gat), .B(G162gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT82), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n261), .A2(new_n255), .A3(G148gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT2), .ZN(new_n264));
  INV_X1    g063(.A(G162gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT83), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT83), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G162gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n264), .B1(new_n269), .B2(G155gat), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT2), .B1(new_n256), .B2(new_n258), .ZN(new_n271));
  OR3_X1    g070(.A1(KEYINPUT81), .A2(G155gat), .A3(G162gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT81), .B1(G155gat), .B2(G162gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  OAI22_X1  g074(.A1(new_n263), .A2(new_n270), .B1(new_n271), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT22), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n277), .A2(KEYINPUT77), .B1(G211gat), .B2(G218gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT77), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT22), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G197gat), .B(G204gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G211gat), .B(G218gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n281), .A2(new_n284), .A3(new_n282), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT29), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n276), .B1(new_n288), .B2(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g088(.A1(G228gat), .A2(G233gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n286), .A2(new_n287), .ZN(new_n293));
  XNOR2_X1  g092(.A(KEYINPUT83), .B(G162gat), .ZN(new_n294));
  INV_X1    g093(.A(G155gat), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT2), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n296), .A2(new_n259), .A3(new_n260), .A4(new_n262), .ZN(new_n297));
  INV_X1    g096(.A(new_n271), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n298), .A2(new_n273), .A3(new_n272), .A4(new_n274), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT3), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT29), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n293), .B1(new_n303), .B2(KEYINPUT88), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT88), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n301), .A2(new_n305), .A3(new_n302), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n292), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n287), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n284), .B1(new_n281), .B2(new_n282), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT87), .ZN(new_n310));
  NOR3_X1   g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n302), .B1(new_n286), .B2(KEYINPUT87), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n300), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n276), .A2(KEYINPUT84), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT84), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n299), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n293), .B1(new_n301), .B2(new_n302), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n291), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(G22gat), .B1(new_n307), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G78gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n303), .A2(KEYINPUT88), .ZN(new_n324));
  INV_X1    g123(.A(new_n293), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(new_n325), .A3(new_n306), .ZN(new_n326));
  INV_X1    g125(.A(new_n292), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G22gat), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT29), .B1(new_n309), .B2(new_n310), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(new_n293), .B2(new_n310), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n331), .A2(new_n300), .B1(new_n314), .B2(new_n316), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n290), .B1(new_n332), .B2(new_n319), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n328), .A2(new_n329), .A3(new_n333), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n322), .A2(new_n323), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n323), .B1(new_n322), .B2(new_n334), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n254), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NOR3_X1   g136(.A1(new_n307), .A2(new_n321), .A3(G22gat), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n329), .B1(new_n328), .B2(new_n333), .ZN(new_n339));
  OAI21_X1  g138(.A(G78gat), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n322), .A2(new_n334), .A3(new_n323), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n341), .A3(new_n253), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT25), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT23), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g146(.A(KEYINPUT64), .B(KEYINPUT23), .C1(G169gat), .C2(G176gat), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT24), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(G183gat), .A3(G190gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(G183gat), .A2(G190gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT24), .ZN(new_n354));
  NOR2_X1   g153(.A1(G183gat), .A2(G190gat), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n350), .B(new_n352), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n344), .B1(new_n349), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n347), .A2(new_n348), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n352), .A2(new_n350), .ZN(new_n359));
  INV_X1    g158(.A(new_n355), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(KEYINPUT24), .A3(new_n353), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n358), .A2(new_n359), .A3(new_n361), .A4(KEYINPUT25), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  XOR2_X1   g162(.A(G127gat), .B(G134gat), .Z(new_n364));
  XNOR2_X1  g163(.A(G113gat), .B(G120gat), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n364), .B(KEYINPUT67), .C1(KEYINPUT1), .C2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT67), .ZN(new_n367));
  INV_X1    g166(.A(G120gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G113gat), .ZN(new_n369));
  INV_X1    g168(.A(G113gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G120gat), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT1), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G127gat), .B(G134gat), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n367), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n364), .A2(KEYINPUT1), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT68), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n370), .A2(KEYINPUT68), .A3(G120gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n369), .A3(new_n378), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n366), .A2(new_n374), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(G183gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT27), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT27), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(G183gat), .ZN(new_n384));
  INV_X1    g183(.A(G190gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT65), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT66), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT28), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT65), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n382), .A2(new_n384), .A3(new_n390), .A4(new_n385), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n387), .A2(new_n388), .A3(new_n389), .A4(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G169gat), .ZN(new_n393));
  INV_X1    g192(.A(G176gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT26), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n353), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT26), .B1(new_n393), .B2(new_n394), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n397), .B1(new_n350), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n392), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT66), .B1(new_n386), .B2(new_n389), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT28), .B1(new_n386), .B2(KEYINPUT65), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n401), .B1(new_n391), .B2(new_n402), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n363), .B(new_n380), .C1(new_n400), .C2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT69), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n387), .A2(new_n389), .A3(new_n391), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n392), .B(new_n399), .C1(new_n407), .C2(new_n401), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n408), .A2(KEYINPUT69), .A3(new_n380), .A4(new_n363), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n363), .B1(new_n400), .B2(new_n403), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n366), .A2(new_n374), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n375), .A2(new_n379), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n406), .A2(new_n409), .A3(new_n414), .ZN(new_n415));
  AND2_X1   g214(.A1(G227gat), .A2(G233gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT32), .ZN(new_n418));
  XNOR2_X1  g217(.A(G15gat), .B(G43gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(G71gat), .B(G99gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT33), .B1(new_n422), .B2(KEYINPUT72), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n423), .B1(KEYINPUT72), .B2(new_n422), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT33), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n421), .B1(new_n417), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT70), .B1(new_n417), .B2(KEYINPUT32), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT70), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT32), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n429), .B(new_n430), .C1(new_n415), .C2(new_n416), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n427), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT71), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT71), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n434), .B(new_n427), .C1(new_n428), .C2(new_n431), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n425), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT74), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n437), .B1(new_n415), .B2(new_n416), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT34), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n343), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n439), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT73), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n441), .B1(new_n436), .B2(new_n442), .ZN(new_n443));
  AOI211_X1 g242(.A(KEYINPUT73), .B(new_n425), .C1(new_n433), .C2(new_n435), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n440), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT94), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT4), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n314), .A2(new_n316), .A3(new_n448), .A4(new_n380), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n411), .A2(new_n297), .A3(new_n299), .A4(new_n412), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT4), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT5), .ZN(new_n453));
  NAND2_X1  g252(.A1(G225gat), .A2(G233gat), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n276), .A2(KEYINPUT3), .B1(new_n411), .B2(new_n412), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n455), .B1(new_n456), .B2(new_n301), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n452), .A2(new_n453), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT86), .ZN(new_n459));
  INV_X1    g258(.A(new_n450), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n411), .A2(new_n412), .B1(new_n297), .B2(new_n299), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n459), .B(KEYINPUT5), .C1(new_n462), .C2(new_n454), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n413), .A2(new_n276), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n454), .B1(new_n464), .B2(new_n450), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT86), .B1(new_n465), .B2(new_n453), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT4), .B1(new_n317), .B2(new_n413), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n460), .A2(KEYINPUT85), .A3(new_n448), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT85), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n470), .B1(new_n450), .B2(KEYINPUT4), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n468), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n457), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n458), .B1(new_n467), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(G1gat), .B(G29gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(KEYINPUT0), .ZN(new_n476));
  XNOR2_X1  g275(.A(G57gat), .B(G85gat), .ZN(new_n477));
  XOR2_X1   g276(.A(new_n476), .B(new_n477), .Z(new_n478));
  AOI21_X1  g277(.A(KEYINPUT6), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n479), .B1(new_n478), .B2(new_n474), .ZN(new_n480));
  INV_X1    g279(.A(new_n478), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n463), .A2(new_n466), .B1(new_n472), .B2(new_n457), .ZN(new_n482));
  OAI211_X1 g281(.A(KEYINPUT6), .B(new_n481), .C1(new_n482), .C2(new_n458), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(G226gat), .A2(G233gat), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n487), .B1(new_n410), .B2(new_n302), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n486), .B1(new_n408), .B2(new_n363), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n325), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n410), .A2(new_n487), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT29), .B1(new_n408), .B2(new_n363), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n491), .B(new_n293), .C1(new_n492), .C2(new_n487), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT78), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n490), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  OAI211_X1 g294(.A(KEYINPUT78), .B(new_n325), .C1(new_n488), .C2(new_n489), .ZN(new_n496));
  XNOR2_X1  g295(.A(G8gat), .B(G36gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(G64gat), .B(G92gat), .ZN(new_n498));
  XOR2_X1   g297(.A(new_n497), .B(new_n498), .Z(new_n499));
  XOR2_X1   g298(.A(new_n499), .B(KEYINPUT79), .Z(new_n500));
  NAND3_X1  g299(.A1(new_n495), .A2(new_n496), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT80), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n501), .A2(new_n502), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT30), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n495), .A2(new_n496), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n505), .B1(new_n506), .B2(new_n499), .ZN(new_n507));
  INV_X1    g306(.A(new_n499), .ZN(new_n508));
  AOI211_X1 g307(.A(KEYINPUT30), .B(new_n508), .C1(new_n495), .C2(new_n496), .ZN(new_n509));
  OAI22_X1  g308(.A1(new_n503), .A2(new_n504), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n485), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n440), .B(KEYINPUT94), .C1(new_n443), .C2(new_n444), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n447), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT35), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT76), .B1(new_n436), .B2(new_n439), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n433), .A2(new_n435), .ZN(new_n516));
  INV_X1    g315(.A(new_n425), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT76), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n519), .A3(new_n441), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT75), .ZN(new_n521));
  AND4_X1   g320(.A1(new_n521), .A2(new_n516), .A3(new_n517), .A4(new_n439), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n521), .B1(new_n436), .B2(new_n439), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n515), .B(new_n520), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n343), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n481), .B1(new_n474), .B2(KEYINPUT91), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT91), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n482), .A2(new_n527), .A3(new_n458), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n479), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n483), .ZN(new_n530));
  INV_X1    g329(.A(new_n510), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT35), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n525), .A2(new_n530), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n524), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n514), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT36), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n524), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n444), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n518), .A2(KEYINPUT73), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(new_n540), .A3(new_n441), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n537), .B1(new_n436), .B2(new_n439), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT37), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n506), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n495), .A2(KEYINPUT37), .A3(new_n496), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(new_n508), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT38), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n545), .B1(new_n490), .B2(new_n493), .ZN(new_n550));
  INV_X1    g349(.A(new_n500), .ZN(new_n551));
  NOR3_X1   g350(.A1(new_n550), .A2(KEYINPUT38), .A3(new_n551), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n546), .A2(new_n552), .B1(new_n506), .B2(new_n499), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n529), .A2(new_n549), .A3(new_n483), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n525), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n526), .A2(new_n528), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n456), .A2(new_n301), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n452), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n559), .A2(KEYINPUT89), .A3(new_n455), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT89), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n449), .A2(new_n451), .B1(new_n301), .B2(new_n456), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n561), .B1(new_n562), .B2(new_n454), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT39), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n565), .B1(new_n462), .B2(new_n454), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n560), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n478), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT90), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT40), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT40), .B1(new_n569), .B2(new_n570), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n510), .B(new_n557), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT92), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n569), .A2(new_n570), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT40), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT40), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n526), .A2(new_n528), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n507), .A2(new_n509), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n501), .B(new_n502), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT92), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n556), .B1(new_n575), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT93), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n574), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n580), .A2(new_n584), .A3(KEYINPUT92), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n555), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT93), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n343), .B1(new_n485), .B2(new_n510), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n544), .A2(new_n588), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n251), .B1(new_n536), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(G71gat), .A2(G78gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT100), .ZN(new_n597));
  NAND2_X1  g396(.A1(G71gat), .A2(G78gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT101), .ZN(new_n600));
  XOR2_X1   g399(.A(G57gat), .B(G64gat), .Z(new_n601));
  INV_X1    g400(.A(new_n598), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n601), .B1(KEYINPUT9), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  OR3_X1    g403(.A1(new_n603), .A2(new_n602), .A3(new_n596), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n606), .A2(KEYINPUT21), .ZN(new_n607));
  XNOR2_X1  g406(.A(G127gat), .B(G155gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n224), .B1(new_n606), .B2(KEYINPUT21), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT102), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n611), .B(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G85gat), .A2(G92gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT7), .ZN(new_n621));
  NAND2_X1  g420(.A1(G99gat), .A2(G106gat), .ZN(new_n622));
  INV_X1    g421(.A(G85gat), .ZN(new_n623));
  INV_X1    g422(.A(G92gat), .ZN(new_n624));
  AOI22_X1  g423(.A1(KEYINPUT8), .A2(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G99gat), .B(G106gat), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n621), .B(new_n625), .C1(KEYINPUT103), .C2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(KEYINPUT103), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n627), .B(new_n628), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n213), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(G190gat), .B(G218gat), .Z(new_n632));
  INV_X1    g431(.A(KEYINPUT104), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT41), .ZN(new_n634));
  NAND2_X1  g433(.A1(G232gat), .A2(G233gat), .ZN(new_n635));
  OAI22_X1  g434(.A1(new_n632), .A2(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n636), .B1(new_n212), .B2(new_n629), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n632), .A2(new_n633), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(G134gat), .B(G162gat), .Z(new_n641));
  NAND2_X1  g440(.A1(new_n635), .A2(new_n634), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n643), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n619), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n606), .B(new_n629), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT105), .ZN(new_n650));
  OR3_X1    g449(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT10), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n650), .B1(new_n649), .B2(KEYINPUT10), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n606), .A2(KEYINPUT10), .A3(new_n629), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(G230gat), .A2(G233gat), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n655), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n649), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G120gat), .B(G148gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(G176gat), .B(G204gat), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n660), .B(new_n661), .Z(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n656), .A2(new_n658), .A3(new_n662), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n595), .A2(new_n648), .A3(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(new_n484), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(G1gat), .Z(G1324gat));
  XNOR2_X1  g468(.A(KEYINPUT16), .B(G8gat), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n667), .A2(new_n531), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(KEYINPUT42), .Z(new_n672));
  OAI21_X1  g471(.A(G8gat), .B1(new_n667), .B2(new_n531), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT106), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(G1325gat));
  OAI21_X1  g474(.A(G15gat), .B1(new_n667), .B2(new_n544), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n524), .A2(G15gat), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n676), .B1(new_n667), .B2(new_n677), .ZN(G1326gat));
  NOR2_X1   g477(.A1(new_n667), .A2(new_n525), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT43), .B(G22gat), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  INV_X1    g480(.A(KEYINPUT107), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n593), .B1(new_n591), .B2(KEYINPUT93), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n524), .A2(new_n537), .B1(new_n541), .B2(new_n542), .ZN(new_n684));
  AOI211_X1 g483(.A(new_n587), .B(new_n555), .C1(new_n589), .C2(new_n590), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n534), .B1(new_n513), .B2(KEYINPUT35), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n682), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n536), .A2(KEYINPUT107), .A3(new_n594), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n646), .A2(KEYINPUT44), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n647), .B1(new_n686), .B2(new_n687), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT44), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n666), .A2(new_n619), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n251), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G29gat), .B1(new_n697), .B2(new_n484), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n646), .B1(new_n536), .B2(new_n594), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n699), .A2(new_n202), .A3(new_n485), .A4(new_n696), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT45), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n698), .A2(new_n701), .ZN(G1328gat));
  OAI21_X1  g501(.A(G36gat), .B1(new_n697), .B2(new_n531), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n695), .A2(new_n646), .ZN(new_n704));
  AOI21_X1  g503(.A(G36gat), .B1(KEYINPUT108), .B2(KEYINPUT46), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n595), .A2(new_n510), .A3(new_n704), .A4(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT109), .ZN(G1329gat));
  INV_X1    g509(.A(G43gat), .ZN(new_n711));
  INV_X1    g510(.A(new_n524), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n595), .A2(new_n711), .A3(new_n712), .A4(new_n704), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(KEYINPUT110), .B2(KEYINPUT47), .ZN(new_n714));
  AOI211_X1 g513(.A(new_n251), .B(new_n695), .C1(new_n691), .C2(new_n693), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n684), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n714), .B1(new_n716), .B2(G43gat), .ZN(new_n717));
  NAND2_X1  g516(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n717), .B(new_n718), .Z(G1330gat));
  NAND2_X1  g518(.A1(new_n715), .A2(new_n343), .ZN(new_n720));
  INV_X1    g519(.A(G50gat), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n343), .A2(new_n721), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n722), .A2(KEYINPUT111), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n704), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n724), .B1(KEYINPUT111), .B2(new_n722), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n720), .A2(G50gat), .B1(new_n595), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g526(.A1(new_n688), .A2(new_n689), .ZN(new_n728));
  INV_X1    g527(.A(new_n666), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n251), .A2(new_n648), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n485), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g533(.A1(new_n731), .A2(new_n531), .ZN(new_n735));
  NOR2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  AND2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n735), .B2(new_n736), .ZN(G1333gat));
  OAI21_X1  g538(.A(G71gat), .B1(new_n731), .B2(new_n544), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n524), .A2(G71gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n731), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1334gat));
  NOR2_X1   g543(.A1(new_n731), .A2(new_n525), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(new_n323), .ZN(G1335gat));
  INV_X1    g545(.A(KEYINPUT114), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n251), .A2(new_n619), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n748), .A2(KEYINPUT113), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n748), .A2(KEYINPUT113), .ZN(new_n750));
  OR2_X1    g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n729), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n747), .B1(new_n694), .B2(new_n753), .ZN(new_n754));
  AOI211_X1 g553(.A(KEYINPUT114), .B(new_n752), .C1(new_n691), .C2(new_n693), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(G85gat), .B1(new_n757), .B2(new_n484), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n749), .A2(new_n750), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n759), .B1(new_n699), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n692), .A2(KEYINPUT115), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT51), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n729), .A2(new_n623), .A3(new_n485), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n758), .B1(new_n764), .B2(new_n765), .ZN(G1336gat));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n694), .A2(new_n753), .ZN(new_n768));
  OAI21_X1  g567(.A(G92gat), .B1(new_n768), .B2(new_n531), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n666), .A2(G92gat), .A3(new_n531), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n767), .B(new_n769), .C1(new_n764), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n510), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n751), .B1(new_n692), .B2(KEYINPUT115), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n536), .A2(new_n594), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n760), .B1(new_n775), .B2(new_n647), .ZN(new_n776));
  NOR2_X1   g575(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n774), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n777), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n761), .B2(new_n762), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  AOI22_X1  g580(.A1(new_n773), .A2(G92gat), .B1(new_n781), .B2(new_n770), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n772), .B1(new_n782), .B2(new_n767), .ZN(G1337gat));
  OAI21_X1  g582(.A(G99gat), .B1(new_n757), .B2(new_n544), .ZN(new_n784));
  OR3_X1    g583(.A1(new_n524), .A2(G99gat), .A3(new_n666), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n764), .B2(new_n785), .ZN(G1338gat));
  NOR3_X1   g585(.A1(new_n666), .A2(G106gat), .A3(new_n525), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(new_n778), .B2(new_n780), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT118), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI211_X1 g589(.A(KEYINPUT118), .B(new_n787), .C1(new_n778), .C2(new_n780), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XOR2_X1   g591(.A(KEYINPUT117), .B(G106gat), .Z(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(new_n756), .B2(new_n343), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT53), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n768), .A2(new_n525), .ZN(new_n797));
  INV_X1    g596(.A(new_n787), .ZN(new_n798));
  OAI221_X1 g597(.A(new_n796), .B1(new_n797), .B2(new_n793), .C1(new_n764), .C2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n795), .A2(new_n799), .ZN(G1339gat));
  NOR2_X1   g599(.A1(new_n656), .A2(KEYINPUT54), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n662), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n651), .A2(new_n657), .A3(new_n652), .A4(new_n653), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n656), .A2(KEYINPUT54), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n802), .A2(KEYINPUT55), .A3(new_n804), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n805), .A2(new_n665), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n249), .A2(new_n250), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n804), .B(new_n663), .C1(KEYINPUT54), .C2(new_n656), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n806), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n225), .A2(new_n226), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n230), .A2(new_n231), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n245), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n248), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n729), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n647), .B1(new_n811), .B2(new_n817), .ZN(new_n818));
  AND4_X1   g617(.A1(new_n647), .A2(new_n806), .A3(new_n816), .A4(new_n810), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n619), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n251), .A2(new_n648), .A3(new_n666), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n343), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n484), .A2(new_n510), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n712), .A3(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n824), .A2(new_n370), .A3(new_n251), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n484), .B1(new_n820), .B2(new_n821), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n447), .A2(new_n512), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n531), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n807), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n825), .B1(new_n830), .B2(new_n370), .ZN(G1340gat));
  NOR3_X1   g630(.A1(new_n824), .A2(new_n368), .A3(new_n666), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n829), .A2(new_n729), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(new_n833), .B2(new_n368), .ZN(G1341gat));
  OAI21_X1  g633(.A(G127gat), .B1(new_n824), .B2(new_n619), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n619), .A2(G127gat), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n828), .B2(new_n836), .ZN(G1342gat));
  NOR3_X1   g636(.A1(new_n828), .A2(G134gat), .A3(new_n646), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT56), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  OAI21_X1  g640(.A(G134gat), .B1(new_n824), .B2(new_n646), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n842), .A2(KEYINPUT119), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(KEYINPUT119), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n840), .B(new_n841), .C1(new_n843), .C2(new_n844), .ZN(G1343gat));
  NOR2_X1   g644(.A1(new_n684), .A2(new_n525), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n826), .A2(new_n531), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n255), .A3(new_n807), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT120), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n808), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n802), .A2(KEYINPUT120), .A3(new_n804), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n852), .A3(new_n809), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n806), .A2(new_n807), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n647), .B1(new_n854), .B2(new_n817), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n619), .B1(new_n855), .B2(new_n819), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI211_X1 g657(.A(KEYINPUT121), .B(new_n619), .C1(new_n855), .C2(new_n819), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n858), .A2(new_n821), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n849), .B1(new_n860), .B2(new_n343), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n820), .A2(new_n821), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n849), .A3(new_n343), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n544), .A2(new_n823), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n861), .A2(new_n251), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n848), .B1(new_n867), .B2(new_n255), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT58), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n848), .B(new_n870), .C1(new_n867), .C2(new_n255), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(G1344gat));
  NAND3_X1  g671(.A1(new_n847), .A2(new_n257), .A3(new_n729), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n861), .A2(new_n866), .ZN(new_n874));
  AOI211_X1 g673(.A(KEYINPUT59), .B(new_n257), .C1(new_n874), .C2(new_n729), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n862), .A2(new_n343), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n856), .A2(new_n821), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n525), .A2(KEYINPUT57), .ZN(new_n879));
  AOI22_X1  g678(.A1(new_n877), .A2(KEYINPUT57), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n729), .A3(new_n865), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n876), .B1(new_n881), .B2(G148gat), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n873), .B1(new_n875), .B2(new_n882), .ZN(G1345gat));
  INV_X1    g682(.A(new_n874), .ZN(new_n884));
  OAI21_X1  g683(.A(G155gat), .B1(new_n884), .B2(new_n619), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n847), .A2(new_n295), .A3(new_n618), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1346gat));
  OAI21_X1  g686(.A(new_n269), .B1(new_n884), .B2(new_n646), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n847), .A2(new_n294), .A3(new_n647), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(G1347gat));
  AOI21_X1  g689(.A(new_n485), .B1(new_n820), .B2(new_n821), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n891), .A2(new_n510), .A3(new_n827), .ZN(new_n892));
  AOI21_X1  g691(.A(G169gat), .B1(new_n892), .B2(new_n807), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n822), .A2(new_n484), .A3(new_n510), .A4(new_n712), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n894), .A2(new_n393), .A3(new_n251), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n893), .A2(new_n895), .ZN(G1348gat));
  NAND3_X1  g695(.A1(new_n892), .A2(new_n394), .A3(new_n729), .ZN(new_n897));
  OAI21_X1  g696(.A(G176gat), .B1(new_n894), .B2(new_n666), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1349gat));
  NAND4_X1  g698(.A1(new_n892), .A2(new_n382), .A3(new_n384), .A4(new_n618), .ZN(new_n900));
  OAI21_X1  g699(.A(G183gat), .B1(new_n894), .B2(new_n619), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g702(.A1(new_n892), .A2(new_n385), .A3(new_n647), .ZN(new_n904));
  OAI21_X1  g703(.A(G190gat), .B1(new_n894), .B2(new_n646), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(KEYINPUT61), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(KEYINPUT61), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(G1351gat));
  NAND2_X1  g707(.A1(new_n846), .A2(new_n510), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n909), .A2(KEYINPUT122), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n891), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(KEYINPUT122), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n251), .A2(G197gat), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT123), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n544), .A2(new_n484), .A3(new_n510), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT124), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n880), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(G197gat), .B1(new_n918), .B2(new_n251), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n915), .A2(new_n919), .ZN(G1352gat));
  INV_X1    g719(.A(G204gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n880), .A2(new_n729), .A3(new_n917), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n924), .B1(new_n923), .B2(new_n922), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n911), .A2(new_n912), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n729), .A2(new_n921), .ZN(new_n927));
  XOR2_X1   g726(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  OR3_X1    g728(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n929), .B1(new_n926), .B2(new_n927), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n925), .A2(new_n930), .A3(new_n931), .ZN(G1353gat));
  OR3_X1    g731(.A1(new_n926), .A2(G211gat), .A3(new_n619), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n880), .A2(new_n618), .A3(new_n917), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n934), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT63), .B1(new_n934), .B2(G211gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(G1354gat));
  INV_X1    g736(.A(G218gat), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n918), .A2(new_n938), .A3(new_n646), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n926), .B2(new_n646), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n940), .A2(KEYINPUT127), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(KEYINPUT127), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(G1355gat));
endmodule


