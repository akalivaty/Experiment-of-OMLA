//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n551, new_n553,
    new_n554, new_n555, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n564, new_n565, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1137, new_n1138;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT65), .Z(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n451), .ZN(new_n456));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  AOI22_X1  g032(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  XNOR2_X1  g033(.A(KEYINPUT66), .B(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT67), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n460), .A2(new_n463), .A3(G101), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT3), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G137), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n465), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n476), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  OR2_X1    g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  AOI21_X1  g056(.A(new_n470), .B1(new_n459), .B2(KEYINPUT3), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n473), .A2(G136), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n478), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  OR2_X1    g065(.A1(new_n478), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n483), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n482), .A2(new_n497), .A3(G138), .A4(new_n478), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n468), .A2(G138), .A3(new_n478), .A4(new_n471), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT68), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n498), .A2(new_n500), .A3(KEYINPUT4), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n476), .A2(new_n502), .A3(G138), .A4(new_n478), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n496), .B1(new_n501), .B2(new_n503), .ZN(G164));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT6), .B1(new_n510), .B2(KEYINPUT69), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT69), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(G651), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n509), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n511), .A2(new_n514), .A3(G543), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n520), .A2(new_n510), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n519), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XOR2_X1   g099(.A(new_n524), .B(KEYINPUT7), .Z(new_n525));
  NAND2_X1  g100(.A1(new_n509), .A2(KEYINPUT70), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n506), .A2(new_n508), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n525), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n511), .A2(new_n514), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n527), .ZN(new_n534));
  INV_X1    g109(.A(new_n518), .ZN(new_n535));
  AOI22_X1  g110(.A1(G89), .A2(new_n534), .B1(new_n535), .B2(G51), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n532), .A2(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  AOI22_X1  g113(.A1(new_n530), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n510), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT71), .B(G90), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n534), .A2(new_n541), .B1(new_n535), .B2(G52), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  XNOR2_X1  g119(.A(KEYINPUT72), .B(G81), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n534), .A2(new_n545), .B1(new_n535), .B2(G43), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n530), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n547), .B2(new_n510), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  XOR2_X1   g127(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n553));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(new_n535), .A2(G53), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n527), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(G91), .A2(new_n534), .B1(new_n561), .B2(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(G299));
  OAI21_X1  g138(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n564));
  INV_X1    g139(.A(G87), .ZN(new_n565));
  OR3_X1    g140(.A1(new_n515), .A2(KEYINPUT74), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n535), .A2(G49), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT74), .B1(new_n515), .B2(new_n565), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n564), .A2(new_n566), .A3(new_n567), .A4(new_n568), .ZN(G288));
  NAND2_X1  g144(.A1(new_n534), .A2(G86), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n535), .A2(G48), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n570), .B(new_n571), .C1(new_n510), .C2(new_n572), .ZN(new_n573));
  XOR2_X1   g148(.A(new_n573), .B(KEYINPUT75), .Z(G305));
  AOI22_X1  g149(.A1(new_n530), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n510), .ZN(new_n576));
  INV_X1    g151(.A(G85), .ZN(new_n577));
  INV_X1    g152(.A(G47), .ZN(new_n578));
  OAI22_X1  g153(.A1(new_n515), .A2(new_n577), .B1(new_n578), .B2(new_n518), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G290));
  INV_X1    g156(.A(G868), .ZN(new_n582));
  NOR2_X1   g157(.A1(G171), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n534), .A2(G92), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n584), .B(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n510), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(G54), .B2(new_n535), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(G868), .ZN(new_n592));
  OAI21_X1  g167(.A(KEYINPUT76), .B1(new_n583), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(KEYINPUT76), .B2(new_n583), .ZN(G284));
  OAI21_X1  g169(.A(new_n593), .B1(KEYINPUT76), .B2(new_n583), .ZN(G321));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  XOR2_X1   g171(.A(G299), .B(KEYINPUT77), .Z(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G297));
  OAI21_X1  g173(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n591), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n548), .A2(new_n582), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n590), .A2(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(new_n582), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n460), .A2(new_n476), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT13), .Z(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(G2100), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n473), .A2(G135), .ZN(new_n610));
  INV_X1    g185(.A(G123), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n478), .A2(G111), .ZN(new_n612));
  OAI21_X1  g187(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n613));
  OAI221_X1 g188(.A(new_n610), .B1(new_n611), .B2(new_n483), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(KEYINPUT78), .B(G2096), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n608), .A2(G2100), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n609), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT79), .ZN(G156));
  INV_X1    g194(.A(KEYINPUT14), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT15), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2435), .ZN(new_n622));
  XNOR2_X1  g197(.A(G2427), .B(G2438), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n623), .B2(new_n622), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2451), .B(G2454), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT16), .B(G1341), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2443), .B(G2446), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G1348), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n628), .B(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(G14), .B1(new_n625), .B2(new_n631), .ZN(new_n632));
  AND2_X1   g207(.A1(new_n625), .A2(new_n631), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n632), .A2(new_n633), .ZN(G401));
  XOR2_X1   g209(.A(G2084), .B(G2090), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT80), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2072), .B(G2078), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2067), .B(G2678), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT18), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n639), .B(KEYINPUT81), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT82), .B(KEYINPUT17), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n638), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n637), .A2(new_n642), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n646), .B(new_n647), .C1(new_n638), .C2(new_n643), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n641), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2096), .B(G2100), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(G227));
  XOR2_X1   g226(.A(G1956), .B(G2474), .Z(new_n652));
  XOR2_X1   g227(.A(G1961), .B(G1966), .Z(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n652), .A2(new_n653), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT20), .ZN(new_n662));
  OAI221_X1 g237(.A(new_n659), .B1(new_n657), .B2(new_n655), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(new_n661), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT21), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT22), .ZN(new_n666));
  XOR2_X1   g241(.A(G1991), .B(G1996), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT83), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1981), .B(G1986), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G229));
  MUX2_X1   g246(.A(G6), .B(G305), .S(G16), .Z(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT32), .B(G1981), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(G16), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(G22), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(G166), .B2(new_n675), .ZN(new_n677));
  INV_X1    g252(.A(G1971), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n675), .A2(G23), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(G288), .B2(G16), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT33), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT85), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n683), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n679), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n674), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT34), .ZN(new_n688));
  NOR2_X1   g263(.A1(G25), .A2(G29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n473), .A2(G131), .ZN(new_n690));
  INV_X1    g265(.A(G119), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n478), .A2(G107), .ZN(new_n692));
  OAI21_X1  g267(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n693));
  OAI221_X1 g268(.A(new_n690), .B1(new_n691), .B2(new_n483), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT84), .Z(new_n695));
  AOI21_X1  g270(.A(new_n689), .B1(new_n695), .B2(G29), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT35), .B(G1991), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n696), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n675), .A2(G24), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n580), .B2(new_n675), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(G1986), .Z(new_n702));
  NAND3_X1  g277(.A1(new_n688), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT36), .Z(new_n704));
  NOR2_X1   g279(.A1(G29), .A2(G33), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT89), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n473), .A2(G139), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT25), .Z(new_n709));
  AOI22_X1  g284(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n707), .B(new_n709), .C1(new_n478), .C2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT90), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n706), .B1(new_n712), .B2(G29), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(G2072), .Z(new_n714));
  INV_X1    g289(.A(G2084), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT24), .B(G34), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT91), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n480), .B2(new_n717), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n714), .B1(new_n715), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT27), .B(G1996), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n473), .A2(G141), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT92), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n484), .A2(G129), .ZN(new_n725));
  NAND3_X1  g300(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT26), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n460), .A2(G105), .ZN(new_n728));
  NOR4_X1   g303(.A1(new_n724), .A2(new_n725), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G29), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT93), .Z(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G29), .B2(G32), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n721), .B1(new_n722), .B2(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT94), .Z(new_n734));
  AND2_X1   g309(.A1(new_n717), .A2(G26), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n473), .A2(G140), .ZN(new_n736));
  INV_X1    g311(.A(G128), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n478), .A2(G116), .ZN(new_n738));
  OAI21_X1  g313(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n739));
  OAI221_X1 g314(.A(new_n736), .B1(new_n737), .B2(new_n483), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n735), .B1(new_n740), .B2(G29), .ZN(new_n741));
  MUX2_X1   g316(.A(new_n735), .B(new_n741), .S(KEYINPUT28), .Z(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT88), .B(G2067), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n732), .B2(new_n722), .ZN(new_n745));
  NOR2_X1   g320(.A1(G4), .A2(G16), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT86), .Z(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n590), .B2(new_n675), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT87), .B(G1348), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G28), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n751), .A2(KEYINPUT30), .ZN(new_n752));
  AOI21_X1  g327(.A(G29), .B1(new_n751), .B2(KEYINPUT30), .ZN(new_n753));
  OR2_X1    g328(.A1(KEYINPUT31), .A2(G11), .ZN(new_n754));
  NAND2_X1  g329(.A1(KEYINPUT31), .A2(G11), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n752), .A2(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n614), .B2(new_n717), .ZN(new_n757));
  NOR2_X1   g332(.A1(G168), .A2(new_n675), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n675), .B2(G21), .ZN(new_n759));
  INV_X1    g334(.A(G1966), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n757), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n750), .B(new_n761), .C1(new_n760), .C2(new_n759), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT23), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n675), .A2(G20), .ZN(new_n764));
  AOI211_X1 g339(.A(new_n763), .B(new_n764), .C1(G299), .C2(G16), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n763), .B2(new_n764), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT97), .B(G1956), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n675), .A2(G19), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n549), .B2(new_n675), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(G1341), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n720), .A2(new_n715), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n717), .A2(G35), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G162), .B2(new_n717), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT29), .Z(new_n775));
  INV_X1    g350(.A(G2090), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n771), .B(new_n772), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NOR4_X1   g352(.A1(new_n745), .A2(new_n762), .A3(new_n768), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n775), .A2(new_n776), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n675), .A2(G5), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G171), .B2(new_n675), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT95), .ZN(new_n782));
  INV_X1    g357(.A(G1961), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n779), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n783), .B2(new_n782), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT96), .ZN(new_n786));
  INV_X1    g361(.A(new_n503), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n502), .B1(new_n499), .B2(KEYINPUT68), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n498), .ZN(new_n789));
  OAI21_X1  g364(.A(G29), .B1(new_n789), .B2(new_n496), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n717), .A2(G27), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n786), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n786), .B2(new_n791), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G2078), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n778), .A2(new_n785), .A3(new_n794), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n704), .A2(new_n734), .A3(new_n795), .ZN(G311));
  INV_X1    g371(.A(KEYINPUT98), .ZN(new_n797));
  XNOR2_X1  g372(.A(G311), .B(new_n797), .ZN(G150));
  AOI22_X1  g373(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(new_n510), .ZN(new_n800));
  INV_X1    g375(.A(G93), .ZN(new_n801));
  INV_X1    g376(.A(G55), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n515), .A2(new_n801), .B1(new_n802), .B2(new_n518), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(KEYINPUT99), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT99), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n548), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n805), .A2(KEYINPUT99), .A3(new_n548), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n591), .A2(G559), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n815));
  AOI21_X1  g390(.A(G860), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n815), .B2(new_n814), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n805), .A2(G860), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT37), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n819), .ZN(G145));
  NAND2_X1  g395(.A1(new_n501), .A2(new_n503), .ZN(new_n821));
  INV_X1    g396(.A(new_n496), .ZN(new_n822));
  AOI21_X1  g397(.A(KEYINPUT100), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT100), .ZN(new_n824));
  NOR3_X1   g399(.A1(new_n789), .A2(new_n824), .A3(new_n496), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n740), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n729), .ZN(new_n828));
  INV_X1    g403(.A(new_n712), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n711), .B2(new_n828), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n480), .B(new_n614), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n473), .A2(G142), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n478), .A2(G118), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(G130), .B2(new_n484), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G162), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n832), .B(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n694), .B(new_n607), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(G37), .B1(new_n831), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n831), .B2(new_n841), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT101), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g420(.A(G303), .B(KEYINPUT103), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n580), .ZN(new_n847));
  XNOR2_X1  g422(.A(G305), .B(G288), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT42), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n849), .B(KEYINPUT104), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n851), .B1(new_n852), .B2(KEYINPUT42), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n590), .B(G299), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT102), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT41), .ZN(new_n856));
  INV_X1    g431(.A(G299), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(new_n590), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n855), .B(new_n856), .C1(KEYINPUT102), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n854), .A2(KEYINPUT41), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n811), .B(new_n603), .ZN(new_n862));
  MUX2_X1   g437(.A(new_n854), .B(new_n861), .S(new_n862), .Z(new_n863));
  AND2_X1   g438(.A1(new_n853), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT105), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(new_n863), .B2(new_n853), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n864), .A2(KEYINPUT105), .ZN(new_n867));
  OAI21_X1  g442(.A(G868), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(G868), .B2(new_n804), .ZN(G295));
  OAI21_X1  g444(.A(new_n868), .B1(G868), .B2(new_n804), .ZN(G331));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n871));
  XNOR2_X1  g446(.A(G301), .B(G286), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n873), .A2(new_n810), .A3(new_n809), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n811), .A2(new_n872), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n861), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT106), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n811), .A2(KEYINPUT106), .A3(new_n872), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n854), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n849), .B(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n878), .A2(new_n879), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n854), .A2(new_n856), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n855), .B1(KEYINPUT102), .B2(new_n858), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n887), .B1(new_n888), .B2(new_n856), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n874), .A2(new_n875), .ZN(new_n890));
  OAI22_X1  g465(.A1(new_n886), .A2(new_n889), .B1(new_n854), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n852), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n884), .A2(new_n885), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n871), .B1(new_n893), .B2(KEYINPUT43), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n881), .A2(new_n883), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT107), .B1(new_n895), .B2(G37), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n897), .B(new_n885), .C1(new_n881), .C2(new_n883), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n898), .A3(new_n884), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n894), .B1(new_n899), .B2(KEYINPUT43), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(KEYINPUT43), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n893), .A2(KEYINPUT43), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n901), .B1(new_n905), .B2(new_n871), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n903), .B1(new_n899), .B2(KEYINPUT43), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n907), .A2(KEYINPUT108), .A3(KEYINPUT44), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n900), .B1(new_n906), .B2(new_n908), .ZN(G397));
  XOR2_X1   g484(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(new_n826), .B2(G1384), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n465), .A2(G40), .A3(new_n479), .A4(new_n474), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n914), .B(KEYINPUT110), .Z(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n740), .B(G2067), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n915), .A2(new_n729), .ZN(new_n919));
  INV_X1    g494(.A(G1996), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n914), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT46), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n918), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT47), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n919), .A2(new_n920), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n914), .A2(new_n920), .A3(new_n729), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n694), .B(new_n697), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n916), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n925), .A2(new_n926), .A3(new_n918), .A4(new_n928), .ZN(new_n929));
  NOR4_X1   g504(.A1(new_n912), .A2(G1986), .A3(G290), .A4(new_n913), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT48), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n924), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n695), .A2(new_n698), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n925), .A2(new_n926), .A3(new_n918), .A4(new_n933), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n740), .A2(G2067), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n915), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT127), .ZN(new_n938));
  AOI21_X1  g513(.A(G1384), .B1(new_n821), .B2(new_n822), .ZN(new_n939));
  INV_X1    g514(.A(new_n913), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G8), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G1976), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n944), .B1(new_n945), .B2(G288), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT52), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT52), .B1(G288), .B2(new_n945), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n944), .B(new_n948), .C1(new_n945), .C2(G288), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT113), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(KEYINPUT113), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n573), .A2(G1981), .ZN(new_n952));
  XOR2_X1   g527(.A(new_n952), .B(KEYINPUT116), .Z(new_n953));
  XNOR2_X1  g528(.A(KEYINPUT114), .B(G1981), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n573), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT115), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT49), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n953), .A2(KEYINPUT49), .A3(new_n956), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n944), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n951), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n950), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(G303), .A2(G8), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT55), .ZN(new_n965));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n789), .B2(new_n496), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n913), .B1(new_n967), .B2(KEYINPUT50), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n969), .B(new_n966), .C1(new_n789), .C2(new_n496), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n971), .A2(G2090), .ZN(new_n972));
  OAI211_X1 g547(.A(KEYINPUT45), .B(new_n966), .C1(new_n823), .C2(new_n825), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT111), .B1(new_n939), .B2(new_n910), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n975), .B(new_n911), .C1(G164), .C2(G1384), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n973), .A2(new_n974), .A3(new_n940), .A4(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n972), .B1(new_n678), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n965), .B1(new_n978), .B2(new_n943), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n940), .B1(new_n939), .B2(new_n969), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n970), .A2(KEYINPUT112), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n970), .A2(KEYINPUT112), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n776), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n977), .A2(new_n678), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n943), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n965), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n963), .A2(new_n979), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n940), .B1(new_n939), .B2(KEYINPUT45), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n913), .B1(new_n967), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT117), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n939), .A2(new_n910), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n993), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n998), .A2(new_n760), .B1(new_n983), .B2(new_n715), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT124), .B1(new_n999), .B2(new_n943), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n997), .B1(new_n995), .B2(KEYINPUT117), .ZN(new_n1001));
  AOI211_X1 g576(.A(new_n992), .B(new_n913), .C1(new_n967), .C2(new_n994), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n760), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n970), .A2(KEYINPUT112), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n970), .A2(KEYINPUT112), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n715), .B(new_n968), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n943), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT124), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(G168), .A2(new_n943), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(KEYINPUT51), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1000), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1013));
  OAI211_X1 g588(.A(KEYINPUT51), .B(G8), .C1(new_n1013), .C2(G286), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT123), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g591(.A(KEYINPUT123), .B(KEYINPUT51), .C1(new_n1007), .C2(new_n1010), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1012), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT62), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1013), .A2(new_n1010), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1019), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n977), .B2(G2078), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n968), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n783), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1023), .A2(G2078), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n993), .A2(new_n996), .A3(new_n997), .A4(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1024), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(G171), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT125), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT125), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n1032), .A3(G171), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1021), .A2(new_n1022), .A3(new_n1035), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n976), .A2(new_n940), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT56), .B(G2072), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1037), .A2(new_n973), .A3(new_n974), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1956), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n971), .A2(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n558), .A2(KEYINPUT57), .A3(new_n562), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT57), .B1(new_n558), .B2(new_n562), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1039), .A2(new_n1041), .A3(new_n1046), .ZN(new_n1047));
  OR3_X1    g622(.A1(new_n1042), .A2(new_n1044), .A3(KEYINPUT119), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT119), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1050), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1051), .B(KEYINPUT120), .ZN(new_n1052));
  INV_X1    g627(.A(G1348), .ZN(new_n1053));
  INV_X1    g628(.A(G2067), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1025), .A2(new_n1053), .B1(new_n1054), .B2(new_n942), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(new_n590), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1047), .B1(new_n1052), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT61), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1047), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1046), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1037), .A2(new_n920), .A3(new_n973), .A4(new_n974), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT58), .B(G1341), .Z(new_n1063));
  NAND2_X1  g638(.A1(new_n941), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT59), .B1(new_n1065), .B2(new_n549), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n1067));
  AOI211_X1 g642(.A(new_n1067), .B(new_n548), .C1(new_n1062), .C2(new_n1064), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1025), .A2(new_n1053), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n942), .A2(new_n1054), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1070), .A2(KEYINPUT122), .A3(KEYINPUT60), .A4(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n591), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT122), .B1(new_n1055), .B2(KEYINPUT60), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g650(.A(KEYINPUT60), .B(new_n1071), .C1(new_n983), .C2(G1348), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT122), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(new_n1077), .A3(new_n590), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT60), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1061), .B(new_n1069), .C1(new_n1075), .C2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1047), .A2(KEYINPUT121), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1039), .A2(new_n1085), .A3(new_n1041), .A4(new_n1046), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(KEYINPUT61), .A3(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1052), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1057), .B1(new_n1083), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT54), .B1(new_n1029), .B2(G171), .ZN(new_n1090));
  INV_X1    g665(.A(G2078), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1037), .A2(new_n1091), .A3(new_n973), .A4(new_n974), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1092), .A2(new_n1023), .B1(new_n783), .B2(new_n1025), .ZN(new_n1093));
  XOR2_X1   g668(.A(new_n475), .B(KEYINPUT126), .Z(new_n1094));
  AND3_X1   g669(.A1(new_n479), .A2(G40), .A3(new_n1027), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n912), .A2(new_n973), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(G301), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1090), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1093), .A2(G301), .A3(new_n1096), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1031), .A2(new_n1033), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1098), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1089), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n990), .B1(new_n1036), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT63), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1007), .A2(G168), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1106), .B1(new_n989), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n963), .B1(new_n987), .B2(new_n986), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n988), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1112), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1108), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n963), .A2(new_n1112), .ZN(new_n1116));
  INV_X1    g691(.A(new_n961), .ZN(new_n1117));
  OR2_X1    g692(.A1(G288), .A2(G1976), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n956), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n944), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1116), .A2(new_n1120), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1115), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1105), .A2(new_n1122), .ZN(new_n1123));
  XOR2_X1   g698(.A(new_n580), .B(G1986), .Z(new_n1124));
  AOI21_X1  g699(.A(new_n929), .B1(new_n914), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n938), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1103), .A2(KEYINPUT62), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1127), .A2(new_n1034), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1089), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n989), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1115), .A2(new_n1121), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n938), .B(new_n1125), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n937), .B1(new_n1126), .B2(new_n1134), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g710(.A(G319), .B1(new_n632), .B2(new_n633), .ZN(new_n1137));
  OR3_X1    g711(.A1(G229), .A2(G227), .A3(new_n1137), .ZN(new_n1138));
  NOR3_X1   g712(.A1(new_n1138), .A2(new_n907), .A3(new_n844), .ZN(G308));
  INV_X1    g713(.A(G308), .ZN(G225));
endmodule


