

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786;

  BUF_X1 U369 ( .A(n745), .Z(n750) );
  XOR2_X1 U370 ( .A(n370), .B(n675), .Z(n359) );
  BUF_X1 U371 ( .A(n452), .Z(n432) );
  NOR2_X1 U372 ( .A1(n586), .A2(n719), .ZN(n717) );
  OR2_X1 U373 ( .A1(n748), .A2(G902), .ZN(n382) );
  XNOR2_X1 U374 ( .A(n497), .B(G110), .ZN(n465) );
  BUF_X1 U375 ( .A(n742), .Z(n348) );
  INV_X2 U376 ( .A(G953), .ZN(n534) );
  XNOR2_X2 U377 ( .A(n583), .B(n582), .ZN(n592) );
  INV_X1 U378 ( .A(n584), .ZN(n639) );
  XNOR2_X1 U379 ( .A(n767), .B(n505), .ZN(n526) );
  INV_X2 U380 ( .A(G143), .ZN(n555) );
  XNOR2_X1 U381 ( .A(n505), .B(G125), .ZN(n537) );
  BUF_X2 U382 ( .A(n534), .Z(n771) );
  NAND2_X1 U383 ( .A1(n436), .A2(n434), .ZN(n422) );
  AND2_X1 U384 ( .A1(n607), .A2(n483), .ZN(n395) );
  NOR2_X1 U385 ( .A1(n674), .A2(n596), .ZN(n484) );
  XNOR2_X1 U386 ( .A(n657), .B(KEYINPUT40), .ZN(n786) );
  NAND2_X1 U387 ( .A1(n592), .A2(n591), .ZN(n486) );
  AND2_X1 U388 ( .A1(n459), .A2(n455), .ZN(n454) );
  NOR2_X1 U389 ( .A1(n653), .A2(n652), .ZN(n656) );
  NOR2_X1 U390 ( .A1(n491), .A2(n487), .ZN(n621) );
  NOR2_X1 U391 ( .A1(n639), .A2(n720), .ZN(n598) );
  AND2_X1 U392 ( .A1(n425), .A2(n424), .ZN(n366) );
  XNOR2_X1 U393 ( .A(n506), .B(n526), .ZN(n742) );
  XNOR2_X1 U394 ( .A(n567), .B(n566), .ZN(n605) );
  XNOR2_X1 U395 ( .A(n539), .B(n501), .ZN(n506) );
  XNOR2_X1 U396 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U397 ( .A(n538), .B(n502), .ZN(n571) );
  XNOR2_X1 U398 ( .A(n445), .B(n537), .ZN(n769) );
  NAND2_X1 U399 ( .A1(n771), .A2(G234), .ZN(n451) );
  XNOR2_X1 U400 ( .A(G140), .B(KEYINPUT80), .ZN(n499) );
  XOR2_X1 U401 ( .A(KEYINPUT69), .B(G131), .Z(n556) );
  XNOR2_X2 U402 ( .A(n612), .B(KEYINPUT45), .ZN(n379) );
  NAND2_X2 U403 ( .A1(n393), .A2(n390), .ZN(n612) );
  AND2_X1 U404 ( .A1(n408), .A2(n407), .ZN(n634) );
  NAND2_X1 U405 ( .A1(n692), .A2(KEYINPUT47), .ZN(n407) );
  NOR2_X1 U406 ( .A1(n737), .A2(G953), .ZN(n549) );
  NOR2_X1 U407 ( .A1(G953), .A2(G237), .ZN(n527) );
  NAND2_X1 U408 ( .A1(n378), .A2(n377), .ZN(n665) );
  INV_X1 U409 ( .A(KEYINPUT2), .ZN(n377) );
  NAND2_X1 U410 ( .A1(n457), .A2(n349), .ZN(n453) );
  INV_X1 U411 ( .A(G146), .ZN(n505) );
  XNOR2_X1 U412 ( .A(n409), .B(KEYINPUT28), .ZN(n620) );
  NAND2_X1 U413 ( .A1(n635), .A2(n410), .ZN(n409) );
  NOR2_X1 U414 ( .A1(n622), .A2(n411), .ZN(n410) );
  NOR2_X1 U415 ( .A1(n452), .A2(n472), .ZN(n471) );
  NAND2_X1 U416 ( .A1(n470), .A2(n642), .ZN(n469) );
  NAND2_X1 U417 ( .A1(n466), .A2(G902), .ZN(n424) );
  NAND2_X1 U418 ( .A1(n507), .A2(n541), .ZN(n423) );
  INV_X1 U419 ( .A(KEYINPUT48), .ZN(n441) );
  AND2_X1 U420 ( .A1(n646), .A2(n442), .ZN(n440) );
  XNOR2_X1 U421 ( .A(n504), .B(n571), .ZN(n767) );
  XNOR2_X1 U422 ( .A(n412), .B(n351), .ZN(n586) );
  OR2_X1 U423 ( .A1(n751), .A2(G902), .ZN(n412) );
  XNOR2_X1 U424 ( .A(G101), .B(G116), .ZN(n523) );
  AND2_X1 U425 ( .A1(n668), .A2(n667), .ZN(n770) );
  XNOR2_X1 U426 ( .A(n429), .B(n769), .ZN(n564) );
  NAND2_X1 U427 ( .A1(n350), .A2(n352), .ZN(n414) );
  OR2_X2 U428 ( .A1(n770), .A2(KEYINPUT2), .ZN(n436) );
  NAND2_X1 U429 ( .A1(n638), .A2(n639), .ZN(n660) );
  XNOR2_X1 U430 ( .A(n623), .B(KEYINPUT110), .ZN(n624) );
  NOR2_X1 U431 ( .A1(n494), .A2(n546), .ZN(n490) );
  INV_X1 U432 ( .A(G472), .ZN(n385) );
  OR2_X1 U433 ( .A1(n671), .A2(G902), .ZN(n386) );
  XNOR2_X1 U434 ( .A(n446), .B(n413), .ZN(n751) );
  XNOR2_X1 U435 ( .A(n448), .B(n447), .ZN(n446) );
  XNOR2_X1 U436 ( .A(n518), .B(n769), .ZN(n413) );
  XNOR2_X1 U437 ( .A(n515), .B(n517), .ZN(n447) );
  XNOR2_X1 U438 ( .A(n383), .B(n575), .ZN(n748) );
  XNOR2_X1 U439 ( .A(n426), .B(KEYINPUT107), .ZN(n607) );
  NOR2_X1 U440 ( .A1(n471), .A2(n469), .ZN(n468) );
  NAND2_X1 U441 ( .A1(n366), .A2(n367), .ZN(n364) );
  INV_X1 U442 ( .A(KEYINPUT46), .ZN(n443) );
  NAND2_X1 U443 ( .A1(n786), .A2(n784), .ZN(n444) );
  INV_X1 U444 ( .A(n666), .ZN(n420) );
  INV_X1 U445 ( .A(G237), .ZN(n540) );
  XNOR2_X1 U446 ( .A(G902), .B(KEYINPUT15), .ZN(n666) );
  INV_X1 U447 ( .A(KEYINPUT8), .ZN(n450) );
  INV_X1 U448 ( .A(G104), .ZN(n554) );
  XNOR2_X1 U449 ( .A(G113), .B(G122), .ZN(n558) );
  XOR2_X1 U450 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n559) );
  INV_X1 U451 ( .A(KEYINPUT77), .ZN(n434) );
  INV_X1 U452 ( .A(KEYINPUT1), .ZN(n508) );
  NAND2_X1 U453 ( .A1(n454), .A2(n453), .ZN(n461) );
  INV_X1 U454 ( .A(KEYINPUT34), .ZN(n460) );
  NAND2_X1 U455 ( .A1(n616), .A2(G953), .ZN(n617) );
  INV_X1 U456 ( .A(n651), .ZN(n411) );
  NOR2_X1 U457 ( .A1(n614), .A2(n719), .ZN(n635) );
  XNOR2_X1 U458 ( .A(n622), .B(n384), .ZN(n584) );
  INV_X1 U459 ( .A(KEYINPUT6), .ZN(n384) );
  XNOR2_X1 U460 ( .A(G107), .B(G104), .ZN(n464) );
  XNOR2_X1 U461 ( .A(n533), .B(n476), .ZN(n481) );
  INV_X1 U462 ( .A(KEYINPUT16), .ZN(n479) );
  XNOR2_X1 U463 ( .A(G128), .B(G110), .ZN(n517) );
  XNOR2_X1 U464 ( .A(n514), .B(n516), .ZN(n448) );
  XNOR2_X1 U465 ( .A(n428), .B(n427), .ZN(n445) );
  INV_X1 U466 ( .A(G140), .ZN(n427) );
  XNOR2_X1 U467 ( .A(KEYINPUT68), .B(KEYINPUT10), .ZN(n428) );
  XOR2_X1 U468 ( .A(KEYINPUT104), .B(KEYINPUT7), .Z(n569) );
  XNOR2_X1 U469 ( .A(G107), .B(KEYINPUT9), .ZN(n568) );
  INV_X1 U470 ( .A(G134), .ZN(n502) );
  NAND2_X1 U471 ( .A1(G234), .A2(G237), .ZN(n547) );
  XNOR2_X1 U472 ( .A(n565), .B(G475), .ZN(n566) );
  NOR2_X1 U473 ( .A1(G902), .A2(n746), .ZN(n567) );
  INV_X1 U474 ( .A(G478), .ZN(n381) );
  XNOR2_X1 U475 ( .A(n437), .B(KEYINPUT99), .ZN(n627) );
  XNOR2_X1 U476 ( .A(n430), .B(n526), .ZN(n671) );
  XNOR2_X1 U477 ( .A(n530), .B(n525), .ZN(n430) );
  NAND2_X1 U478 ( .A1(G953), .A2(G224), .ZN(n754) );
  NAND2_X1 U479 ( .A1(n756), .A2(G953), .ZN(n763) );
  INV_X1 U480 ( .A(n436), .ZN(n435) );
  AND2_X1 U481 ( .A1(n388), .A2(n387), .ZN(n641) );
  NAND2_X1 U482 ( .A1(n649), .A2(n621), .ZN(n692) );
  NAND2_X1 U483 ( .A1(n775), .A2(G953), .ZN(n776) );
  XNOR2_X1 U484 ( .A(n752), .B(n751), .ZN(n375) );
  XNOR2_X1 U485 ( .A(n749), .B(n748), .ZN(n376) );
  INV_X1 U486 ( .A(KEYINPUT60), .ZN(n398) );
  XNOR2_X1 U487 ( .A(n744), .B(n743), .ZN(n374) );
  INV_X1 U488 ( .A(KEYINPUT56), .ZN(n400) );
  NOR2_X1 U489 ( .A1(n584), .A2(n358), .ZN(n349) );
  AND2_X1 U490 ( .A1(n421), .A2(KEYINPUT64), .ZN(n350) );
  XNOR2_X1 U491 ( .A(n520), .B(KEYINPUT25), .ZN(n351) );
  AND2_X1 U492 ( .A1(n419), .A2(n665), .ZN(n352) );
  XOR2_X1 U493 ( .A(n543), .B(n542), .Z(n353) );
  XNOR2_X1 U494 ( .A(n613), .B(KEYINPUT83), .ZN(n354) );
  NAND2_X1 U495 ( .A1(n618), .A2(n551), .ZN(n355) );
  AND2_X1 U496 ( .A1(n380), .A2(n670), .ZN(n356) );
  AND2_X1 U497 ( .A1(n459), .A2(n458), .ZN(n357) );
  XOR2_X1 U498 ( .A(n532), .B(KEYINPUT88), .Z(n358) );
  XNOR2_X1 U499 ( .A(n746), .B(KEYINPUT59), .ZN(n360) );
  XOR2_X1 U500 ( .A(n671), .B(KEYINPUT62), .Z(n361) );
  AND2_X1 U501 ( .A1(n597), .A2(KEYINPUT86), .ZN(n362) );
  INV_X1 U502 ( .A(n753), .ZN(n404) );
  XNOR2_X1 U503 ( .A(n612), .B(KEYINPUT45), .ZN(n363) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n439) );
  NAND2_X1 U505 ( .A1(n440), .A2(n439), .ZN(n438) );
  XNOR2_X1 U506 ( .A(n438), .B(n441), .ZN(n668) );
  XNOR2_X1 U507 ( .A(n473), .B(KEYINPUT106), .ZN(n462) );
  NAND2_X1 U508 ( .A1(n489), .A2(n355), .ZN(n488) );
  NOR2_X1 U509 ( .A1(n771), .A2(G952), .ZN(n753) );
  NAND2_X1 U510 ( .A1(n534), .A2(G224), .ZN(n372) );
  NAND2_X1 U511 ( .A1(n391), .A2(n611), .ZN(n390) );
  NAND2_X1 U512 ( .A1(n366), .A2(n367), .ZN(n619) );
  INV_X1 U513 ( .A(n396), .ZN(n365) );
  INV_X1 U514 ( .A(n396), .ZN(n463) );
  XNOR2_X1 U515 ( .A(n449), .B(n574), .ZN(n383) );
  XNOR2_X1 U516 ( .A(n557), .B(n554), .ZN(n429) );
  OR2_X1 U517 ( .A1(n742), .A2(n423), .ZN(n367) );
  NAND2_X1 U518 ( .A1(n474), .A2(n598), .ZN(n473) );
  NOR2_X2 U519 ( .A1(n628), .A2(n630), .ZN(n695) );
  BUF_X1 U520 ( .A(n462), .Z(n368) );
  INV_X1 U521 ( .A(n463), .ZN(n369) );
  BUF_X1 U522 ( .A(n676), .Z(n370) );
  NAND2_X1 U523 ( .A1(n419), .A2(n665), .ZN(n418) );
  XNOR2_X1 U524 ( .A(n619), .B(n508), .ZN(n371) );
  XNOR2_X1 U525 ( .A(n364), .B(n508), .ZN(n585) );
  BUF_X1 U526 ( .A(n610), .Z(n781) );
  NOR2_X1 U527 ( .A1(n456), .A2(n603), .ZN(n455) );
  NOR2_X1 U528 ( .A1(n604), .A2(n603), .ZN(n683) );
  INV_X1 U529 ( .A(n706), .ZN(n494) );
  NAND2_X1 U530 ( .A1(n494), .A2(n546), .ZN(n492) );
  XNOR2_X1 U531 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n546) );
  XNOR2_X1 U532 ( .A(n373), .B(n372), .ZN(n536) );
  XNOR2_X2 U533 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n373) );
  NAND2_X2 U534 ( .A1(n415), .A2(n414), .ZN(n745) );
  NOR2_X1 U535 ( .A1(n374), .A2(n753), .ZN(G54) );
  NOR2_X1 U536 ( .A1(n375), .A2(n753), .ZN(G66) );
  NOR2_X1 U537 ( .A1(n376), .A2(n753), .ZN(G63) );
  NAND2_X1 U538 ( .A1(n392), .A2(KEYINPUT86), .ZN(n391) );
  NAND2_X1 U539 ( .A1(n379), .A2(n496), .ZN(n664) );
  NAND2_X1 U540 ( .A1(n379), .A2(n770), .ZN(n669) );
  INV_X1 U541 ( .A(n363), .ZN(n378) );
  NAND2_X1 U542 ( .A1(n363), .A2(n771), .ZN(n759) );
  NAND2_X1 U543 ( .A1(n380), .A2(n422), .ZN(n421) );
  NAND2_X1 U544 ( .A1(n669), .A2(KEYINPUT77), .ZN(n380) );
  XNOR2_X2 U545 ( .A(n382), .B(n381), .ZN(n606) );
  XNOR2_X2 U546 ( .A(n386), .B(n385), .ZN(n622) );
  INV_X1 U547 ( .A(n640), .ZN(n387) );
  XNOR2_X1 U548 ( .A(n389), .B(KEYINPUT36), .ZN(n388) );
  NOR2_X1 U549 ( .A1(n660), .A2(n463), .ZN(n389) );
  NAND2_X1 U550 ( .A1(n609), .A2(n608), .ZN(n392) );
  NAND2_X1 U551 ( .A1(n394), .A2(n482), .ZN(n393) );
  NAND2_X1 U552 ( .A1(n395), .A2(n484), .ZN(n394) );
  NAND2_X1 U553 ( .A1(n396), .A2(n490), .ZN(n489) );
  XNOR2_X2 U554 ( .A(n544), .B(n353), .ZN(n396) );
  NAND2_X1 U555 ( .A1(n365), .A2(n546), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n463), .B(KEYINPUT38), .ZN(n707) );
  NAND2_X1 U557 ( .A1(n631), .A2(n369), .ZN(n632) );
  XNOR2_X1 U558 ( .A(n539), .B(n480), .ZN(n676) );
  XNOR2_X1 U559 ( .A(n397), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U560 ( .A1(n402), .A2(n404), .ZN(n397) );
  XNOR2_X1 U561 ( .A(n399), .B(n398), .ZN(G60) );
  NAND2_X1 U562 ( .A1(n403), .A2(n404), .ZN(n399) );
  XNOR2_X1 U563 ( .A(n401), .B(n400), .ZN(G51) );
  NAND2_X1 U564 ( .A1(n405), .A2(n404), .ZN(n401) );
  XNOR2_X1 U565 ( .A(n672), .B(n361), .ZN(n402) );
  XNOR2_X1 U566 ( .A(n747), .B(n360), .ZN(n403) );
  XNOR2_X1 U567 ( .A(n677), .B(n359), .ZN(n405) );
  XNOR2_X2 U568 ( .A(n406), .B(n521), .ZN(n599) );
  NAND2_X1 U569 ( .A1(n585), .A2(n717), .ZN(n406) );
  NAND2_X1 U570 ( .A1(n462), .A2(n475), .ZN(n426) );
  AND2_X2 U571 ( .A1(n664), .A2(n420), .ZN(n419) );
  NOR2_X1 U572 ( .A1(n633), .A2(n354), .ZN(n408) );
  AND2_X2 U573 ( .A1(n416), .A2(n417), .ZN(n415) );
  NAND2_X1 U574 ( .A1(n356), .A2(n422), .ZN(n416) );
  NAND2_X1 U575 ( .A1(n418), .A2(n670), .ZN(n417) );
  NAND2_X1 U576 ( .A1(n665), .A2(n664), .ZN(n700) );
  NAND2_X1 U577 ( .A1(n742), .A2(n466), .ZN(n425) );
  XNOR2_X2 U578 ( .A(n601), .B(KEYINPUT31), .ZN(n452) );
  XNOR2_X1 U579 ( .A(n461), .B(n460), .ZN(n578) );
  NOR2_X2 U580 ( .A1(n491), .A2(n488), .ZN(n553) );
  XNOR2_X2 U581 ( .A(n431), .B(KEYINPUT35), .ZN(n610) );
  NAND2_X1 U582 ( .A1(n578), .A2(n577), .ZN(n431) );
  XNOR2_X1 U583 ( .A(n433), .B(n481), .ZN(n480) );
  XNOR2_X1 U584 ( .A(n478), .B(n477), .ZN(n433) );
  NOR2_X1 U585 ( .A1(n700), .A2(n435), .ZN(n704) );
  NAND2_X1 U586 ( .A1(n717), .A2(n602), .ZN(n437) );
  XNOR2_X1 U587 ( .A(n634), .B(KEYINPUT82), .ZN(n442) );
  NAND2_X1 U588 ( .A1(n573), .A2(G217), .ZN(n449) );
  XNOR2_X2 U589 ( .A(n451), .B(n450), .ZN(n573) );
  NAND2_X1 U590 ( .A1(n432), .A2(KEYINPUT101), .ZN(n467) );
  NAND2_X1 U591 ( .A1(n432), .A2(n697), .ZN(n698) );
  NAND2_X1 U592 ( .A1(n432), .A2(n695), .ZN(n696) );
  NAND2_X1 U593 ( .A1(n357), .A2(n453), .ZN(n702) );
  INV_X1 U594 ( .A(n458), .ZN(n456) );
  INV_X1 U595 ( .A(n531), .ZN(n457) );
  NAND2_X1 U596 ( .A1(n584), .A2(n358), .ZN(n458) );
  NAND2_X1 U597 ( .A1(n531), .A2(n358), .ZN(n459) );
  XNOR2_X1 U598 ( .A(n368), .B(G101), .ZN(G3) );
  AND2_X1 U599 ( .A1(n463), .A2(n662), .ZN(n673) );
  INV_X1 U600 ( .A(n486), .ZN(n474) );
  XNOR2_X2 U601 ( .A(n465), .B(n464), .ZN(n760) );
  INV_X1 U602 ( .A(n507), .ZN(n466) );
  NAND2_X1 U603 ( .A1(n468), .A2(n467), .ZN(n475) );
  NAND2_X1 U604 ( .A1(n683), .A2(KEYINPUT101), .ZN(n470) );
  OR2_X1 U605 ( .A1(n683), .A2(KEYINPUT101), .ZN(n472) );
  XNOR2_X1 U606 ( .A(n572), .B(n479), .ZN(n476) );
  XNOR2_X1 U607 ( .A(n537), .B(n538), .ZN(n477) );
  XNOR2_X1 U608 ( .A(n536), .B(n535), .ZN(n478) );
  INV_X1 U609 ( .A(n481), .ZN(n762) );
  NAND2_X1 U610 ( .A1(n607), .A2(n362), .ZN(n482) );
  NAND2_X1 U611 ( .A1(n610), .A2(KEYINPUT86), .ZN(n483) );
  XNOR2_X1 U612 ( .A(n486), .B(n485), .ZN(n593) );
  INV_X1 U613 ( .A(KEYINPUT108), .ZN(n485) );
  INV_X1 U614 ( .A(n489), .ZN(n487) );
  NAND2_X1 U615 ( .A1(n493), .A2(n492), .ZN(n491) );
  XNOR2_X1 U616 ( .A(n564), .B(n563), .ZN(n746) );
  XOR2_X1 U617 ( .A(n552), .B(KEYINPUT0), .Z(n495) );
  AND2_X1 U618 ( .A1(n668), .A2(n663), .ZN(n496) );
  INV_X1 U619 ( .A(KEYINPUT109), .ZN(n522) );
  XNOR2_X1 U620 ( .A(n556), .B(n503), .ZN(n504) );
  INV_X1 U621 ( .A(KEYINPUT75), .ZN(n521) );
  XNOR2_X1 U622 ( .A(n529), .B(n533), .ZN(n530) );
  XNOR2_X1 U623 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U624 ( .A(n348), .B(n741), .ZN(n743) );
  XNOR2_X2 U625 ( .A(G101), .B(KEYINPUT76), .ZN(n497) );
  XNOR2_X2 U626 ( .A(n760), .B(KEYINPUT71), .ZN(n539) );
  NAND2_X1 U627 ( .A1(G227), .A2(n771), .ZN(n498) );
  XNOR2_X1 U628 ( .A(n498), .B(KEYINPUT94), .ZN(n500) );
  XNOR2_X2 U629 ( .A(n555), .B(G128), .ZN(n538) );
  XOR2_X1 U630 ( .A(G137), .B(KEYINPUT4), .Z(n503) );
  XNOR2_X1 U631 ( .A(KEYINPUT70), .B(G469), .ZN(n507) );
  NAND2_X1 U632 ( .A1(G234), .A2(n666), .ZN(n509) );
  XNOR2_X1 U633 ( .A(KEYINPUT20), .B(n509), .ZN(n519) );
  AND2_X1 U634 ( .A1(n519), .A2(G221), .ZN(n511) );
  INV_X1 U635 ( .A(KEYINPUT21), .ZN(n510) );
  XNOR2_X1 U636 ( .A(n511), .B(n510), .ZN(n719) );
  XOR2_X1 U637 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n513) );
  XNOR2_X1 U638 ( .A(G137), .B(G119), .ZN(n512) );
  XNOR2_X1 U639 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U640 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n516) );
  XNOR2_X1 U641 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n515) );
  NAND2_X1 U642 ( .A1(G221), .A2(n573), .ZN(n518) );
  NAND2_X1 U643 ( .A1(G217), .A2(n519), .ZN(n520) );
  XNOR2_X1 U644 ( .A(n599), .B(n522), .ZN(n531) );
  XOR2_X1 U645 ( .A(KEYINPUT5), .B(KEYINPUT100), .Z(n524) );
  XOR2_X1 U646 ( .A(n524), .B(n523), .Z(n525) );
  XNOR2_X1 U647 ( .A(n527), .B(KEYINPUT78), .ZN(n560) );
  NAND2_X1 U648 ( .A1(G210), .A2(n560), .ZN(n529) );
  XNOR2_X1 U649 ( .A(G113), .B(KEYINPUT3), .ZN(n528) );
  XNOR2_X1 U650 ( .A(n528), .B(G119), .ZN(n533) );
  XNOR2_X1 U651 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n532) );
  XOR2_X2 U652 ( .A(G116), .B(G122), .Z(n572) );
  XOR2_X1 U653 ( .A(KEYINPUT89), .B(KEYINPUT18), .Z(n535) );
  NAND2_X1 U654 ( .A1(n676), .A2(n666), .ZN(n544) );
  INV_X1 U655 ( .A(G902), .ZN(n541) );
  NAND2_X1 U656 ( .A1(n541), .A2(n540), .ZN(n545) );
  NAND2_X1 U657 ( .A1(n545), .A2(G210), .ZN(n543) );
  INV_X1 U658 ( .A(KEYINPUT91), .ZN(n542) );
  NAND2_X1 U659 ( .A1(n545), .A2(G214), .ZN(n706) );
  XNOR2_X1 U660 ( .A(n547), .B(KEYINPUT14), .ZN(n550) );
  NAND2_X1 U661 ( .A1(G952), .A2(n550), .ZN(n737) );
  INV_X1 U662 ( .A(KEYINPUT92), .ZN(n548) );
  XNOR2_X1 U663 ( .A(n549), .B(n548), .ZN(n618) );
  NAND2_X1 U664 ( .A1(G902), .A2(n550), .ZN(n615) );
  XNOR2_X1 U665 ( .A(KEYINPUT93), .B(G898), .ZN(n756) );
  OR2_X1 U666 ( .A1(n615), .A2(n763), .ZN(n551) );
  INV_X1 U667 ( .A(KEYINPUT87), .ZN(n552) );
  XNOR2_X2 U668 ( .A(n553), .B(n495), .ZN(n603) );
  XNOR2_X1 U669 ( .A(G143), .B(n556), .ZN(n557) );
  XOR2_X1 U670 ( .A(n559), .B(n558), .Z(n562) );
  NAND2_X1 U671 ( .A1(G214), .A2(n560), .ZN(n561) );
  XNOR2_X1 U672 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U673 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n565) );
  INV_X1 U674 ( .A(n605), .ZN(n630) );
  XNOR2_X1 U675 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U676 ( .A(n571), .B(n570), .ZN(n575) );
  XOR2_X1 U677 ( .A(n572), .B(KEYINPUT103), .Z(n574) );
  NOR2_X1 U678 ( .A1(n630), .A2(n606), .ZN(n576) );
  XOR2_X1 U679 ( .A(KEYINPUT81), .B(n576), .Z(n577) );
  INV_X1 U680 ( .A(n606), .ZN(n628) );
  NOR2_X1 U681 ( .A1(n605), .A2(n628), .ZN(n579) );
  XNOR2_X1 U682 ( .A(n579), .B(KEYINPUT105), .ZN(n709) );
  OR2_X2 U683 ( .A1(n709), .A2(n719), .ZN(n580) );
  NOR2_X2 U684 ( .A1(n603), .A2(n580), .ZN(n583) );
  XNOR2_X1 U685 ( .A(KEYINPUT74), .B(KEYINPUT22), .ZN(n581) );
  XNOR2_X1 U686 ( .A(n581), .B(KEYINPUT66), .ZN(n582) );
  INV_X1 U687 ( .A(n371), .ZN(n591) );
  XNOR2_X1 U688 ( .A(KEYINPUT90), .B(n591), .ZN(n640) );
  OR2_X1 U689 ( .A1(n639), .A2(n640), .ZN(n587) );
  INV_X1 U690 ( .A(n586), .ZN(n614) );
  NOR2_X1 U691 ( .A1(n587), .A2(n614), .ZN(n588) );
  NAND2_X1 U692 ( .A1(n592), .A2(n588), .ZN(n590) );
  INV_X1 U693 ( .A(KEYINPUT32), .ZN(n589) );
  XNOR2_X1 U694 ( .A(n590), .B(n589), .ZN(n783) );
  INV_X1 U695 ( .A(KEYINPUT44), .ZN(n597) );
  OR2_X1 U696 ( .A1(n783), .A2(n597), .ZN(n596) );
  NAND2_X1 U697 ( .A1(n593), .A2(n622), .ZN(n594) );
  XNOR2_X1 U698 ( .A(n594), .B(KEYINPUT65), .ZN(n595) );
  INV_X1 U699 ( .A(n614), .ZN(n720) );
  AND2_X2 U700 ( .A1(n595), .A2(n720), .ZN(n674) );
  NOR2_X1 U701 ( .A1(n599), .A2(n622), .ZN(n727) );
  INV_X1 U702 ( .A(n603), .ZN(n600) );
  NAND2_X1 U703 ( .A1(n727), .A2(n600), .ZN(n601) );
  INV_X1 U704 ( .A(n619), .ZN(n602) );
  NAND2_X1 U705 ( .A1(n622), .A2(n627), .ZN(n604) );
  NOR2_X1 U706 ( .A1(n606), .A2(n605), .ZN(n697) );
  INV_X1 U707 ( .A(n697), .ZN(n686) );
  INV_X1 U708 ( .A(n695), .ZN(n691) );
  NAND2_X1 U709 ( .A1(n686), .A2(n691), .ZN(n642) );
  INV_X1 U710 ( .A(n674), .ZN(n609) );
  NOR2_X1 U711 ( .A1(n783), .A2(KEYINPUT44), .ZN(n608) );
  INV_X1 U712 ( .A(n781), .ZN(n611) );
  INV_X1 U713 ( .A(n642), .ZN(n712) );
  NAND2_X1 U714 ( .A1(n712), .A2(KEYINPUT47), .ZN(n613) );
  NOR2_X1 U715 ( .A1(G900), .A2(n615), .ZN(n616) );
  NAND2_X1 U716 ( .A1(n618), .A2(n617), .ZN(n651) );
  NOR2_X1 U717 ( .A1(n620), .A2(n619), .ZN(n649) );
  INV_X1 U718 ( .A(n622), .ZN(n716) );
  NAND2_X1 U719 ( .A1(n716), .A2(n706), .ZN(n625) );
  INV_X1 U720 ( .A(KEYINPUT30), .ZN(n623) );
  NAND2_X1 U721 ( .A1(n627), .A2(n626), .ZN(n652) );
  NAND2_X1 U722 ( .A1(n628), .A2(n651), .ZN(n629) );
  NOR2_X1 U723 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U724 ( .A1(n652), .A2(n632), .ZN(n690) );
  XNOR2_X1 U725 ( .A(n690), .B(KEYINPUT84), .ZN(n633) );
  NAND2_X1 U726 ( .A1(n706), .A2(n651), .ZN(n637) );
  NAND2_X1 U727 ( .A1(n695), .A2(n635), .ZN(n636) );
  NOR2_X1 U728 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U729 ( .A(KEYINPUT112), .B(n641), .ZN(n778) );
  XNOR2_X1 U730 ( .A(KEYINPUT67), .B(KEYINPUT47), .ZN(n643) );
  NAND2_X1 U731 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U732 ( .A1(n692), .A2(n644), .ZN(n645) );
  NOR2_X1 U733 ( .A1(n778), .A2(n645), .ZN(n646) );
  NAND2_X1 U734 ( .A1(n707), .A2(n706), .ZN(n711) );
  NOR2_X1 U735 ( .A1(n709), .A2(n711), .ZN(n648) );
  XNOR2_X1 U736 ( .A(KEYINPUT41), .B(KEYINPUT111), .ZN(n647) );
  XNOR2_X1 U737 ( .A(n648), .B(n647), .ZN(n701) );
  NAND2_X1 U738 ( .A1(n701), .A2(n649), .ZN(n650) );
  XNOR2_X1 U739 ( .A(n650), .B(KEYINPUT42), .ZN(n784) );
  NAND2_X1 U740 ( .A1(n707), .A2(n651), .ZN(n653) );
  XOR2_X1 U741 ( .A(KEYINPUT73), .B(KEYINPUT85), .Z(n654) );
  XNOR2_X1 U742 ( .A(KEYINPUT39), .B(n654), .ZN(n655) );
  XNOR2_X1 U743 ( .A(n656), .B(n655), .ZN(n658) );
  NAND2_X1 U744 ( .A1(n658), .A2(n695), .ZN(n657) );
  NAND2_X1 U745 ( .A1(n697), .A2(n658), .ZN(n659) );
  XNOR2_X1 U746 ( .A(n659), .B(KEYINPUT113), .ZN(n782) );
  OR2_X1 U747 ( .A1(n660), .A2(n371), .ZN(n661) );
  XNOR2_X1 U748 ( .A(n661), .B(KEYINPUT43), .ZN(n662) );
  NOR2_X1 U749 ( .A1(n782), .A2(n673), .ZN(n667) );
  AND2_X1 U750 ( .A1(n667), .A2(KEYINPUT2), .ZN(n663) );
  INV_X1 U751 ( .A(KEYINPUT64), .ZN(n670) );
  NAND2_X1 U752 ( .A1(n745), .A2(G472), .ZN(n672) );
  XOR2_X1 U753 ( .A(n673), .B(G140), .Z(G42) );
  XOR2_X1 U754 ( .A(n674), .B(G110), .Z(G12) );
  NAND2_X1 U755 ( .A1(n745), .A2(G210), .ZN(n677) );
  XNOR2_X1 U756 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n675) );
  NAND2_X1 U757 ( .A1(n683), .A2(n695), .ZN(n678) );
  XNOR2_X1 U758 ( .A(n678), .B(KEYINPUT114), .ZN(n679) );
  XNOR2_X1 U759 ( .A(G104), .B(n679), .ZN(G6) );
  XOR2_X1 U760 ( .A(KEYINPUT27), .B(KEYINPUT116), .Z(n681) );
  XNOR2_X1 U761 ( .A(G107), .B(KEYINPUT26), .ZN(n680) );
  XNOR2_X1 U762 ( .A(n681), .B(n680), .ZN(n682) );
  XOR2_X1 U763 ( .A(KEYINPUT115), .B(n682), .Z(n685) );
  NAND2_X1 U764 ( .A1(n683), .A2(n697), .ZN(n684) );
  XNOR2_X1 U765 ( .A(n685), .B(n684), .ZN(G9) );
  NOR2_X1 U766 ( .A1(n692), .A2(n686), .ZN(n688) );
  XNOR2_X1 U767 ( .A(KEYINPUT29), .B(KEYINPUT117), .ZN(n687) );
  XNOR2_X1 U768 ( .A(n688), .B(n687), .ZN(n689) );
  XOR2_X1 U769 ( .A(G128), .B(n689), .Z(G30) );
  XOR2_X1 U770 ( .A(G143), .B(n690), .Z(G45) );
  NOR2_X1 U771 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U772 ( .A(KEYINPUT118), .B(n693), .Z(n694) );
  XNOR2_X1 U773 ( .A(G146), .B(n694), .ZN(G48) );
  XNOR2_X1 U774 ( .A(n696), .B(G113), .ZN(G15) );
  XOR2_X1 U775 ( .A(G116), .B(KEYINPUT119), .Z(n699) );
  XNOR2_X1 U776 ( .A(n699), .B(n698), .ZN(G18) );
  INV_X1 U777 ( .A(n701), .ZN(n730) );
  NOR2_X1 U778 ( .A1(n730), .A2(n702), .ZN(n703) );
  NOR2_X1 U779 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U780 ( .A1(n705), .A2(n771), .ZN(n739) );
  NOR2_X1 U781 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U782 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U783 ( .A(KEYINPUT123), .B(n710), .Z(n714) );
  NOR2_X1 U784 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U785 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U786 ( .A1(n702), .A2(n715), .ZN(n733) );
  NOR2_X1 U787 ( .A1(n717), .A2(n371), .ZN(n718) );
  XOR2_X1 U788 ( .A(KEYINPUT50), .B(n718), .Z(n724) );
  NAND2_X1 U789 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U790 ( .A(n721), .B(KEYINPUT49), .ZN(n722) );
  XNOR2_X1 U791 ( .A(KEYINPUT121), .B(n722), .ZN(n723) );
  NAND2_X1 U792 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U793 ( .A1(n716), .A2(n725), .ZN(n726) );
  NOR2_X1 U794 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U795 ( .A(n728), .B(KEYINPUT122), .Z(n729) );
  XNOR2_X1 U796 ( .A(KEYINPUT51), .B(n729), .ZN(n731) );
  NOR2_X1 U797 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U798 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U799 ( .A(n734), .B(KEYINPUT124), .ZN(n735) );
  XNOR2_X1 U800 ( .A(KEYINPUT52), .B(n735), .ZN(n736) );
  NOR2_X1 U801 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U802 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U803 ( .A(n740), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U804 ( .A1(n750), .A2(G469), .ZN(n744) );
  XOR2_X1 U805 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n741) );
  NAND2_X1 U806 ( .A1(n745), .A2(G475), .ZN(n747) );
  NAND2_X1 U807 ( .A1(n750), .A2(G478), .ZN(n749) );
  NAND2_X1 U808 ( .A1(n750), .A2(G217), .ZN(n752) );
  XOR2_X1 U809 ( .A(KEYINPUT61), .B(n754), .Z(n755) );
  NOR2_X1 U810 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U811 ( .A(n757), .B(KEYINPUT125), .ZN(n758) );
  NAND2_X1 U812 ( .A1(n759), .A2(n758), .ZN(n766) );
  XNOR2_X1 U813 ( .A(n760), .B(KEYINPUT126), .ZN(n761) );
  XNOR2_X1 U814 ( .A(n762), .B(n761), .ZN(n764) );
  NAND2_X1 U815 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U816 ( .A(n766), .B(n765), .Z(G69) );
  XOR2_X1 U817 ( .A(n767), .B(KEYINPUT94), .Z(n768) );
  XOR2_X1 U818 ( .A(n769), .B(n768), .Z(n773) );
  XOR2_X1 U819 ( .A(n773), .B(n770), .Z(n772) );
  NAND2_X1 U820 ( .A1(n772), .A2(n771), .ZN(n777) );
  XNOR2_X1 U821 ( .A(G227), .B(n773), .ZN(n774) );
  NAND2_X1 U822 ( .A1(n774), .A2(G900), .ZN(n775) );
  NAND2_X1 U823 ( .A1(n777), .A2(n776), .ZN(G72) );
  XNOR2_X1 U824 ( .A(KEYINPUT120), .B(KEYINPUT37), .ZN(n779) );
  XNOR2_X1 U825 ( .A(n779), .B(n778), .ZN(n780) );
  XNOR2_X1 U826 ( .A(G125), .B(n780), .ZN(G27) );
  XOR2_X1 U827 ( .A(G122), .B(n781), .Z(G24) );
  XOR2_X1 U828 ( .A(G134), .B(n782), .Z(G36) );
  XOR2_X1 U829 ( .A(G119), .B(n783), .Z(G21) );
  XOR2_X1 U830 ( .A(G137), .B(n784), .Z(n785) );
  XNOR2_X1 U831 ( .A(KEYINPUT127), .B(n785), .ZN(G39) );
  XNOR2_X1 U832 ( .A(G131), .B(n786), .ZN(G33) );
endmodule

