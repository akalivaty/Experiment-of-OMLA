//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304, new_n1305;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(new_n206));
  AOI22_X1  g0006(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n208));
  NAND3_X1  g0008(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT66), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(KEYINPUT66), .B1(new_n207), .B2(new_n208), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n206), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT1), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n202), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT65), .ZN(new_n222));
  INV_X1    g0022(.A(new_n206), .ZN(new_n223));
  INV_X1    g0023(.A(G13), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NOR3_X1   g0025(.A1(new_n206), .A2(KEYINPUT65), .A3(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  INV_X1    g0029(.A(KEYINPUT0), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n221), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n215), .B(new_n231), .C1(new_n230), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT67), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n238), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(new_n236), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NOR2_X1   g0049(.A1(new_n224), .A2(G1), .ZN(new_n250));
  INV_X1    g0050(.A(G68), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n250), .A2(G20), .A3(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(KEYINPUT12), .ZN(new_n253));
  AND2_X1   g0053(.A1(new_n252), .A2(KEYINPUT12), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n253), .B1(new_n254), .B2(KEYINPUT76), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(KEYINPUT76), .B2(new_n254), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n218), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n257), .A2(G20), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(G68), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n256), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n261), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n219), .A2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G77), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G20), .A2(G33), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n270), .A2(G50), .B1(G20), .B2(new_n251), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n266), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n272), .B(KEYINPUT11), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n265), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n278), .B(KEYINPUT75), .ZN(new_n279));
  INV_X1    g0079(.A(G238), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n276), .A2(KEYINPUT69), .ZN(new_n282));
  INV_X1    g0082(.A(G41), .ZN(new_n283));
  INV_X1    g0083(.A(G45), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT69), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(new_n286), .A3(new_n257), .ZN(new_n287));
  AOI211_X1 g0087(.A(new_n280), .B(new_n281), .C1(new_n282), .C2(new_n287), .ZN(new_n288));
  OR2_X1    g0088(.A1(new_n279), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n218), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT71), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G41), .ZN(new_n292));
  AND3_X1   g0092(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n291), .B1(new_n290), .B2(new_n292), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(KEYINPUT3), .A2(G33), .ZN(new_n297));
  NOR2_X1   g0097(.A1(KEYINPUT3), .A2(G33), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G1698), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n300), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n301));
  INV_X1    g0101(.A(G1698), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT3), .ZN(new_n303));
  INV_X1    g0103(.A(G33), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(KEYINPUT3), .A2(G33), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n302), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G232), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n296), .B1(new_n301), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT13), .B1(new_n289), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n301), .A2(new_n308), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n295), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT13), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n279), .A2(new_n288), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n310), .A2(new_n315), .A3(G179), .ZN(new_n316));
  INV_X1    g0116(.A(G169), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(new_n310), .B2(new_n315), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT14), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AOI211_X1 g0120(.A(KEYINPUT14), .B(new_n317), .C1(new_n310), .C2(new_n315), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n275), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n310), .ZN(new_n323));
  INV_X1    g0123(.A(new_n315), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n323), .A2(new_n324), .A3(G190), .ZN(new_n325));
  AOI21_X1  g0125(.A(G200), .B1(new_n310), .B2(new_n315), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n274), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n263), .A2(G50), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G50), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n262), .A2(new_n331), .B1(new_n332), .B2(new_n259), .ZN(new_n333));
  OAI21_X1  g0133(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n334));
  INV_X1    g0134(.A(G150), .ZN(new_n335));
  INV_X1    g0135(.A(new_n270), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT8), .B(G58), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT72), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G58), .ZN(new_n341));
  OR3_X1    g0141(.A1(new_n339), .A2(new_n341), .A3(KEYINPUT8), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n337), .B1(new_n343), .B2(new_n268), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n333), .B1(new_n344), .B2(new_n266), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n300), .A2(G222), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n307), .A2(G223), .ZN(new_n348));
  INV_X1    g0148(.A(G77), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n305), .A2(new_n306), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n347), .B(new_n348), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n351), .A2(KEYINPUT70), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n295), .B1(new_n351), .B2(KEYINPUT70), .ZN(new_n353));
  OR2_X1    g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n281), .B1(new_n287), .B2(new_n282), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n278), .B1(new_n355), .B2(G226), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(G179), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n356), .B1(new_n352), .B2(new_n353), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G169), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n346), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n354), .A2(G190), .A3(new_n356), .ZN(new_n361));
  XNOR2_X1  g0161(.A(new_n345), .B(KEYINPUT9), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n358), .A2(G200), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT10), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT10), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n361), .A2(new_n362), .A3(new_n366), .A4(new_n363), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n360), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n300), .A2(G232), .B1(G107), .B2(new_n299), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n307), .A2(G238), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n295), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n278), .B1(new_n355), .B2(G244), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G190), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G200), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n262), .A2(G77), .A3(new_n263), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT74), .ZN(new_n382));
  INV_X1    g0182(.A(G87), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT15), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT15), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G87), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT73), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g0189(.A(KEYINPUT15), .B(G87), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n390), .A2(KEYINPUT73), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n268), .ZN(new_n393));
  INV_X1    g0193(.A(new_n338), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(new_n270), .B1(G20), .B2(G77), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n266), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n349), .B2(new_n259), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n380), .A2(new_n382), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n375), .A2(G179), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n374), .A2(G169), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n399), .A2(new_n400), .B1(new_n382), .B2(new_n397), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n329), .A2(new_n368), .A3(new_n398), .A4(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT78), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G87), .ZN(new_n405));
  OAI211_X1 g0205(.A(G223), .B(new_n302), .C1(new_n297), .C2(new_n298), .ZN(new_n406));
  OAI211_X1 g0206(.A(G226), .B(G1698), .C1(new_n297), .C2(new_n298), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT77), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n405), .B(new_n406), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT77), .B1(new_n307), .B2(G226), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n295), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n278), .B1(new_n355), .B2(G232), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n376), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n290), .A2(new_n292), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n286), .B1(new_n285), .B2(new_n257), .ZN(new_n415));
  NOR2_X1   g0215(.A1(G41), .A2(G45), .ZN(new_n416));
  NOR3_X1   g0216(.A1(new_n416), .A2(KEYINPUT69), .A3(G1), .ZN(new_n417));
  OAI211_X1 g0217(.A(G232), .B(new_n414), .C1(new_n415), .C2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n278), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n307), .A2(KEYINPUT77), .A3(G226), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n407), .A2(new_n408), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(new_n405), .A4(new_n406), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n420), .B1(new_n423), .B2(new_n295), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n413), .B1(new_n424), .B2(G200), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n305), .A2(new_n219), .A3(new_n306), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT7), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n305), .A2(KEYINPUT7), .A3(new_n219), .A4(new_n306), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n251), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n341), .A2(new_n251), .ZN(new_n431));
  OAI21_X1  g0231(.A(G20), .B1(new_n431), .B2(new_n201), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n270), .A2(G159), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT16), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT7), .B1(new_n299), .B2(new_n219), .ZN(new_n436));
  INV_X1    g0236(.A(new_n429), .ZN(new_n437));
  OAI21_X1  g0237(.A(G68), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT16), .ZN(new_n439));
  INV_X1    g0239(.A(new_n434), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n435), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n261), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n343), .A2(new_n263), .ZN(new_n444));
  INV_X1    g0244(.A(new_n262), .ZN(new_n445));
  OAI22_X1  g0245(.A1(new_n444), .A2(new_n445), .B1(new_n258), .B2(new_n343), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n425), .A2(new_n443), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n404), .B1(new_n448), .B2(KEYINPUT17), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n446), .B1(new_n442), .B2(new_n261), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT17), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n450), .A2(KEYINPUT78), .A3(new_n451), .A4(new_n425), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n448), .A2(KEYINPUT17), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n266), .B1(new_n435), .B2(new_n441), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n411), .A2(G179), .A3(new_n412), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n317), .B1(new_n411), .B2(new_n412), .ZN(new_n458));
  OAI22_X1  g0258(.A1(new_n456), .A2(new_n446), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g0259(.A(new_n459), .B(KEYINPUT18), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n403), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT90), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n257), .B(G45), .C1(new_n283), .C2(KEYINPUT5), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT82), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n283), .A2(KEYINPUT5), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(new_n465), .B2(new_n466), .ZN(new_n470));
  OAI211_X1 g0270(.A(G270), .B(new_n414), .C1(new_n468), .C2(new_n470), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n465), .A2(new_n466), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n281), .A2(new_n277), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n472), .A2(new_n473), .A3(new_n467), .A4(new_n469), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(G264), .B(G1698), .C1(new_n297), .C2(new_n298), .ZN(new_n476));
  OAI211_X1 g0276(.A(G257), .B(new_n302), .C1(new_n297), .C2(new_n298), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n305), .A2(G303), .A3(new_n306), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT86), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT86), .A4(new_n478), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(new_n295), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n378), .B1(new_n475), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G283), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n304), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G97), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n487), .B(new_n219), .C1(G33), .C2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(G116), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G20), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n261), .A2(KEYINPUT88), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT88), .B1(new_n261), .B2(new_n491), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT20), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n489), .B(KEYINPUT20), .C1(new_n492), .C2(new_n493), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n257), .A2(G33), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n258), .A2(new_n499), .A3(new_n218), .A4(new_n260), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n500), .A2(KEYINPUT87), .A3(new_n490), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT87), .B1(new_n500), .B2(new_n490), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n502), .A2(new_n503), .B1(new_n490), .B2(new_n259), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n464), .B1(new_n484), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n259), .A2(new_n490), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT87), .ZN(new_n508));
  AND4_X1   g0308(.A1(new_n218), .A2(new_n258), .A3(new_n260), .A4(new_n499), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n508), .B1(new_n509), .B2(G116), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n507), .B1(new_n510), .B2(new_n501), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(new_n496), .B2(new_n497), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n481), .A2(new_n295), .A3(new_n482), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n471), .A2(new_n474), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n512), .B(KEYINPUT90), .C1(new_n515), .C2(new_n378), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(G190), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n506), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT21), .ZN(new_n519));
  OAI21_X1  g0319(.A(G169), .B1(new_n513), .B2(new_n514), .ZN(new_n520));
  OAI211_X1 g0320(.A(KEYINPUT89), .B(new_n519), .C1(new_n520), .C2(new_n512), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT89), .B1(new_n520), .B2(new_n512), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT21), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n505), .A2(new_n515), .A3(G179), .ZN(new_n524));
  AND4_X1   g0324(.A1(new_n518), .A2(new_n521), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n259), .A2(new_n488), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n500), .B2(new_n488), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT6), .ZN(new_n528));
  INV_X1    g0328(.A(G107), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n488), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(G97), .A2(G107), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n529), .A2(KEYINPUT6), .A3(G97), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n534), .A2(G20), .B1(G77), .B2(new_n270), .ZN(new_n535));
  OAI21_X1  g0335(.A(G107), .B1(new_n436), .B2(new_n437), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n527), .B1(new_n537), .B2(new_n261), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(G244), .B(new_n302), .C1(new_n297), .C2(new_n298), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT79), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT4), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n541), .B1(new_n540), .B2(new_n542), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT80), .B1(new_n540), .B2(new_n542), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n486), .B1(new_n307), .B2(G250), .ZN(new_n547));
  INV_X1    g0347(.A(G244), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n305), .B2(new_n306), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT80), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(KEYINPUT4), .A4(new_n302), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n546), .A2(new_n547), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n295), .B1(new_n545), .B2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(G257), .B(new_n414), .C1(new_n468), .C2(new_n470), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n554), .A2(new_n474), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(G190), .A3(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT83), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n553), .A2(KEYINPUT83), .A3(G190), .A4(new_n555), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n539), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT81), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n553), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(KEYINPUT81), .B(new_n295), .C1(new_n545), .C2(new_n552), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n563), .A3(new_n555), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G200), .ZN(new_n565));
  INV_X1    g0365(.A(G179), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n562), .A2(new_n566), .A3(new_n563), .A4(new_n555), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n553), .A2(new_n555), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n538), .B1(new_n568), .B2(new_n317), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n560), .A2(new_n565), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n250), .A2(G20), .A3(new_n529), .ZN(new_n571));
  XNOR2_X1  g0371(.A(new_n571), .B(KEYINPUT25), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(G107), .B2(new_n509), .ZN(new_n573));
  OAI21_X1  g0373(.A(KEYINPUT23), .B1(new_n219), .B2(G107), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT23), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n575), .A2(new_n529), .A3(G20), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n219), .A2(G33), .A3(G116), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT91), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n574), .A2(new_n576), .A3(new_n577), .A4(KEYINPUT91), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n219), .B(G87), .C1(new_n297), .C2(new_n298), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT22), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OR2_X1    g0385(.A1(new_n583), .A2(new_n584), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n582), .A2(KEYINPUT24), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n261), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n583), .B(KEYINPUT22), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT24), .B1(new_n589), .B2(new_n582), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n573), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT92), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT92), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n593), .B(new_n573), .C1(new_n588), .C2(new_n590), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n350), .A2(G250), .A3(new_n302), .ZN(new_n595));
  OAI211_X1 g0395(.A(G257), .B(G1698), .C1(new_n297), .C2(new_n298), .ZN(new_n596));
  NAND2_X1  g0396(.A1(G33), .A2(G294), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n295), .ZN(new_n599));
  OAI211_X1 g0399(.A(G264), .B(new_n414), .C1(new_n468), .C2(new_n470), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n474), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n317), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n599), .A2(new_n566), .A3(new_n600), .A4(new_n474), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n592), .A2(new_n594), .A3(new_n604), .ZN(new_n605));
  OR2_X1    g0405(.A1(new_n601), .A2(G190), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n601), .A2(new_n378), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n591), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n509), .A2(G87), .ZN(new_n611));
  XNOR2_X1  g0411(.A(new_n611), .B(KEYINPUT85), .ZN(new_n612));
  NAND2_X1  g0412(.A1(G33), .A2(G97), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT19), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n219), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n383), .A2(new_n488), .A3(new_n529), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n219), .B(G68), .C1(new_n297), .C2(new_n298), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n614), .B1(new_n613), .B2(G20), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n261), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n259), .B1(new_n389), .B2(new_n391), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n612), .A2(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(G238), .B(new_n302), .C1(new_n297), .C2(new_n298), .ZN(new_n625));
  OAI211_X1 g0425(.A(G244), .B(G1698), .C1(new_n297), .C2(new_n298), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n625), .B(new_n626), .C1(new_n304), .C2(new_n490), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n295), .ZN(new_n628));
  OAI21_X1  g0428(.A(G250), .B1(new_n284), .B2(G1), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n257), .A2(G45), .A3(G274), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n281), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n628), .A2(G190), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n628), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G200), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n624), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n387), .A2(new_n388), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n390), .A2(KEYINPUT73), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n509), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n621), .A2(new_n622), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT84), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT84), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n621), .A2(new_n622), .A3(new_n642), .A4(new_n639), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n634), .A2(G169), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n628), .A2(G179), .A3(new_n632), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  AND4_X1   g0448(.A1(new_n605), .A2(new_n610), .A3(new_n636), .A4(new_n648), .ZN(new_n649));
  AND4_X1   g0449(.A1(new_n463), .A2(new_n525), .A3(new_n570), .A4(new_n649), .ZN(G372));
  NAND2_X1  g0450(.A1(new_n365), .A2(new_n367), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n322), .A2(new_n402), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n652), .A2(new_n455), .A3(new_n327), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n651), .B1(new_n653), .B2(new_n460), .ZN(new_n654));
  INV_X1    g0454(.A(new_n360), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n647), .A2(new_n640), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n569), .A2(new_n567), .A3(new_n636), .A4(new_n648), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n658), .B1(new_n659), .B2(KEYINPUT26), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n569), .A2(new_n567), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n591), .B1(new_n606), .B2(new_n607), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n560), .B2(new_n565), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n604), .A2(new_n591), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n523), .A2(new_n521), .A3(new_n524), .A4(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n662), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n636), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n660), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n656), .B1(new_n463), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT93), .ZN(G369));
  INV_X1    g0472(.A(KEYINPUT89), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n317), .B1(new_n475), .B2(new_n483), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n673), .B1(new_n674), .B2(new_n505), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n524), .B1(new_n675), .B2(new_n519), .ZN(new_n676));
  INV_X1    g0476(.A(new_n521), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n250), .ZN(new_n679));
  OR3_X1    g0479(.A1(new_n679), .A2(KEYINPUT27), .A3(G20), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT27), .B1(new_n679), .B2(G20), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G213), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n512), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n678), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n525), .B2(new_n686), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT94), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n605), .A2(new_n685), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n592), .A2(new_n594), .A3(new_n684), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n605), .A2(new_n692), .A3(new_n610), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n685), .B1(new_n676), .B2(new_n677), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(new_n693), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n604), .A2(new_n591), .A3(new_n685), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n697), .A2(new_n702), .ZN(G399));
  NOR2_X1   g0503(.A1(new_n227), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR4_X1   g0505(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G1), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n216), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n605), .A2(new_n523), .A3(new_n521), .A4(new_n524), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n636), .A2(new_n657), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n663), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n570), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n659), .A2(new_n668), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n569), .A2(new_n567), .A3(KEYINPUT26), .A4(new_n636), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n658), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI211_X1 g0517(.A(new_n710), .B(new_n684), .C1(new_n714), .C2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n670), .A2(new_n685), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n718), .B1(new_n710), .B2(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n525), .A2(new_n649), .A3(new_n570), .A4(new_n685), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n475), .A2(new_n483), .ZN(new_n722));
  AOI21_X1  g0522(.A(G179), .B1(new_n628), .B2(new_n632), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n564), .A2(new_n722), .A3(new_n601), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n599), .A2(new_n600), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n722), .A2(new_n725), .A3(new_n646), .ZN(new_n726));
  INV_X1    g0526(.A(new_n568), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT95), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(KEYINPUT30), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  AOI211_X1 g0530(.A(KEYINPUT95), .B(new_n730), .C1(new_n726), .C2(new_n727), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n724), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n684), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n721), .A2(new_n733), .A3(KEYINPUT31), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT31), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n732), .A2(new_n735), .A3(new_n684), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n720), .B1(G330), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n709), .B1(new_n738), .B2(G1), .ZN(G364));
  OR2_X1    g0539(.A1(new_n689), .A2(G330), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n224), .A2(G20), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G45), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n705), .A2(G1), .A3(new_n742), .ZN(new_n743));
  AND3_X1   g0543(.A1(new_n740), .A2(new_n690), .A3(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n743), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n745), .A2(KEYINPUT96), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(KEYINPUT96), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n228), .A2(G355), .A3(new_n350), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n228), .A2(new_n299), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n217), .A2(G45), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n752), .B1(new_n245), .B2(G45), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n750), .B1(G116), .B2(new_n228), .C1(new_n751), .C2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n290), .B1(new_n219), .B2(G169), .ZN(new_n755));
  XOR2_X1   g0555(.A(new_n755), .B(KEYINPUT97), .Z(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n219), .A2(new_n376), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n566), .A2(G200), .ZN(new_n763));
  AND3_X1   g0563(.A1(new_n762), .A2(KEYINPUT98), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(KEYINPUT98), .B1(new_n762), .B2(new_n763), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G58), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n219), .A2(G190), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G179), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G159), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT32), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n762), .A2(new_n566), .A3(G200), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n350), .B1(new_n775), .B2(new_n383), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT99), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n768), .A2(new_n774), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n566), .A2(new_n378), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n762), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n769), .A2(new_n566), .A3(G200), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n783), .A2(G50), .B1(new_n785), .B2(G107), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n781), .A2(new_n769), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n763), .A2(new_n769), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI22_X1  g0590(.A1(G68), .A2(new_n788), .B1(new_n790), .B2(G77), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n219), .B1(new_n770), .B2(G190), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G97), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n786), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n767), .A2(G322), .ZN(new_n796));
  XNOR2_X1  g0596(.A(KEYINPUT33), .B(G317), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n350), .B1(new_n788), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n775), .ZN(new_n799));
  INV_X1    g0599(.A(new_n771), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n799), .A2(G303), .B1(new_n800), .B2(G329), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G283), .A2(new_n785), .B1(new_n790), .B2(G311), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n796), .A2(new_n798), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G326), .ZN(new_n804));
  INV_X1    g0604(.A(G294), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n782), .A2(new_n804), .B1(new_n792), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT100), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n780), .A2(new_n795), .B1(new_n803), .B2(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n754), .A2(new_n761), .B1(new_n757), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n749), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT101), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(new_n688), .B2(new_n760), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n744), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(G396));
  NAND2_X1  g0614(.A1(new_n737), .A2(G330), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n397), .A2(new_n382), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n684), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n398), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n402), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n401), .A2(new_n685), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n719), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n401), .B1(new_n398), .B2(new_n817), .ZN(new_n823));
  INV_X1    g0623(.A(new_n820), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n664), .A2(new_n666), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n669), .B1(new_n826), .B2(new_n661), .ZN(new_n827));
  INV_X1    g0627(.A(new_n660), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n685), .B(new_n825), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n822), .A2(new_n829), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n815), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n815), .A2(new_n830), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n831), .A2(new_n743), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n756), .A2(new_n759), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT102), .Z(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n748), .B1(new_n349), .B2(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G137), .A2(new_n783), .B1(new_n790), .B2(G159), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n335), .B2(new_n787), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(G143), .B2(new_n767), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n840), .A2(KEYINPUT34), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(KEYINPUT34), .ZN(new_n842));
  INV_X1    g0642(.A(G132), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n784), .A2(new_n251), .B1(new_n771), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n350), .B1(new_n775), .B2(new_n332), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n844), .B(new_n845), .C1(G58), .C2(new_n793), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n841), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(G311), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n789), .A2(new_n490), .B1(new_n771), .B2(new_n848), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n350), .B(new_n849), .C1(G87), .C2(new_n785), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n767), .A2(G294), .ZN(new_n851));
  XOR2_X1   g0651(.A(KEYINPUT103), .B(G283), .Z(new_n852));
  OAI22_X1  g0652(.A1(new_n529), .A2(new_n775), .B1(new_n852), .B2(new_n787), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(G303), .B2(new_n783), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n850), .A2(new_n794), .A3(new_n851), .A4(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT104), .B1(new_n847), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n847), .A2(KEYINPUT104), .A3(new_n855), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n757), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n837), .B1(new_n856), .B2(new_n858), .C1(new_n825), .C2(new_n759), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n833), .A2(new_n859), .ZN(G384));
  OAI211_X1 g0660(.A(G116), .B(new_n220), .C1(new_n534), .C2(KEYINPUT35), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(KEYINPUT35), .B2(new_n534), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT36), .ZN(new_n863));
  OR3_X1    g0663(.A1(new_n216), .A2(new_n349), .A3(new_n431), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n332), .A2(G68), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n257), .B(G13), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n450), .A2(new_n682), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n449), .A2(new_n452), .B1(KEYINPUT17), .B2(new_n448), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n868), .B1(new_n869), .B2(new_n460), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n448), .A2(new_n459), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT37), .B1(new_n871), .B2(new_n868), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT105), .B1(new_n450), .B2(new_n682), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT105), .ZN(new_n874));
  INV_X1    g0674(.A(new_n682), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n874), .B(new_n875), .C1(new_n456), .C2(new_n446), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n448), .A2(new_n459), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n872), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n870), .A2(KEYINPUT38), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT107), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n871), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n448), .A2(new_n459), .A3(KEYINPUT107), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n873), .A2(new_n876), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n878), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n448), .A2(new_n878), .A3(new_n459), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n889), .A2(KEYINPUT108), .A3(new_n873), .A4(new_n876), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT108), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n877), .B2(new_n879), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT109), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n448), .A2(KEYINPUT107), .A3(new_n459), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT107), .B1(new_n448), .B2(new_n459), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n887), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT37), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT109), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n898), .A2(new_n899), .A3(new_n892), .A4(new_n890), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n887), .B1(new_n455), .B2(new_n461), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n894), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT38), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n882), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n328), .A2(new_n275), .A3(new_n684), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n322), .B(new_n327), .C1(new_n274), .C2(new_n685), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n821), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n737), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT40), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n908), .A2(new_n734), .A3(new_n736), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT40), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n870), .A2(new_n880), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n904), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n881), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n911), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n910), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n737), .A2(new_n463), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n917), .B(new_n918), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n919), .A2(G330), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n829), .A2(new_n820), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n906), .A2(new_n907), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(new_n915), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n460), .A2(new_n682), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n914), .B2(new_n881), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n905), .B2(new_n925), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n322), .A2(new_n684), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT106), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n923), .B(new_n924), .C1(new_n927), .C2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n656), .B1(new_n720), .B2(new_n463), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n931), .B(new_n932), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n920), .A2(new_n933), .B1(new_n257), .B2(new_n741), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n920), .A2(new_n933), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n867), .B1(new_n934), .B2(new_n935), .ZN(G367));
  OAI21_X1  g0736(.A(new_n570), .B1(new_n538), .B2(new_n685), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n662), .A2(new_n684), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(new_n699), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT42), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n940), .A2(KEYINPUT110), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n661), .B1(new_n937), .B2(new_n605), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n685), .ZN(new_n944));
  OAI21_X1  g0744(.A(KEYINPUT42), .B1(new_n939), .B2(new_n699), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n942), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n940), .A2(new_n941), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT110), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n624), .A2(new_n685), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n657), .ZN(new_n952));
  INV_X1    g0752(.A(new_n712), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n952), .B1(new_n953), .B2(new_n951), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n947), .A2(new_n950), .B1(KEYINPUT43), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(KEYINPUT43), .B2(new_n955), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT43), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n947), .A2(new_n958), .A3(new_n954), .A4(new_n950), .ZN(new_n959));
  INV_X1    g0759(.A(new_n939), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n957), .A2(new_n696), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n957), .A2(new_n959), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n697), .B2(new_n939), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n704), .B(KEYINPUT41), .Z(new_n964));
  NOR2_X1   g0764(.A1(new_n939), .A2(new_n701), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT45), .ZN(new_n966));
  OAI21_X1  g0766(.A(KEYINPUT44), .B1(new_n960), .B2(new_n702), .ZN(new_n967));
  OR3_X1    g0767(.A1(new_n960), .A2(new_n702), .A3(KEYINPUT44), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(KEYINPUT111), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n697), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n699), .A2(KEYINPUT112), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n699), .A2(KEYINPUT112), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n695), .A2(new_n698), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n690), .B(new_n975), .Z(new_n976));
  NAND3_X1  g0776(.A1(new_n969), .A2(KEYINPUT111), .A3(new_n696), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n971), .A2(new_n738), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n964), .B1(new_n978), .B2(new_n738), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n742), .A2(G1), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n961), .B(new_n963), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n954), .A2(new_n760), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n799), .A2(G116), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT46), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n350), .B(new_n985), .C1(G311), .C2(new_n783), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n784), .A2(new_n488), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n852), .A2(new_n789), .B1(new_n787), .B2(new_n805), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(G317), .C2(new_n800), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n983), .A2(new_n984), .B1(new_n793), .B2(G107), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n767), .A2(G303), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n986), .A2(new_n989), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n784), .A2(new_n349), .ZN(new_n993));
  INV_X1    g0793(.A(G137), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n350), .B1(new_n771), .B2(new_n994), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n993), .B(new_n995), .C1(G159), .C2(new_n788), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n793), .A2(G68), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n767), .A2(G150), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n775), .A2(new_n341), .B1(new_n789), .B2(new_n332), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(G143), .B2(new_n783), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n996), .A2(new_n997), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n992), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n756), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n392), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n761), .B1(new_n228), .B2(new_n1006), .C1(new_n751), .C2(new_n241), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n749), .A2(new_n982), .A3(new_n1005), .A4(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n981), .A2(new_n1008), .ZN(G387));
  NAND2_X1  g0809(.A1(new_n976), .A2(new_n738), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1011), .A2(new_n705), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n738), .B2(new_n976), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G322), .A2(new_n783), .B1(new_n790), .B2(G303), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n848), .B2(new_n787), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G317), .B2(new_n767), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT114), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1018), .A2(KEYINPUT48), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1018), .A2(KEYINPUT48), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n775), .A2(new_n805), .B1(new_n852), .B2(new_n792), .ZN(new_n1021));
  NOR3_X1   g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT49), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n299), .B1(new_n771), .B2(new_n804), .C1(new_n490), .C2(new_n784), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n767), .A2(G50), .B1(new_n343), .B2(new_n788), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n1006), .B2(new_n792), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G68), .A2(new_n790), .B1(new_n800), .B2(G150), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n349), .B2(new_n775), .C1(new_n772), .C2(new_n782), .ZN(new_n1029));
  NOR4_X1   g0829(.A1(new_n1027), .A2(new_n1029), .A3(new_n299), .A4(new_n987), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n757), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n236), .A2(G45), .A3(new_n299), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n394), .A2(new_n332), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT50), .ZN(new_n1034));
  AOI211_X1 g0834(.A(G45), .B(new_n1034), .C1(G68), .C2(G77), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n706), .B1(new_n1035), .B2(new_n350), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n227), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n761), .B1(new_n228), .B2(new_n529), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1031), .B(new_n749), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n695), .B2(new_n760), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n976), .B2(new_n980), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1013), .A2(new_n1041), .ZN(G393));
  INV_X1    g0842(.A(KEYINPUT117), .ZN(new_n1043));
  NOR3_X1   g0843(.A1(new_n969), .A2(new_n696), .A3(KEYINPUT115), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n969), .A2(new_n696), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT115), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n969), .A2(new_n696), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1044), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1043), .B1(new_n1050), .B2(new_n1011), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1048), .B1(new_n1046), .B2(new_n1045), .ZN(new_n1052));
  OAI211_X1 g0852(.A(KEYINPUT117), .B(new_n1010), .C1(new_n1052), .C2(new_n1044), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1051), .A2(new_n1053), .A3(new_n704), .A4(new_n978), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n939), .A2(new_n760), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n761), .B1(new_n488), .B2(new_n228), .C1(new_n751), .C2(new_n248), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n749), .A2(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n767), .A2(G311), .B1(G317), .B2(new_n783), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT52), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G303), .A2(new_n788), .B1(new_n800), .B2(G322), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n805), .B2(new_n789), .C1(new_n775), .C2(new_n852), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n299), .B1(new_n792), .B2(new_n490), .C1(new_n784), .C2(new_n529), .ZN(new_n1062));
  OR3_X1    g0862(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n799), .A2(G68), .B1(new_n800), .B2(G143), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1064), .B(new_n350), .C1(new_n383), .C2(new_n784), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT116), .Z(new_n1066));
  OAI22_X1  g0866(.A1(new_n766), .A2(new_n772), .B1(new_n335), .B2(new_n782), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT51), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n793), .A2(G77), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G50), .A2(new_n788), .B1(new_n790), .B2(new_n394), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n756), .B1(new_n1063), .B2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1057), .A2(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1050), .A2(new_n980), .B1(new_n1055), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1054), .A2(new_n1074), .ZN(G390));
  NAND4_X1  g0875(.A1(new_n908), .A2(new_n734), .A3(new_n736), .A4(G330), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  AOI211_X1 g0877(.A(KEYINPUT39), .B(new_n882), .C1(new_n903), .C2(new_n904), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n929), .B1(new_n921), .B2(new_n922), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n1078), .A2(new_n1079), .A3(new_n926), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n684), .B(new_n823), .C1(new_n714), .C2(new_n717), .ZN(new_n1081));
  OAI21_X1  g0881(.A(KEYINPUT118), .B1(new_n1081), .B2(new_n824), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT118), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n714), .A2(new_n717), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n685), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1083), .B(new_n820), .C1(new_n1085), .C2(new_n823), .ZN(new_n1086));
  AND3_X1   g0886(.A1(new_n1082), .A2(new_n922), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n877), .B1(new_n884), .B2(new_n885), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n892), .B(new_n890), .C1(new_n1088), .C2(new_n878), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n901), .B1(new_n1089), .B2(KEYINPUT109), .ZN(new_n1090));
  AOI21_X1  g0890(.A(KEYINPUT38), .B1(new_n1090), .B2(new_n900), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n930), .B1(new_n1091), .B2(new_n882), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1087), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1077), .B1(new_n1080), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1082), .A2(new_n1086), .A3(new_n922), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n903), .A2(new_n904), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n881), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1095), .A2(new_n1097), .A3(new_n930), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n926), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n1097), .B2(KEYINPUT39), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1098), .B(new_n1076), .C1(new_n1100), .C2(new_n1079), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1094), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G1), .B2(new_n742), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G97), .A2(new_n790), .B1(new_n800), .B2(G294), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n485), .B2(new_n782), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(G116), .B2(new_n767), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n785), .A2(G68), .B1(new_n788), .B2(G107), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n350), .B1(new_n799), .B2(G87), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n1107), .A2(new_n1069), .A3(new_n1108), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n350), .B1(new_n792), .B2(new_n772), .C1(new_n784), .C2(new_n332), .ZN(new_n1110));
  INV_X1    g0910(.A(G128), .ZN(new_n1111));
  INV_X1    g0911(.A(G125), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n782), .A2(new_n1111), .B1(new_n771), .B2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(KEYINPUT54), .B(G143), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n787), .A2(new_n994), .B1(new_n789), .B2(new_n1114), .ZN(new_n1115));
  NOR3_X1   g0915(.A1(new_n1110), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n799), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT53), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n775), .B2(new_n335), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n767), .A2(G132), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1106), .A2(new_n1109), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n343), .A2(new_n835), .B1(new_n1121), .B2(new_n756), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n748), .B(new_n1122), .C1(new_n927), .C2(new_n758), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1103), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT120), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n719), .A2(new_n710), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1126), .B(new_n463), .C1(new_n710), .C2(new_n1085), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n656), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n737), .A2(G330), .A3(new_n463), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(KEYINPUT119), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT119), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n932), .A2(new_n1132), .A3(new_n1129), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n734), .A2(new_n736), .A3(G330), .A4(new_n825), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n922), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1137), .A2(new_n1086), .A3(new_n1082), .A4(new_n1076), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1137), .A2(new_n1076), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1138), .B1(new_n1139), .B2(new_n921), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1125), .B1(new_n1134), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1141), .A2(new_n1094), .A3(new_n1101), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1132), .B1(new_n932), .B2(new_n1129), .ZN(new_n1143));
  AND4_X1   g0943(.A1(new_n1132), .A2(new_n1127), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1140), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1147), .A2(new_n1102), .A3(new_n1125), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1142), .A2(new_n1148), .A3(new_n704), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1124), .A2(new_n1149), .ZN(G378));
  NAND2_X1  g0950(.A1(new_n345), .A2(new_n875), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n368), .B(new_n1151), .ZN(new_n1152));
  XOR2_X1   g0952(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1153));
  XOR2_X1   g0953(.A(new_n1152), .B(new_n1153), .Z(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n931), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n929), .B1(new_n1078), .B2(new_n926), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1157), .A2(new_n923), .A3(new_n924), .A4(new_n1154), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n917), .A2(G330), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1156), .A2(new_n1160), .A3(new_n1158), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n980), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1154), .A2(new_n758), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n304), .B(new_n283), .C1(new_n784), .C2(new_n772), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n782), .A2(new_n1112), .B1(new_n789), .B2(new_n994), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n775), .A2(new_n1114), .B1(new_n787), .B2(new_n843), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1168), .B(new_n1169), .C1(G150), .C2(new_n793), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n1111), .B2(new_n766), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1171), .A2(KEYINPUT59), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1167), .B(new_n1172), .C1(G124), .C2(new_n800), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n1171), .A2(KEYINPUT59), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n1006), .A2(new_n789), .B1(new_n529), .B2(new_n766), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n783), .A2(G116), .B1(new_n785), .B2(G58), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G97), .A2(new_n788), .B1(new_n800), .B2(G283), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n299), .A2(new_n283), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n799), .B2(G77), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1177), .A2(new_n1178), .A3(new_n1180), .A4(new_n997), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1176), .A2(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1173), .A2(new_n1174), .B1(new_n1175), .B2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1179), .B(new_n332), .C1(G33), .C2(G41), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n1182), .B2(new_n1175), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT122), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n756), .B1(new_n1183), .B2(new_n1186), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n743), .B(new_n1187), .C1(new_n332), .C2(new_n836), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1166), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1165), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1094), .A2(new_n1101), .A3(new_n1146), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n1145), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1156), .A2(new_n1160), .A3(new_n1158), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1160), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(KEYINPUT57), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT57), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1192), .B(new_n1197), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1190), .B1(new_n1199), .B2(new_n704), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(G375));
  NAND2_X1  g1001(.A1(new_n1146), .A2(new_n980), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G107), .A2(new_n790), .B1(new_n800), .B2(G303), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n488), .B2(new_n775), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n782), .A2(new_n805), .B1(new_n787), .B2(new_n490), .ZN(new_n1205));
  NOR4_X1   g1005(.A1(new_n1204), .A2(new_n350), .A3(new_n1205), .A4(new_n993), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n767), .A2(G283), .B1(new_n392), .B2(new_n793), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n799), .A2(G159), .B1(new_n800), .B2(G128), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n335), .B2(new_n789), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n767), .B2(G137), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n350), .B1(new_n784), .B2(new_n341), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n782), .A2(new_n843), .B1(new_n787), .B2(new_n1114), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(G50), .C2(new_n793), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1206), .A2(new_n1207), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n749), .B1(G68), .B2(new_n835), .C1(new_n756), .C2(new_n1214), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT123), .Z(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n922), .B2(new_n759), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1202), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n964), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1140), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1147), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1219), .A2(new_n1222), .ZN(G381));
  NOR2_X1   g1023(.A1(G375), .A2(G378), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n981), .A2(new_n1054), .A3(new_n1008), .A4(new_n1074), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1013), .A2(new_n1041), .A3(new_n813), .ZN(new_n1226));
  NOR4_X1   g1026(.A1(new_n1225), .A2(G384), .A3(G381), .A4(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1224), .A2(new_n1227), .ZN(G407));
  INV_X1    g1028(.A(G213), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(G343), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1224), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(G407), .A2(new_n1231), .A3(G213), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT124), .ZN(G409));
  INV_X1    g1033(.A(new_n1230), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n704), .B1(new_n1134), .B2(new_n1140), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1221), .A2(KEYINPUT60), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT60), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1134), .A2(new_n1237), .A3(new_n1140), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1235), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(G384), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1239), .A2(new_n1240), .A3(new_n1218), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n705), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1221), .A2(KEYINPUT60), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1237), .B1(new_n1134), .B2(new_n1140), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1242), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(G384), .B1(new_n1245), .B2(new_n1219), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1241), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n705), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1124), .A2(new_n1149), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1248), .A2(new_n1249), .A3(new_n1190), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1164), .A2(new_n980), .B1(new_n1166), .B2(new_n1188), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1164), .A2(new_n1220), .A3(new_n1192), .ZN(new_n1252));
  AOI21_X1  g1052(.A(G378), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1234), .B(new_n1247), .C1(new_n1250), .C2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT63), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(G387), .A2(G390), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G393), .A2(G396), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1226), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1257), .A2(new_n1259), .A3(new_n1225), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1259), .B1(new_n1257), .B2(new_n1225), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1198), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1197), .B1(new_n1164), .B2(new_n1192), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n704), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(G378), .A3(new_n1251), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1253), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1268), .A2(KEYINPUT63), .A3(new_n1234), .A4(new_n1247), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT125), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1240), .B1(new_n1239), .B2(new_n1218), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1245), .A2(G384), .A3(new_n1219), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1230), .A2(G2897), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1271), .A2(new_n1272), .A3(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1274), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1270), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1273), .B1(new_n1241), .B2(new_n1246), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1271), .A2(new_n1272), .A3(new_n1274), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(KEYINPUT125), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1277), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1253), .B1(new_n1200), .B2(G378), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1281), .B1(new_n1282), .B2(new_n1230), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1256), .A2(new_n1262), .A3(new_n1269), .A4(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1262), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT126), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1284), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT127), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1291), .A2(KEYINPUT62), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1254), .A2(new_n1291), .A3(KEYINPUT62), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1291), .A2(KEYINPUT62), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1268), .A2(new_n1234), .A3(new_n1247), .A4(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1292), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1282), .A2(new_n1230), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1298));
  OAI22_X1  g1098(.A1(new_n1297), .A2(new_n1298), .B1(new_n1286), .B2(new_n1289), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1285), .B1(new_n1296), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1290), .A2(new_n1300), .ZN(G405));
  NAND2_X1  g1101(.A1(new_n1262), .A2(new_n1247), .ZN(new_n1302));
  OAI22_X1  g1102(.A1(new_n1260), .A2(new_n1261), .B1(new_n1246), .B2(new_n1241), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(new_n1200), .B(G378), .ZN(new_n1305));
  XOR2_X1   g1105(.A(new_n1304), .B(new_n1305), .Z(G402));
endmodule


