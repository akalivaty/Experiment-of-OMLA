//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT90), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT88), .ZN(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n204), .B1(new_n205), .B2(G1gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G8gat), .ZN(new_n208));
  INV_X1    g007(.A(G1gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT16), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n207), .A2(new_n208), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n211), .ZN(new_n213));
  OAI21_X1  g012(.A(G8gat), .B1(new_n213), .B2(new_n206), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT89), .ZN(new_n215));
  INV_X1    g014(.A(G29gat), .ZN(new_n216));
  INV_X1    g015(.A(G36gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT14), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT14), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(G29gat), .B2(G36gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G43gat), .ZN(new_n223));
  INV_X1    g022(.A(G50gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G43gat), .A2(G50gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT15), .ZN(new_n228));
  NAND2_X1  g027(.A1(G29gat), .A2(G36gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT87), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT15), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n225), .A2(new_n231), .A3(new_n226), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n222), .A2(new_n228), .A3(new_n230), .A4(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234));
  INV_X1    g033(.A(new_n229), .ZN(new_n235));
  OAI211_X1 g034(.A(KEYINPUT15), .B(new_n227), .C1(new_n221), .C2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n233), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n234), .B1(new_n233), .B2(new_n236), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n215), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT89), .B1(new_n212), .B2(new_n214), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n203), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n239), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n237), .ZN(new_n244));
  INV_X1    g043(.A(new_n241), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT90), .A4(new_n215), .ZN(new_n246));
  NAND2_X1  g045(.A1(G229gat), .A2(G233gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n212), .A2(new_n214), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n236), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n242), .A2(new_n246), .A3(new_n247), .A4(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT18), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n202), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G113gat), .B(G141gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(G197gat), .ZN(new_n255));
  XOR2_X1   g054(.A(KEYINPUT11), .B(G169gat), .Z(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT12), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n248), .B(new_n249), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n247), .B(KEYINPUT13), .Z(new_n261));
  AOI22_X1  g060(.A1(new_n251), .A2(new_n252), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n244), .A2(new_n245), .A3(new_n215), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n263), .A2(new_n203), .B1(new_n248), .B2(new_n249), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n264), .A2(KEYINPUT18), .A3(new_n247), .A4(new_n246), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n262), .B(new_n265), .C1(new_n253), .C2(new_n258), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT80), .ZN(new_n270));
  XNOR2_X1  g069(.A(G141gat), .B(G148gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT2), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n272), .B1(G155gat), .B2(G162gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n270), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G155gat), .B(G162gat), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n274), .B(new_n275), .Z(new_n276));
  INV_X1    g075(.A(KEYINPUT3), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT81), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n276), .A2(KEYINPUT81), .A3(new_n277), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT29), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G197gat), .B(G204gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT78), .B(G218gat), .ZN(new_n286));
  INV_X1    g085(.A(G211gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n285), .B1(new_n288), .B2(KEYINPUT22), .ZN(new_n289));
  XNOR2_X1  g088(.A(G211gat), .B(G218gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n284), .A2(KEYINPUT84), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT84), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT29), .B1(new_n280), .B2(new_n281), .ZN(new_n294));
  INV_X1    g093(.A(new_n291), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n277), .B1(new_n291), .B2(KEYINPUT29), .ZN(new_n297));
  INV_X1    g096(.A(new_n276), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n299), .A2(KEYINPUT83), .ZN(new_n300));
  NAND2_X1  g099(.A1(G228gat), .A2(G233gat), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n301), .B1(new_n299), .B2(KEYINPUT83), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n292), .A2(new_n296), .A3(new_n300), .A4(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G22gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n291), .A2(KEYINPUT82), .ZN(new_n305));
  INV_X1    g104(.A(new_n290), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n305), .B(new_n283), .C1(KEYINPUT82), .C2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n276), .B1(new_n308), .B2(new_n277), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n294), .A2(new_n295), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n301), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n303), .A2(new_n304), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n304), .B1(new_n303), .B2(new_n311), .ZN(new_n314));
  OAI21_X1  g113(.A(G78gat), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n303), .A2(new_n311), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G22gat), .ZN(new_n317));
  INV_X1    g116(.A(G78gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n318), .A3(new_n312), .ZN(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT31), .B(G50gat), .ZN(new_n320));
  INV_X1    g119(.A(G106gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n315), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n322), .B1(new_n315), .B2(new_n319), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT25), .ZN(new_n326));
  NAND2_X1  g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT68), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G169gat), .ZN(new_n330));
  INV_X1    g129(.A(G176gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT23), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT69), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G183gat), .A2(G190gat), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT70), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT24), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(new_n337), .B2(new_n336), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT24), .ZN(new_n340));
  INV_X1    g139(.A(G183gat), .ZN(new_n341));
  INV_X1    g140(.A(G190gat), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n342), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n344), .A2(KEYINPUT71), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(KEYINPUT71), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n343), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g146(.A1(G169gat), .A2(G176gat), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n348), .A2(KEYINPUT23), .ZN(new_n349));
  OR2_X1    g148(.A1(new_n349), .A2(KEYINPUT67), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(KEYINPUT67), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n339), .A2(new_n347), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n326), .B1(new_n335), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n343), .A2(KEYINPUT65), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n343), .A2(KEYINPUT65), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n340), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n355), .A2(new_n344), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n350), .A2(new_n351), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT66), .B(G176gat), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(KEYINPUT23), .A3(new_n330), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n329), .A2(new_n326), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n358), .A2(new_n359), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n348), .B(KEYINPUT26), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n329), .ZN(new_n365));
  XOR2_X1   g164(.A(KEYINPUT27), .B(G183gat), .Z(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT72), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n341), .A2(KEYINPUT27), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT72), .ZN(new_n369));
  AOI21_X1  g168(.A(G190gat), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT28), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT28), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n366), .A2(new_n372), .A3(G190gat), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n336), .B(new_n365), .C1(new_n371), .C2(new_n373), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n363), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(G127gat), .B(G134gat), .Z(new_n376));
  XNOR2_X1  g175(.A(G113gat), .B(G120gat), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n376), .B1(KEYINPUT1), .B2(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(new_n378), .B(KEYINPUT73), .Z(new_n379));
  INV_X1    g178(.A(KEYINPUT74), .ZN(new_n380));
  INV_X1    g179(.A(G113gat), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n380), .B1(new_n381), .B2(G120gat), .ZN(new_n382));
  INV_X1    g181(.A(G120gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(KEYINPUT74), .A3(G113gat), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n382), .B(new_n384), .C1(G113gat), .C2(new_n383), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT75), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n376), .A2(KEYINPUT1), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n379), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n354), .A2(new_n375), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n363), .A2(new_n374), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n379), .B(new_n389), .C1(new_n353), .C2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT64), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n391), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT33), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT76), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT76), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n396), .A2(new_n400), .A3(new_n397), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n396), .A2(KEYINPUT32), .ZN(new_n403));
  XNOR2_X1  g202(.A(G15gat), .B(G43gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(KEYINPUT77), .ZN(new_n405));
  XNOR2_X1  g204(.A(G71gat), .B(G99gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n402), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n409));
  INV_X1    g208(.A(new_n395), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OR2_X1    g210(.A1(new_n411), .A2(KEYINPUT34), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(KEYINPUT34), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n407), .A2(KEYINPUT33), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n396), .A2(KEYINPUT32), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n408), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n407), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n419), .B1(new_n401), .B2(new_n399), .ZN(new_n420));
  INV_X1    g219(.A(new_n417), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n414), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n324), .A2(new_n325), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT35), .ZN(new_n425));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(G64gat), .B(G92gat), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  OAI21_X1  g227(.A(new_n283), .B1(new_n353), .B2(new_n392), .ZN(new_n429));
  NAND2_X1  g228(.A1(G226gat), .A2(G233gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g230(.A(G226gat), .B(G233gat), .C1(new_n353), .C2(new_n392), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n295), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(new_n295), .A3(new_n432), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n428), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(new_n428), .A3(new_n435), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n436), .B1(new_n438), .B2(KEYINPUT30), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT30), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT79), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT79), .B1(new_n437), .B2(new_n440), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n439), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G1gat), .B(G29gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT0), .ZN(new_n448));
  XNOR2_X1  g247(.A(G57gat), .B(G85gat), .ZN(new_n449));
  XOR2_X1   g248(.A(new_n448), .B(new_n449), .Z(new_n450));
  OAI211_X1 g249(.A(new_n282), .B(new_n390), .C1(new_n277), .C2(new_n276), .ZN(new_n451));
  NAND2_X1  g250(.A1(G225gat), .A2(G233gat), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n379), .A2(new_n276), .A3(new_n389), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n453), .B(KEYINPUT4), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n390), .A2(new_n298), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n453), .ZN(new_n457));
  INV_X1    g256(.A(new_n452), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT5), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT5), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n455), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n450), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n455), .A2(new_n463), .ZN(new_n466));
  INV_X1    g265(.A(new_n450), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n467), .A3(new_n461), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT6), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n465), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n466), .A2(new_n461), .A3(KEYINPUT6), .A4(new_n467), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n446), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n424), .A2(new_n425), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n315), .A2(new_n319), .ZN(new_n476));
  INV_X1    g275(.A(new_n322), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n423), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n479), .A3(new_n323), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT35), .B1(new_n480), .B2(new_n473), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n452), .B1(new_n451), .B2(new_n454), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT39), .B1(new_n457), .B2(new_n458), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n450), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI211_X1 g284(.A(KEYINPUT39), .B(new_n452), .C1(new_n451), .C2(new_n454), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT40), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n488), .A2(new_n468), .ZN(new_n489));
  XOR2_X1   g288(.A(KEYINPUT85), .B(KEYINPUT40), .Z(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(new_n485), .B2(new_n486), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT86), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT86), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n493), .B(new_n490), .C1(new_n485), .C2(new_n486), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n489), .A2(new_n445), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n435), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT37), .B1(new_n497), .B2(new_n433), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT37), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n434), .A2(new_n499), .A3(new_n435), .ZN(new_n500));
  INV_X1    g299(.A(new_n428), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n438), .B1(new_n502), .B2(KEYINPUT38), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT38), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n498), .A2(new_n500), .A3(new_n504), .A4(new_n501), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n470), .A2(new_n503), .A3(new_n471), .A4(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n496), .A2(new_n478), .A3(new_n506), .A4(new_n323), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n470), .A2(new_n471), .ZN(new_n508));
  OAI22_X1  g307(.A1(new_n324), .A2(new_n325), .B1(new_n508), .B2(new_n445), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n418), .A2(KEYINPUT36), .A3(new_n422), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT36), .B1(new_n418), .B2(new_n422), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n507), .B(new_n509), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n269), .B1(new_n482), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G85gat), .A2(G92gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT7), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT7), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(G85gat), .A3(G92gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G99gat), .A2(G106gat), .ZN(new_n520));
  INV_X1    g319(.A(G85gat), .ZN(new_n521));
  INV_X1    g320(.A(G92gat), .ZN(new_n522));
  AOI22_X1  g321(.A1(KEYINPUT8), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G99gat), .B(G106gat), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n519), .A2(new_n523), .A3(new_n525), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n244), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n528), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n525), .B1(new_n519), .B2(new_n523), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G232gat), .A2(G233gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT96), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n249), .A2(new_n533), .B1(KEYINPUT41), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n530), .A2(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(G190gat), .B(G218gat), .Z(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n536), .A2(KEYINPUT41), .ZN(new_n541));
  XNOR2_X1  g340(.A(G134gat), .B(G162gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n540), .B(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G71gat), .B(G78gat), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n548));
  INV_X1    g347(.A(G57gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(G64gat), .ZN(new_n550));
  INV_X1    g349(.A(G64gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(G57gat), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n548), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  OAI211_X1 g352(.A(KEYINPUT93), .B(new_n547), .C1(new_n553), .C2(KEYINPUT92), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT93), .ZN(new_n555));
  NAND2_X1  g354(.A1(G71gat), .A2(G78gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n551), .A2(G57gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n549), .A2(G64gat), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT92), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n555), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n546), .B1(new_n553), .B2(KEYINPUT93), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n554), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n533), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT10), .ZN(new_n567));
  XNOR2_X1  g366(.A(G57gat), .B(G64gat), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n555), .B1(new_n568), .B2(new_n548), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n550), .A2(new_n552), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT92), .B1(new_n570), .B2(new_n558), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n546), .B(new_n569), .C1(new_n571), .C2(new_n555), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n529), .A2(new_n572), .A3(new_n554), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n566), .A2(new_n567), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n565), .A2(new_n533), .A3(KEYINPUT10), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n574), .A2(KEYINPUT97), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT97), .B1(new_n574), .B2(new_n575), .ZN(new_n577));
  AND2_X1   g376(.A1(G230gat), .A2(G233gat), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n566), .A2(new_n573), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n578), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT98), .ZN(new_n582));
  XNOR2_X1  g381(.A(G120gat), .B(G148gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(G176gat), .B(G204gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NOR3_X1   g385(.A1(new_n579), .A2(new_n582), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT100), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n575), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n578), .B(KEYINPUT99), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n589), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  AOI211_X1 g392(.A(KEYINPUT100), .B(new_n591), .C1(new_n574), .C2(new_n575), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n586), .B1(new_n595), .B2(new_n582), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n588), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G127gat), .B(G155gat), .ZN(new_n598));
  INV_X1    g397(.A(new_n565), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT21), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n603), .A2(new_n604), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n598), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n607), .ZN(new_n609));
  INV_X1    g408(.A(new_n598), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(new_n610), .A3(new_n605), .ZN(new_n611));
  XOR2_X1   g410(.A(G183gat), .B(G211gat), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n608), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n613), .B1(new_n608), .B2(new_n611), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n214), .B(new_n212), .C1(new_n599), .C2(new_n600), .ZN(new_n617));
  XNOR2_X1  g416(.A(KEYINPUT95), .B(KEYINPUT20), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n615), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n619), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n608), .A2(new_n611), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n612), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n621), .B1(new_n623), .B2(new_n614), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n545), .B(new_n597), .C1(new_n620), .C2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n514), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(new_n472), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(new_n209), .ZN(G1324gat));
  XNOR2_X1  g428(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n630));
  INV_X1    g429(.A(new_n627), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n445), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT16), .B(G8gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT102), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n630), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(G8gat), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT42), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n635), .B(new_n636), .C1(new_n632), .C2(new_n638), .ZN(G1325gat));
  AOI21_X1  g438(.A(G15gat), .B1(new_n631), .B2(new_n479), .ZN(new_n640));
  OAI21_X1  g439(.A(KEYINPUT103), .B1(new_n511), .B2(new_n512), .ZN(new_n641));
  INV_X1    g440(.A(new_n512), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT103), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(new_n510), .A3(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(G15gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT104), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n640), .B1(new_n631), .B2(new_n648), .ZN(G1326gat));
  NOR2_X1   g448(.A1(new_n324), .A2(new_n325), .ZN(new_n650));
  OR3_X1    g449(.A1(new_n627), .A2(KEYINPUT105), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT105), .B1(new_n627), .B2(new_n650), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT43), .B(G22gat), .ZN(new_n653));
  AND3_X1   g452(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n653), .B1(new_n651), .B2(new_n652), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n654), .A2(new_n655), .ZN(G1327gat));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n507), .A2(new_n509), .A3(new_n644), .A4(new_n641), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n425), .B1(new_n424), .B2(new_n474), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n480), .A2(KEYINPUT35), .A3(new_n473), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n544), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n545), .A2(new_n663), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(new_n482), .B2(new_n513), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n620), .A2(new_n624), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n597), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n269), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n664), .A2(new_n668), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n657), .B1(new_n675), .B2(new_n472), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT44), .B1(new_n661), .B2(new_n544), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n677), .A2(new_n667), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n678), .A2(KEYINPUT106), .A3(new_n508), .A4(new_n674), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n676), .A2(G29gat), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n673), .A2(new_n545), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n514), .A2(new_n216), .A3(new_n508), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT45), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(G1328gat));
  AND2_X1   g483(.A1(new_n514), .A2(new_n681), .ZN(new_n685));
  AOI21_X1  g484(.A(G36gat), .B1(KEYINPUT107), .B2(KEYINPUT46), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n445), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(G36gat), .B1(new_n675), .B2(new_n446), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(G1329gat));
  XNOR2_X1  g490(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n646), .A2(G43gat), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n675), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(G43gat), .B1(new_n685), .B2(new_n479), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n693), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n685), .A2(new_n479), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n223), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n699), .B(new_n692), .C1(new_n675), .C2(new_n694), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n700), .ZN(G1330gat));
  INV_X1    g500(.A(new_n650), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(G50gat), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n675), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(G50gat), .B1(new_n685), .B2(new_n702), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT48), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n685), .A2(new_n702), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n224), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT48), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n708), .B(new_n709), .C1(new_n675), .C2(new_n703), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n706), .A2(new_n710), .ZN(G1331gat));
  OAI21_X1  g510(.A(new_n619), .B1(new_n615), .B2(new_n616), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n623), .A2(new_n621), .A3(new_n614), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n544), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n714), .A2(new_n269), .A3(new_n671), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n661), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n472), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(new_n549), .ZN(G1332gat));
  AND2_X1   g517(.A1(new_n661), .A2(new_n715), .ZN(new_n719));
  NOR2_X1   g518(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n720));
  AND2_X1   g519(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n719), .B(new_n445), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT109), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n716), .A2(new_n446), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n722), .B(new_n723), .C1(new_n724), .C2(new_n720), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n724), .A2(new_n720), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n723), .B1(new_n727), .B2(new_n722), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n726), .A2(new_n728), .ZN(G1333gat));
  XNOR2_X1  g528(.A(new_n423), .B(KEYINPUT110), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(G71gat), .B1(new_n719), .B2(new_n731), .ZN(new_n732));
  AND4_X1   g531(.A1(G71gat), .A2(new_n661), .A3(new_n646), .A4(new_n715), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1334gat));
  NOR2_X1   g535(.A1(new_n716), .A2(new_n650), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(new_n318), .ZN(G1335gat));
  NAND3_X1  g537(.A1(new_n508), .A2(new_n521), .A3(new_n671), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT112), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n267), .A2(new_n268), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n670), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n661), .A2(new_n544), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n661), .A2(KEYINPUT51), .A3(new_n544), .A4(new_n742), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n745), .A2(KEYINPUT111), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT111), .B1(new_n745), .B2(new_n746), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n740), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n742), .A2(new_n671), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n664), .A2(new_n668), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752), .B2(new_n472), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n749), .A2(new_n753), .ZN(G1336gat));
  NOR3_X1   g553(.A1(new_n677), .A2(new_n667), .A3(new_n750), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n522), .B1(new_n755), .B2(new_n445), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n446), .A2(G92gat), .A3(new_n597), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n758), .B1(new_n745), .B2(new_n746), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT52), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(G92gat), .B1(new_n752), .B2(new_n446), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762));
  INV_X1    g561(.A(new_n759), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n760), .A2(new_n764), .ZN(G1337gat));
  NOR3_X1   g564(.A1(new_n423), .A2(G99gat), .A3(new_n597), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n747), .B2(new_n748), .ZN(new_n767));
  OAI21_X1  g566(.A(G99gat), .B1(new_n752), .B2(new_n645), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(G1338gat));
  AOI21_X1  g568(.A(new_n321), .B1(new_n755), .B2(new_n702), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n597), .A2(G106gat), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n702), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n745), .B2(new_n746), .ZN(new_n773));
  OAI21_X1  g572(.A(KEYINPUT53), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(G106gat), .B1(new_n752), .B2(new_n650), .ZN(new_n775));
  INV_X1    g574(.A(new_n773), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n774), .A2(new_n778), .ZN(G1339gat));
  NAND3_X1  g578(.A1(new_n574), .A2(new_n575), .A3(new_n591), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT54), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT114), .B1(new_n579), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT97), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n578), .B1(new_n590), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n574), .A2(KEYINPUT97), .A3(new_n575), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n787));
  INV_X1    g586(.A(new_n781), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n782), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n593), .B2(new_n594), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n586), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n792), .A2(KEYINPUT55), .A3(new_n586), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n790), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n588), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n587), .B1(new_n790), .B2(new_n799), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT115), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n798), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n247), .B1(new_n264), .B2(new_n246), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n260), .A2(new_n261), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n257), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n258), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n809), .B1(new_n266), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n545), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n806), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n804), .A2(KEYINPUT115), .ZN(new_n814));
  AOI211_X1 g613(.A(new_n802), .B(new_n587), .C1(new_n790), .C2(new_n799), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n741), .B(new_n797), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n597), .A2(new_n811), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n544), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n669), .B1(new_n813), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n821), .B1(new_n625), .B2(new_n741), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n714), .A2(KEYINPUT113), .A3(new_n269), .A4(new_n597), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n472), .A2(new_n445), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n825), .A2(new_n424), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n741), .ZN(new_n828));
  XNOR2_X1  g627(.A(KEYINPUT116), .B(G113gat), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n828), .B(new_n829), .ZN(G1340gat));
  NAND2_X1  g629(.A1(new_n827), .A2(new_n671), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g631(.A1(new_n827), .A2(new_n670), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g633(.A1(new_n827), .A2(new_n544), .ZN(new_n835));
  OR3_X1    g634(.A1(new_n835), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT56), .B1(new_n835), .B2(G134gat), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(G134gat), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(G1343gat));
  INV_X1    g638(.A(KEYINPUT58), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n641), .A2(new_n644), .A3(new_n826), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n269), .A2(G141gat), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n825), .A2(new_n841), .A3(new_n702), .A4(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n840), .B1(new_n843), .B2(KEYINPUT119), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n844), .B1(KEYINPUT119), .B2(new_n843), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT57), .B1(new_n825), .B2(new_n702), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n650), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n793), .B1(new_n782), .B2(new_n789), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n800), .B(new_n588), .C1(new_n850), .C2(KEYINPUT55), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n797), .A2(KEYINPUT117), .A3(new_n804), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n854), .A3(new_n741), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n544), .B1(new_n855), .B2(new_n818), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n669), .B1(new_n856), .B2(new_n813), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n849), .B1(new_n857), .B2(new_n824), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n741), .B(new_n841), .C1(new_n846), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(G141gat), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n843), .B(KEYINPUT118), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n862), .B1(G141gat), .B2(new_n859), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n863), .B2(new_n840), .ZN(G1344gat));
  NOR2_X1   g663(.A1(new_n625), .A2(new_n741), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n650), .B1(new_n857), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n806), .A2(new_n812), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n817), .B1(new_n806), .B2(new_n741), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n868), .B1(new_n869), .B2(new_n544), .ZN(new_n870));
  AOI22_X1  g669(.A1(new_n870), .A2(new_n669), .B1(new_n822), .B2(new_n823), .ZN(new_n871));
  OAI22_X1  g670(.A1(new_n867), .A2(KEYINPUT57), .B1(new_n871), .B2(new_n849), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n872), .A2(new_n671), .A3(new_n841), .ZN(new_n873));
  INV_X1    g672(.A(G148gat), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT59), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n671), .B(new_n841), .C1(new_n846), .C2(new_n858), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n874), .A2(KEYINPUT59), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n876), .A2(new_n878), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT121), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n875), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n825), .A2(new_n702), .A3(new_n841), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n883), .A2(G148gat), .A3(new_n597), .ZN(new_n884));
  XOR2_X1   g683(.A(new_n884), .B(KEYINPUT120), .Z(new_n885));
  NAND2_X1  g684(.A1(new_n882), .A2(new_n885), .ZN(G1345gat));
  OAI21_X1  g685(.A(new_n841), .B1(new_n846), .B2(new_n858), .ZN(new_n887));
  OAI21_X1  g686(.A(G155gat), .B1(new_n887), .B2(new_n669), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n669), .A2(G155gat), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n883), .B2(new_n889), .ZN(G1346gat));
  OAI21_X1  g689(.A(KEYINPUT122), .B1(new_n887), .B2(new_n545), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G162gat), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n887), .A2(KEYINPUT122), .A3(new_n545), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n545), .A2(G162gat), .ZN(new_n894));
  OAI22_X1  g693(.A1(new_n892), .A2(new_n893), .B1(new_n883), .B2(new_n894), .ZN(G1347gat));
  NAND2_X1  g694(.A1(new_n472), .A2(new_n445), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n702), .A2(new_n730), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n825), .A2(new_n897), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n898), .A2(new_n330), .A3(new_n269), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n480), .A2(new_n446), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n825), .A2(new_n472), .A3(new_n900), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT123), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n741), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n899), .B1(new_n903), .B2(new_n330), .ZN(G1348gat));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n905));
  AOI21_X1  g704(.A(G176gat), .B1(new_n902), .B2(new_n671), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n898), .A2(new_n360), .A3(new_n597), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n901), .B(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n331), .B1(new_n910), .B2(new_n597), .ZN(new_n911));
  INV_X1    g710(.A(new_n907), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(KEYINPUT124), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n908), .A2(new_n913), .ZN(G1349gat));
  OR3_X1    g713(.A1(new_n901), .A2(new_n366), .A3(new_n669), .ZN(new_n915));
  OAI21_X1  g714(.A(G183gat), .B1(new_n898), .B2(new_n669), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n915), .A2(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n919), .B(new_n920), .ZN(G1350gat));
  NAND3_X1  g720(.A1(new_n902), .A2(new_n342), .A3(new_n544), .ZN(new_n922));
  OAI21_X1  g721(.A(G190gat), .B1(new_n898), .B2(new_n545), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT61), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1351gat));
  NOR3_X1   g724(.A1(new_n646), .A2(new_n650), .A3(new_n446), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n926), .A2(new_n472), .A3(new_n825), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n269), .A2(G197gat), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n645), .A2(new_n472), .A3(new_n445), .A4(new_n741), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n269), .B1(new_n851), .B2(new_n852), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n817), .B1(new_n931), .B2(new_n854), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n868), .B1(new_n932), .B2(new_n544), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n865), .B1(new_n933), .B2(new_n669), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n847), .B1(new_n934), .B2(new_n650), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n825), .A2(new_n848), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n930), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT126), .ZN(new_n938));
  OAI21_X1  g737(.A(G197gat), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI211_X1 g738(.A(KEYINPUT126), .B(new_n930), .C1(new_n935), .C2(new_n936), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n929), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI211_X1 g742(.A(KEYINPUT127), .B(new_n929), .C1(new_n939), .C2(new_n940), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1352gat));
  NOR2_X1   g744(.A1(new_n597), .A2(G204gat), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n926), .A2(new_n472), .A3(new_n825), .A4(new_n946), .ZN(new_n947));
  XOR2_X1   g746(.A(new_n947), .B(KEYINPUT62), .Z(new_n948));
  NOR2_X1   g747(.A1(new_n646), .A2(new_n896), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n872), .A2(new_n671), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G204gat), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n948), .A2(new_n951), .ZN(G1353gat));
  NAND3_X1  g751(.A1(new_n927), .A2(new_n287), .A3(new_n670), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n872), .A2(new_n949), .A3(new_n670), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n954), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT63), .B1(new_n954), .B2(G211gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(G1354gat));
  AOI21_X1  g756(.A(G218gat), .B1(new_n927), .B2(new_n544), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n872), .A2(new_n949), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n545), .A2(new_n286), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(G1355gat));
endmodule


