//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n547,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n555,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n587,
    new_n588, new_n589, new_n590, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n633, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g023(.A(G2106), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT66), .Z(new_n453));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n455), .A2(new_n449), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G101), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n470), .B1(new_n471), .B2(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n464), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT69), .B1(new_n468), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n472), .A2(new_n473), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n477), .A2(new_n478), .A3(new_n467), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n465), .A2(new_n466), .ZN(new_n481));
  INV_X1    g056(.A(G125), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n475), .A2(new_n479), .B1(G2105), .B2(new_n483), .ZN(G160));
  OR2_X1    g059(.A1(new_n465), .A2(new_n466), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n485), .A2(KEYINPUT70), .A3(new_n464), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n487), .B1(new_n481), .B2(G2105), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G112), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n481), .A2(new_n464), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G124), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G162));
  OAI211_X1 g072(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n464), .A2(G114), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g076(.A(G138), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n502));
  OR2_X1    g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(G164));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT71), .B1(new_n506), .B2(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(new_n509), .A3(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n511), .A2(G50), .A3(G543), .A4(new_n512), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n513), .A2(KEYINPUT72), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(KEYINPUT72), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT73), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n522), .A2(new_n506), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT75), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n516), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n511), .A2(new_n521), .A3(new_n512), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT74), .B(G88), .Z(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n530), .B1(new_n523), .B2(new_n524), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n526), .A2(new_n531), .ZN(G166));
  NAND3_X1  g107(.A1(new_n511), .A2(G543), .A3(new_n512), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n507), .A2(new_n510), .B1(KEYINPUT6), .B2(new_n506), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n536), .A2(KEYINPUT76), .A3(G543), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n538), .A2(G51), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n541), .A2(KEYINPUT7), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(KEYINPUT7), .ZN(new_n543));
  INV_X1    g118(.A(G89), .ZN(new_n544));
  OAI221_X1 g119(.A(new_n540), .B1(new_n542), .B2(new_n543), .C1(new_n527), .C2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n539), .A2(new_n545), .ZN(G168));
  AOI22_X1  g121(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n506), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n549), .B2(new_n527), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n550), .B1(G52), .B2(new_n538), .ZN(G171));
  AOI22_X1  g126(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n552), .A2(new_n506), .B1(new_n527), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n554), .B1(G43), .B2(new_n538), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  INV_X1    g135(.A(KEYINPUT80), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n511), .A2(G53), .A3(G543), .A4(new_n512), .ZN(new_n562));
  NAND2_X1  g137(.A1(KEYINPUT77), .A2(KEYINPUT9), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n536), .A2(G91), .A3(new_n521), .ZN(new_n565));
  AND3_X1   g140(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n566));
  AOI21_X1  g141(.A(KEYINPUT5), .B1(KEYINPUT73), .B2(G543), .ZN(new_n567));
  OAI21_X1  g142(.A(G65), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT78), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n571), .A2(G78), .A3(G543), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n568), .A2(KEYINPUT79), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G651), .ZN(new_n575));
  AOI21_X1  g150(.A(KEYINPUT79), .B1(new_n568), .B2(new_n573), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n565), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n561), .B1(new_n564), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n562), .A2(KEYINPUT77), .A3(KEYINPUT9), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n536), .A2(G53), .A3(G543), .A4(new_n563), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n576), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n582), .A2(G651), .A3(new_n574), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n581), .A2(new_n583), .A3(KEYINPUT80), .A4(new_n565), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G299));
  AND4_X1   g161(.A1(KEYINPUT76), .A2(new_n511), .A3(G543), .A4(new_n512), .ZN(new_n587));
  AOI21_X1  g162(.A(KEYINPUT76), .B1(new_n536), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(G52), .ZN(new_n590));
  OAI221_X1 g165(.A(new_n548), .B1(new_n549), .B2(new_n527), .C1(new_n589), .C2(new_n590), .ZN(G301));
  INV_X1    g166(.A(G168), .ZN(G286));
  INV_X1    g167(.A(G166), .ZN(G303));
  NAND3_X1  g168(.A1(new_n536), .A2(G87), .A3(new_n521), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n536), .A2(G49), .A3(G543), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT81), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n566), .A2(new_n567), .ZN(new_n599));
  INV_X1    g174(.A(G74), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(KEYINPUT81), .B1(new_n601), .B2(G651), .ZN(new_n602));
  OAI211_X1 g177(.A(new_n594), .B(new_n595), .C1(new_n598), .C2(new_n602), .ZN(G288));
  INV_X1    g178(.A(G48), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n533), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(G86), .B2(new_n528), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT82), .ZN(new_n607));
  INV_X1    g182(.A(G61), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(new_n519), .B2(new_n520), .ZN(new_n609));
  AND2_X1   g184(.A1(G73), .A2(G543), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n607), .B1(new_n611), .B2(new_n506), .ZN(new_n612));
  OAI211_X1 g187(.A(KEYINPUT82), .B(G651), .C1(new_n609), .C2(new_n610), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n606), .A2(new_n612), .A3(new_n613), .ZN(G305));
  AOI22_X1  g189(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G85), .ZN(new_n616));
  OAI22_X1  g191(.A1(new_n615), .A2(new_n506), .B1(new_n527), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(G47), .B2(new_n538), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(G290));
  NAND2_X1  g194(.A1(G301), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(G66), .B1(new_n566), .B2(new_n567), .ZN(new_n621));
  NAND2_X1  g196(.A1(G79), .A2(G543), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n506), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND4_X1  g198(.A1(new_n511), .A2(new_n521), .A3(G92), .A4(new_n512), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT10), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g201(.A1(new_n536), .A2(KEYINPUT10), .A3(G92), .A4(new_n521), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(G54), .B1(new_n587), .B2(new_n588), .ZN(new_n629));
  AND2_X1   g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n620), .B1(G868), .B2(new_n630), .ZN(G284));
  OAI21_X1  g206(.A(new_n620), .B1(G868), .B2(new_n630), .ZN(G321));
  NAND2_X1  g207(.A1(G286), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n585), .ZN(G297));
  XNOR2_X1  g209(.A(G297), .B(KEYINPUT83), .ZN(G280));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n630), .B1(new_n636), .B2(G860), .ZN(G148));
  NAND2_X1  g212(.A1(new_n630), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G868), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n639), .A2(KEYINPUT84), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(KEYINPUT84), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n640), .B(new_n641), .C1(G868), .C2(new_n555), .ZN(G323));
  XNOR2_X1  g217(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g218(.A1(new_n489), .A2(G135), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT85), .Z(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n646));
  INV_X1    g221(.A(G111), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n646), .B1(new_n647), .B2(G2105), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(new_n494), .B2(G123), .ZN(new_n649));
  AND2_X1   g224(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(G2096), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n485), .A2(new_n476), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT12), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT13), .ZN(new_n656));
  INV_X1    g231(.A(G2100), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n652), .A2(new_n653), .A3(new_n658), .ZN(G156));
  XNOR2_X1  g234(.A(G2427), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2430), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT15), .B(G2435), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(KEYINPUT14), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT86), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2451), .B(G2454), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT16), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2443), .B(G2446), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n666), .A2(new_n668), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n666), .A2(new_n668), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n673), .A2(new_n670), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1341), .B(G1348), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n677), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n672), .A2(new_n679), .A3(new_n675), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT87), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  OAI211_X1 g258(.A(G14), .B(new_n678), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT88), .ZN(G401));
  INV_X1    g260(.A(KEYINPUT18), .ZN(new_n686));
  XOR2_X1   g261(.A(G2084), .B(G2090), .Z(new_n687));
  XNOR2_X1  g262(.A(G2067), .B(G2678), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(KEYINPUT17), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n687), .A2(new_n688), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n686), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(new_n657), .ZN(new_n693));
  XOR2_X1   g268(.A(G2072), .B(G2078), .Z(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n689), .B2(KEYINPUT18), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(new_n651), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n693), .B(new_n696), .ZN(G227));
  XNOR2_X1  g272(.A(G1971), .B(G1976), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT19), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(G1956), .B(G2474), .Z(new_n701));
  XOR2_X1   g276(.A(G1961), .B(G1966), .Z(new_n702));
  AND2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT20), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n701), .A2(new_n702), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  MUX2_X1   g283(.A(new_n708), .B(new_n707), .S(new_n700), .Z(new_n709));
  NOR2_X1   g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1991), .B(G1996), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(G1981), .B(G1986), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(G229));
  INV_X1    g291(.A(KEYINPUT95), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n718), .A2(G33), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT25), .Z(new_n721));
  AOI22_X1  g296(.A1(new_n485), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n486), .A2(new_n488), .ZN(new_n723));
  INV_X1    g298(.A(G139), .ZN(new_n724));
  OAI221_X1 g299(.A(new_n721), .B1(new_n722), .B2(new_n464), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n719), .B1(new_n725), .B2(G29), .ZN(new_n726));
  INV_X1    g301(.A(G2072), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n718), .A2(G32), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n494), .A2(G129), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n476), .A2(G105), .ZN(new_n731));
  NAND3_X1  g306(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT26), .Z(new_n733));
  AND3_X1   g308(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G141), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n723), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n729), .B1(new_n736), .B2(G29), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT27), .B(G1996), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n650), .B2(G29), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT31), .B(G11), .Z(new_n741));
  INV_X1    g316(.A(G28), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(KEYINPUT30), .ZN(new_n743));
  AOI21_X1  g318(.A(G29), .B1(new_n742), .B2(KEYINPUT30), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT92), .B(KEYINPUT24), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(G29), .B1(new_n747), .B2(G34), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G34), .B2(new_n747), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G160), .B2(new_n718), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(G2084), .Z(new_n751));
  AND4_X1   g326(.A1(new_n728), .A2(new_n740), .A3(new_n745), .A4(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G2078), .ZN(new_n753));
  NAND2_X1  g328(.A1(G164), .A2(G29), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G27), .B2(G29), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n737), .A2(new_n738), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  OAI221_X1 g331(.A(new_n756), .B1(new_n727), .B2(new_n726), .C1(new_n753), .C2(new_n755), .ZN(new_n757));
  INV_X1    g332(.A(G16), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G21), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G168), .B2(new_n758), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n757), .B1(G1966), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n758), .A2(G5), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G171), .B2(new_n758), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1961), .ZN(new_n764));
  INV_X1    g339(.A(G1966), .ZN(new_n765));
  INV_X1    g340(.A(new_n760), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AND3_X1   g342(.A1(new_n752), .A2(new_n761), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(KEYINPUT93), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n758), .A2(G4), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n630), .B2(new_n758), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1348), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n718), .A2(G26), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT28), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n489), .A2(G140), .ZN(new_n775));
  OAI21_X1  g350(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n776));
  INV_X1    g351(.A(G116), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(G2105), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n494), .B2(G128), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n774), .B1(new_n780), .B2(G29), .ZN(new_n781));
  INV_X1    g356(.A(G2067), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n758), .A2(G19), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n555), .B2(new_n758), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1341), .ZN(new_n786));
  OR3_X1    g361(.A1(new_n772), .A2(new_n783), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(KEYINPUT91), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n769), .A2(new_n788), .ZN(new_n789));
  OAI22_X1  g364(.A1(new_n768), .A2(KEYINPUT93), .B1(KEYINPUT91), .B2(new_n787), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n718), .A2(G35), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G162), .B2(new_n718), .ZN(new_n793));
  INV_X1    g368(.A(G2090), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n758), .A2(G20), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT23), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n585), .B2(new_n758), .ZN(new_n800));
  INV_X1    g375(.A(G1956), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n717), .B1(new_n791), .B2(new_n803), .ZN(new_n804));
  OR4_X1    g379(.A1(new_n717), .A2(new_n789), .A3(new_n790), .A4(new_n803), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n758), .A2(G23), .ZN(new_n806));
  INV_X1    g381(.A(G288), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(new_n758), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT90), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT33), .B(G1976), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n809), .B(new_n810), .Z(new_n811));
  NOR2_X1   g386(.A1(G6), .A2(G16), .ZN(new_n812));
  INV_X1    g387(.A(G86), .ZN(new_n813));
  OAI221_X1 g388(.A(new_n613), .B1(new_n527), .B2(new_n813), .C1(new_n604), .C2(new_n533), .ZN(new_n814));
  INV_X1    g389(.A(new_n612), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n812), .B1(new_n816), .B2(G16), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT32), .B(G1981), .Z(new_n818));
  XOR2_X1   g393(.A(new_n817), .B(new_n818), .Z(new_n819));
  NOR2_X1   g394(.A1(G16), .A2(G22), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G166), .B2(G16), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G1971), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n811), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT34), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n494), .A2(G119), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT89), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n489), .A2(G131), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n464), .A2(G107), .ZN(new_n830));
  OAI21_X1  g405(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n828), .B(new_n829), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  MUX2_X1   g407(.A(G25), .B(new_n832), .S(G29), .Z(new_n833));
  XOR2_X1   g408(.A(KEYINPUT35), .B(G1991), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(G1986), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n618), .A2(new_n758), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n758), .B2(G24), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n835), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(new_n836), .B2(new_n838), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n825), .A2(new_n826), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(KEYINPUT36), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n841), .A2(KEYINPUT36), .ZN(new_n843));
  AOI22_X1  g418(.A1(new_n804), .A2(new_n805), .B1(new_n842), .B2(new_n843), .ZN(G311));
  NAND2_X1  g419(.A1(new_n804), .A2(new_n805), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n841), .B(KEYINPUT36), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(G150));
  NAND2_X1  g422(.A1(new_n630), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n538), .A2(G55), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n521), .A2(G67), .ZN(new_n851));
  AND2_X1   g426(.A1(G80), .A2(G543), .ZN(new_n852));
  OAI21_X1  g427(.A(KEYINPUT96), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n852), .B1(new_n521), .B2(G67), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(G651), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n528), .A2(G93), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n850), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n554), .ZN(new_n860));
  INV_X1    g435(.A(G43), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n589), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n555), .A2(new_n857), .A3(new_n850), .A4(new_n858), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n849), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT97), .ZN(new_n869));
  AOI21_X1  g444(.A(G860), .B1(new_n866), .B2(new_n867), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT98), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n859), .A2(G860), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT37), .Z(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(G145));
  XNOR2_X1  g450(.A(new_n832), .B(new_n655), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n725), .A2(KEYINPUT99), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n736), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n876), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n503), .A2(new_n504), .ZN(new_n880));
  INV_X1    g455(.A(new_n501), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n780), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(G118), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n884), .A2(KEYINPUT100), .A3(G2105), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT100), .B1(new_n884), .B2(G2105), .ZN(new_n886));
  OAI21_X1  g461(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI22_X1  g463(.A1(new_n494), .A2(G130), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(G142), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n889), .B1(new_n723), .B2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n883), .B(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n879), .B(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n496), .B(G160), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n650), .B(new_n894), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(G37), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n893), .A2(new_n895), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g475(.A(new_n865), .B(new_n638), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n630), .B1(new_n578), .B2(new_n584), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n578), .A2(new_n630), .A3(new_n584), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n578), .A2(new_n630), .A3(KEYINPUT101), .A4(new_n584), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n903), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT41), .B1(new_n910), .B2(new_n904), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n906), .A2(new_n907), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n903), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT102), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n912), .A2(KEYINPUT102), .A3(new_n914), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n909), .B1(new_n919), .B2(new_n902), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n816), .B1(new_n526), .B2(new_n531), .ZN(new_n921));
  INV_X1    g496(.A(new_n531), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n514), .A2(new_n515), .B1(new_n523), .B2(new_n524), .ZN(new_n923));
  NAND3_X1  g498(.A1(G305), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(G290), .A2(new_n807), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n618), .A2(G288), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT42), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n921), .A2(new_n924), .A3(new_n926), .A4(new_n927), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n929), .A2(KEYINPUT103), .A3(new_n931), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT103), .B1(new_n929), .B2(new_n931), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n932), .B1(new_n935), .B2(new_n930), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n920), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n936), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n912), .A2(KEYINPUT102), .A3(new_n914), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT102), .B1(new_n912), .B2(new_n914), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n942), .A2(new_n943), .A3(new_n911), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n944), .A2(new_n901), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n940), .B(new_n941), .C1(new_n945), .C2(new_n909), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n920), .A2(KEYINPUT104), .A3(new_n936), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT105), .B1(new_n920), .B2(new_n936), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n939), .A2(new_n946), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(G868), .ZN(new_n950));
  INV_X1    g525(.A(G868), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n859), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(G295));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n954), .B1(new_n950), .B2(new_n952), .ZN(new_n955));
  INV_X1    g530(.A(new_n952), .ZN(new_n956));
  AOI211_X1 g531(.A(KEYINPUT106), .B(new_n956), .C1(new_n949), .C2(G868), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n955), .A2(new_n957), .ZN(G331));
  OR2_X1    g533(.A1(new_n933), .A2(new_n934), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n863), .A2(new_n864), .A3(G301), .ZN(new_n960));
  AOI21_X1  g535(.A(G301), .B1(new_n863), .B2(new_n864), .ZN(new_n961));
  OAI21_X1  g536(.A(G286), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n865), .A2(G171), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n863), .A2(new_n864), .A3(G301), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(G168), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n908), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n959), .B(new_n968), .C1(new_n944), .C2(new_n966), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n897), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n968), .B1(new_n944), .B2(new_n966), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n959), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI211_X1 g548(.A(KEYINPUT107), .B(new_n968), .C1(new_n944), .C2(new_n966), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n970), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n908), .B1(new_n962), .B2(new_n965), .ZN(new_n978));
  INV_X1    g553(.A(new_n966), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n978), .B1(new_n919), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(G37), .B1(new_n980), .B2(new_n959), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n914), .A2(new_n904), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(new_n908), .B2(KEYINPUT41), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n979), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n968), .A2(KEYINPUT108), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n967), .A2(new_n913), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n966), .B1(new_n987), .B2(new_n983), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n985), .B(new_n935), .C1(new_n986), .C2(new_n988), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n981), .A2(new_n989), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n977), .B(KEYINPUT44), .C1(new_n976), .C2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n981), .A2(new_n976), .A3(new_n989), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(new_n975), .B2(new_n976), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT109), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n966), .B1(new_n917), .B2(new_n918), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n972), .B1(new_n996), .B2(new_n978), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n997), .A2(new_n974), .A3(new_n935), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n976), .B1(new_n998), .B2(new_n981), .ZN(new_n999));
  AND4_X1   g574(.A1(new_n976), .A2(new_n989), .A3(new_n897), .A4(new_n969), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT109), .B(new_n994), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n991), .B1(new_n995), .B2(new_n1002), .ZN(G397));
  NAND2_X1  g578(.A1(new_n483), .A2(G2105), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n468), .A2(new_n474), .A3(KEYINPUT69), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n478), .B1(new_n477), .B2(new_n467), .ZN(new_n1006));
  OAI211_X1 g581(.A(G40), .B(new_n1004), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(G160), .A2(KEYINPUT110), .A3(G40), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(G164), .B2(G1384), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n780), .A2(G2067), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n775), .A2(new_n782), .A3(new_n779), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT112), .ZN(new_n1019));
  INV_X1    g594(.A(new_n736), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1015), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT46), .B1(new_n1015), .B2(G1996), .ZN(new_n1022));
  OR3_X1    g597(.A1(new_n1015), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1024), .B(KEYINPUT47), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1014), .A2(G1996), .A3(new_n736), .ZN(new_n1026));
  XOR2_X1   g601(.A(new_n1026), .B(KEYINPUT111), .Z(new_n1027));
  OAI21_X1  g602(.A(new_n1019), .B1(G1996), .B2(new_n736), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1027), .B1(new_n1014), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n834), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n832), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1015), .B1(new_n1032), .B2(new_n1017), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n832), .B(new_n834), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1029), .B1(new_n1015), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(G290), .A2(G1986), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1014), .A2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1038), .B(KEYINPUT48), .ZN(new_n1039));
  AOI211_X1 g614(.A(new_n1025), .B(new_n1033), .C1(new_n1036), .C2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1042));
  INV_X1    g617(.A(G1384), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n882), .A2(KEYINPUT45), .A3(new_n1043), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1044), .A2(new_n1013), .ZN(new_n1045));
  AOI21_X1  g620(.A(G1971), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n882), .A2(new_n1047), .A3(new_n1043), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1009), .A2(new_n1010), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(G2090), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1041), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n526), .B2(new_n531), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1053), .B(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1009), .A2(new_n1010), .A3(new_n1044), .A4(new_n1013), .ZN(new_n1057));
  INV_X1    g632(.A(G1971), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1059), .B(KEYINPUT113), .C1(G2090), .C2(new_n1050), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1052), .A2(G8), .A3(new_n1056), .A4(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G8), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1050), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1065), .A2(new_n794), .B1(new_n1058), .B2(new_n1057), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1064), .B1(new_n1066), .B2(KEYINPUT113), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1067), .A2(KEYINPUT115), .A3(new_n1056), .A4(new_n1052), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1063), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(G164), .A2(G1384), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1009), .A2(new_n1010), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1072), .A2(new_n1064), .ZN(new_n1073));
  OAI21_X1  g648(.A(G1981), .B1(new_n814), .B2(new_n815), .ZN(new_n1074));
  INV_X1    g649(.A(G1981), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n606), .A2(new_n612), .A3(new_n1075), .A4(new_n613), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1074), .A2(new_n1076), .A3(KEYINPUT49), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT49), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n1080));
  INV_X1    g655(.A(G1976), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(G288), .B2(new_n1081), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n598), .A2(new_n602), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n594), .A2(new_n595), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1083), .A2(KEYINPUT116), .A3(new_n1084), .A4(G1976), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(G8), .A3(new_n1071), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1073), .A2(new_n1079), .B1(new_n1087), .B2(KEYINPUT52), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT52), .B1(G288), .B2(new_n1081), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1086), .A2(G8), .A3(new_n1071), .A4(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1088), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1048), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1070), .A2(KEYINPUT119), .A3(new_n1047), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1009), .A2(new_n1010), .A3(new_n1049), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1059), .B1(new_n1100), .B2(G2090), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1056), .B1(new_n1101), .B2(G8), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1094), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1069), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT126), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1069), .A2(new_n1103), .A3(KEYINPUT126), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n581), .A2(new_n583), .A3(new_n565), .ZN(new_n1109));
  XOR2_X1   g684(.A(new_n1109), .B(KEYINPUT57), .Z(new_n1110));
  OAI21_X1  g685(.A(new_n801), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT56), .B(G2072), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1042), .A2(new_n1045), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1110), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1111), .A2(new_n1110), .A3(new_n1113), .ZN(new_n1115));
  INV_X1    g690(.A(new_n630), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1072), .A2(new_n782), .ZN(new_n1117));
  INV_X1    g692(.A(G1348), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1050), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1116), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1114), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(G1996), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1042), .A2(new_n1122), .A3(new_n1045), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT58), .B(G1341), .Z(new_n1124));
  NAND2_X1  g699(.A1(new_n1071), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1126), .A2(KEYINPUT123), .A3(new_n555), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n1128));
  AOI211_X1 g703(.A(new_n1128), .B(new_n862), .C1(new_n1123), .C2(new_n1125), .ZN(new_n1129));
  OAI211_X1 g704(.A(KEYINPUT59), .B(new_n1127), .C1(new_n1129), .C2(KEYINPUT123), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1115), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1131), .B1(new_n1132), .B2(new_n1114), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1126), .A2(KEYINPUT124), .A3(new_n555), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1117), .A2(new_n1116), .A3(new_n1119), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT60), .B1(new_n1138), .B2(new_n1120), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1130), .A2(new_n1133), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1114), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1141), .A2(KEYINPUT61), .A3(new_n1115), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1116), .A2(KEYINPUT60), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1117), .A2(new_n1119), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1121), .B1(new_n1140), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n1147));
  OR3_X1    g722(.A1(new_n1050), .A2(new_n1147), .A3(G2084), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1147), .B1(new_n1050), .B2(G2084), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1057), .A2(new_n765), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(G286), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1148), .A2(G168), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(G8), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT51), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1155), .A2(KEYINPUT51), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1057), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT53), .B1(new_n1160), .B2(new_n753), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n1161), .A2(KEYINPUT125), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(KEYINPUT125), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1065), .A2(G1961), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(G301), .B(KEYINPUT54), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT53), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1007), .A2(new_n1167), .A3(G2078), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1166), .B1(new_n1045), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1160), .A2(KEYINPUT53), .A3(new_n753), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .A4(new_n1170), .ZN(new_n1171));
  AOI22_X1  g746(.A1(new_n1165), .A2(new_n1169), .B1(new_n1171), .B2(new_n1166), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1146), .A2(new_n1159), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT51), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1154), .A2(G8), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1174), .B1(new_n1175), .B2(new_n1152), .ZN(new_n1176));
  OAI21_X1  g751(.A(KEYINPUT62), .B1(new_n1176), .B2(new_n1157), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1156), .A2(new_n1158), .A3(new_n1178), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1171), .A2(G171), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1177), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1108), .B1(new_n1173), .B2(new_n1181), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1151), .A2(G8), .A3(G168), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1069), .A2(new_n1103), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT121), .ZN(new_n1185));
  AOI21_X1  g760(.A(KEYINPUT63), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1069), .A2(new_n1103), .A3(KEYINPUT121), .A4(new_n1183), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1056), .B1(new_n1067), .B2(new_n1052), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT122), .ZN(new_n1189));
  OR3_X1    g764(.A1(new_n1188), .A2(new_n1094), .A3(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1189), .B1(new_n1188), .B2(new_n1094), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1069), .A2(KEYINPUT63), .A3(new_n1183), .ZN(new_n1193));
  AOI22_X1  g768(.A1(new_n1186), .A2(new_n1187), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(G288), .A2(G1976), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1195), .B(KEYINPUT118), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1196), .B1(new_n1079), .B2(new_n1073), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1076), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1073), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1199), .B1(new_n1069), .B2(new_n1094), .ZN(new_n1200));
  NOR3_X1   g775(.A1(new_n1182), .A2(new_n1194), .A3(new_n1200), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n618), .A2(new_n836), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1014), .B1(new_n1037), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1036), .A2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1040), .B1(new_n1201), .B2(new_n1204), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g780(.A(new_n899), .ZN(new_n1207));
  NOR3_X1   g781(.A1(G229), .A2(new_n462), .A3(G227), .ZN(new_n1208));
  NAND2_X1  g782(.A1(new_n1208), .A2(new_n684), .ZN(new_n1209));
  INV_X1    g783(.A(KEYINPUT127), .ZN(new_n1210));
  NAND2_X1  g784(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g785(.A1(new_n1208), .A2(new_n684), .A3(KEYINPUT127), .ZN(new_n1212));
  AOI21_X1  g786(.A(new_n1207), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AND2_X1   g787(.A1(new_n1213), .A2(new_n993), .ZN(G308));
  NAND2_X1  g788(.A1(new_n1213), .A2(new_n993), .ZN(G225));
endmodule


