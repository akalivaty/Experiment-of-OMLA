//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n591, new_n592, new_n593, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n791, new_n793,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT27), .B(G183gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(KEYINPUT28), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n209), .ZN(new_n211));
  NOR2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(KEYINPUT26), .ZN(new_n213));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n212), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n210), .A2(new_n211), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n212), .B(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n220), .B(new_n214), .C1(KEYINPUT24), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(KEYINPUT24), .ZN(new_n223));
  INV_X1    g022(.A(G183gat), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n223), .B1(new_n224), .B2(new_n207), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT64), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT25), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT25), .ZN(new_n228));
  OAI211_X1 g027(.A(KEYINPUT64), .B(new_n228), .C1(new_n222), .C2(new_n225), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n218), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G226gat), .A2(G233gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(KEYINPUT74), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(new_n230), .B2(KEYINPUT29), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n232), .B1(new_n235), .B2(KEYINPUT75), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n227), .A2(new_n229), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(new_n217), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT29), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT75), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(new_n241), .A3(new_n234), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n236), .A2(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(KEYINPUT71), .B(G197gat), .Z(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G204gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT22), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT72), .B(G218gat), .ZN(new_n247));
  INV_X1    g046(.A(G211gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT71), .B(G197gat), .ZN(new_n250));
  INV_X1    g049(.A(G204gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n245), .A2(new_n249), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G211gat), .B(G218gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(KEYINPUT73), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n253), .B(new_n255), .Z(new_n256));
  NAND2_X1  g055(.A1(new_n243), .A2(new_n256), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n240), .A2(new_n231), .B1(new_n238), .B2(new_n233), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n253), .B(new_n255), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n205), .B1(new_n261), .B2(KEYINPUT37), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT37), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n263), .B1(new_n257), .B2(new_n260), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT38), .ZN(new_n266));
  XOR2_X1   g065(.A(G141gat), .B(G148gat), .Z(new_n267));
  INV_X1    g066(.A(G155gat), .ZN(new_n268));
  INV_X1    g067(.A(G162gat), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT2), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G155gat), .B(G162gat), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n271), .B(new_n272), .Z(new_n273));
  XNOR2_X1  g072(.A(G127gat), .B(G134gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT66), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT1), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(G113gat), .B(G120gat), .Z(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(new_n276), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n277), .B(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n273), .B(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G225gat), .A2(G233gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  OR3_X1    g083(.A1(new_n273), .A2(new_n280), .A3(KEYINPUT4), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT77), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT4), .B1(new_n273), .B2(new_n280), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n271), .B(new_n272), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT3), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n289), .A2(new_n280), .A3(new_n292), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n293), .B(new_n282), .C1(new_n287), .C2(new_n286), .ZN(new_n294));
  OAI211_X1 g093(.A(KEYINPUT5), .B(new_n284), .C1(new_n288), .C2(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n283), .A2(KEYINPUT5), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT78), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n285), .A2(new_n297), .A3(new_n287), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n297), .B1(new_n285), .B2(new_n287), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n293), .B(new_n296), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G1gat), .B(G29gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n302), .B(KEYINPUT0), .ZN(new_n303));
  XNOR2_X1  g102(.A(G57gat), .B(G85gat), .ZN(new_n304));
  XOR2_X1   g103(.A(new_n303), .B(new_n304), .Z(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT6), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n295), .A2(new_n300), .A3(new_n305), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n301), .A2(KEYINPUT6), .A3(new_n306), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n257), .A2(new_n260), .A3(new_n204), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n263), .B1(new_n258), .B2(new_n256), .ZN(new_n315));
  INV_X1    g114(.A(new_n243), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n315), .B1(new_n316), .B2(new_n256), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT82), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n262), .A2(KEYINPUT38), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n266), .A2(new_n313), .A3(new_n314), .A4(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G78gat), .B(G106gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n322), .B(G22gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n259), .B1(new_n239), .B2(new_n292), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n291), .B1(new_n256), .B2(KEYINPUT29), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n325), .B1(new_n326), .B2(new_n273), .ZN(new_n327));
  INV_X1    g126(.A(G228gat), .ZN(new_n328));
  INV_X1    g127(.A(G233gat), .ZN(new_n329));
  NOR3_X1   g128(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT29), .B1(new_n253), .B2(new_n254), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(new_n254), .B2(new_n253), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n290), .B1(new_n332), .B2(new_n291), .ZN(new_n333));
  AOI211_X1 g132(.A(new_n333), .B(new_n325), .C1(G228gat), .C2(G233gat), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT79), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NOR3_X1   g135(.A1(new_n330), .A2(new_n334), .A3(KEYINPUT79), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT31), .B(G50gat), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n338), .ZN(new_n340));
  OR3_X1    g139(.A1(new_n330), .A2(new_n334), .A3(KEYINPUT79), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n340), .B1(new_n341), .B2(new_n335), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n324), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n338), .B1(new_n336), .B2(new_n337), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n341), .A2(new_n335), .A3(new_n340), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(new_n323), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n293), .B1(new_n298), .B2(new_n299), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT39), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(new_n283), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n350), .A2(new_n305), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(new_n283), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n352), .B(KEYINPUT39), .C1(new_n283), .C2(new_n281), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT40), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT80), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n351), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n307), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n355), .B1(new_n351), .B2(new_n353), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT30), .ZN(new_n360));
  OR2_X1    g159(.A1(new_n314), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n314), .A2(new_n360), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n261), .A2(new_n205), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n365), .A2(KEYINPUT81), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT81), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(new_n359), .B2(new_n364), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n321), .B(new_n347), .C1(new_n366), .C2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n363), .B1(new_n314), .B2(new_n360), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT76), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT76), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n361), .A2(new_n372), .A3(new_n363), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n371), .A2(new_n373), .A3(new_n312), .A4(new_n362), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n343), .A2(new_n346), .ZN(new_n375));
  XOR2_X1   g174(.A(G15gat), .B(G43gat), .Z(new_n376));
  XNOR2_X1  g175(.A(G71gat), .B(G99gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(G227gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(new_n329), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n238), .A2(new_n280), .ZN(new_n384));
  INV_X1    g183(.A(new_n280), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n230), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n383), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT32), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n380), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OR3_X1    g188(.A1(new_n387), .A2(KEYINPUT67), .A3(KEYINPUT33), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT67), .B1(new_n387), .B2(KEYINPUT33), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n384), .A2(new_n383), .A3(new_n386), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT34), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n380), .A2(KEYINPUT70), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n380), .A2(KEYINPUT70), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n396), .A2(KEYINPUT33), .ZN(new_n397));
  AOI211_X1 g196(.A(new_n388), .B(new_n387), .C1(new_n395), .C2(new_n397), .ZN(new_n398));
  OR3_X1    g197(.A1(new_n392), .A2(new_n394), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n394), .B1(new_n392), .B2(new_n398), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT36), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n399), .A2(new_n400), .A3(KEYINPUT36), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n374), .A2(new_n375), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n369), .A2(new_n405), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n399), .A2(new_n400), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n347), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT35), .B1(new_n408), .B2(new_n374), .ZN(new_n409));
  INV_X1    g208(.A(new_n364), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n313), .A2(KEYINPUT35), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n407), .A2(new_n347), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n406), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G15gat), .B(G22gat), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT16), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n415), .B1(new_n416), .B2(G1gat), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n417), .B(KEYINPUT87), .C1(G1gat), .C2(new_n415), .ZN(new_n418));
  INV_X1    g217(.A(G8gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT91), .ZN(new_n422));
  XNOR2_X1  g221(.A(G57gat), .B(G64gat), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G71gat), .B(G78gat), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n422), .B(new_n426), .C1(new_n423), .C2(new_n424), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n421), .B1(KEYINPUT21), .B2(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(new_n268), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n433), .B(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n430), .A2(KEYINPUT21), .ZN(new_n437));
  NAND2_X1  g236(.A1(G231gat), .A2(G233gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(G127gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(G183gat), .B(G211gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n436), .B(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT17), .ZN(new_n445));
  INV_X1    g244(.A(G29gat), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n446), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT14), .B(G29gat), .ZN(new_n448));
  INV_X1    g247(.A(G36gat), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AND2_X1   g249(.A1(G43gat), .A2(G50gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(G43gat), .A2(G50gat), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT15), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(G43gat), .ZN(new_n454));
  INV_X1    g253(.A(G50gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT15), .ZN(new_n457));
  NAND2_X1  g256(.A1(G43gat), .A2(G50gat), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT85), .B1(new_n450), .B2(new_n460), .ZN(new_n461));
  AND2_X1   g260(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n462));
  NOR2_X1   g261(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n449), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n446), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT85), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n466), .A2(new_n467), .A3(new_n453), .A4(new_n459), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n461), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT84), .B1(new_n466), .B2(new_n453), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT84), .ZN(new_n471));
  INV_X1    g270(.A(new_n453), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n450), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n445), .B1(new_n475), .B2(KEYINPUT88), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT88), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n461), .A2(new_n468), .B1(new_n470), .B2(new_n473), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n477), .B1(new_n478), .B2(KEYINPUT86), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n477), .B(new_n445), .C1(new_n478), .C2(KEYINPUT86), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(G99gat), .A2(G106gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT8), .ZN(new_n484));
  NAND2_X1  g283(.A1(G85gat), .A2(G92gat), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT7), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(G85gat), .ZN(new_n488));
  INV_X1    g287(.A(G92gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n484), .A2(new_n487), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G99gat), .B(G106gat), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AOI22_X1  g294(.A1(KEYINPUT8), .A2(new_n483), .B1(new_n488), .B2(new_n489), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n496), .A2(new_n493), .A3(new_n487), .A4(new_n491), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n498), .ZN(new_n500));
  NAND2_X1  g299(.A1(G232gat), .A2(G233gat), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n475), .A2(new_n500), .B1(KEYINPUT41), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G190gat), .B(G218gat), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n505), .B(KEYINPUT94), .Z(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n502), .A2(KEYINPUT41), .ZN(new_n508));
  XNOR2_X1  g307(.A(G134gat), .B(G162gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n506), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n499), .A2(new_n511), .A3(new_n503), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n507), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n510), .B1(new_n507), .B2(new_n512), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n444), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT86), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT88), .B1(new_n475), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT17), .B1(new_n478), .B2(new_n477), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n481), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n420), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G229gat), .A2(G233gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n420), .A2(new_n478), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n523), .A2(KEYINPUT18), .A3(new_n524), .A4(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT89), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n525), .B1(new_n482), .B2(new_n420), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n530), .A2(KEYINPUT89), .A3(KEYINPUT18), .A4(new_n524), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n524), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT18), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT90), .B1(new_n421), .B2(new_n475), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(new_n526), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n524), .B(KEYINPUT13), .Z(new_n537));
  AOI22_X1  g336(.A1(new_n533), .A2(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G113gat), .B(G141gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(G197gat), .ZN(new_n540));
  XOR2_X1   g339(.A(KEYINPUT11), .B(G169gat), .Z(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n542), .B(new_n543), .Z(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n532), .A2(new_n538), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n545), .B1(new_n532), .B2(new_n538), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G230gat), .A2(G233gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT95), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n493), .B1(new_n492), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT96), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n496), .A2(KEYINPUT95), .A3(new_n487), .A4(new_n491), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n551), .A2(new_n553), .B1(new_n552), .B2(new_n497), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n430), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n430), .A2(new_n498), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT10), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n500), .A2(new_n430), .A3(KEYINPUT10), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n549), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n549), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n556), .A2(new_n558), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G120gat), .B(G148gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(G176gat), .B(G204gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n565), .A2(new_n568), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR3_X1   g371(.A1(new_n517), .A2(new_n548), .A3(new_n572), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n414), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n313), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(G1gat), .ZN(G1324gat));
  AND3_X1   g375(.A1(new_n414), .A2(new_n364), .A3(new_n573), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(new_n419), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT97), .ZN(new_n579));
  XOR2_X1   g378(.A(KEYINPUT16), .B(G8gat), .Z(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT42), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(new_n582), .ZN(G1325gat));
  INV_X1    g382(.A(G15gat), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n574), .A2(new_n584), .A3(new_n407), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n403), .A2(new_n404), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n574), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n585), .B1(new_n588), .B2(new_n584), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n589), .B(KEYINPUT98), .Z(G1326gat));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n375), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT99), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT43), .B(G22gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(G1327gat));
  AOI22_X1  g393(.A1(new_n369), .A2(new_n405), .B1(new_n409), .B2(new_n412), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(new_n516), .ZN(new_n596));
  NOR3_X1   g395(.A1(new_n548), .A2(new_n444), .A3(new_n572), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n596), .A2(new_n446), .A3(new_n313), .A4(new_n597), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n598), .A2(KEYINPUT100), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT45), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(KEYINPUT100), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n600), .B1(new_n599), .B2(new_n601), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT44), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n604), .B1(new_n595), .B2(new_n516), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n374), .A2(new_n375), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n586), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n365), .B(KEYINPUT81), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n313), .A2(new_n314), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n609), .B1(new_n265), .B2(KEYINPUT38), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n375), .B1(new_n610), .B2(new_n320), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n607), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n409), .A2(new_n412), .ZN(new_n613));
  OAI211_X1 g412(.A(KEYINPUT44), .B(new_n515), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  AND4_X1   g413(.A1(new_n313), .A2(new_n605), .A3(new_n614), .A4(new_n597), .ZN(new_n615));
  OAI22_X1  g414(.A1(new_n602), .A2(new_n603), .B1(new_n446), .B2(new_n615), .ZN(G1328gat));
  NOR2_X1   g415(.A1(new_n410), .A2(G36gat), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n414), .A2(new_n515), .A3(new_n597), .A4(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT101), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n596), .A2(KEYINPUT101), .A3(new_n597), .A4(new_n617), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT46), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT102), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n622), .B1(new_n620), .B2(new_n621), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n605), .A2(new_n614), .A3(new_n364), .A4(new_n597), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n626), .B1(G36gat), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(G1329gat));
  NAND4_X1  g428(.A1(new_n605), .A2(new_n614), .A3(new_n587), .A4(new_n597), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(G43gat), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT103), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT47), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n596), .A2(new_n597), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(new_n454), .A3(new_n407), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n631), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n633), .B(new_n636), .ZN(G1330gat));
  INV_X1    g436(.A(KEYINPUT104), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n634), .A2(new_n455), .A3(new_n375), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n605), .A2(new_n614), .A3(new_n375), .A4(new_n597), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(G50gat), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n638), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT105), .B(KEYINPUT48), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n642), .B(new_n644), .ZN(G1331gat));
  NAND2_X1  g444(.A1(new_n532), .A2(new_n538), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n544), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n532), .A2(new_n538), .A3(new_n545), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n517), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n572), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT106), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n414), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(new_n312), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT107), .B(G57gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1332gat));
  NOR2_X1   g455(.A1(new_n653), .A2(new_n410), .ZN(new_n657));
  NOR2_X1   g456(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n658));
  AND2_X1   g457(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n660), .B1(new_n657), .B2(new_n658), .ZN(G1333gat));
  INV_X1    g460(.A(new_n653), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n662), .A2(G71gat), .A3(new_n587), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n401), .B(KEYINPUT108), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n653), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n663), .B1(G71gat), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g466(.A1(new_n662), .A2(new_n375), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G78gat), .ZN(G1335gat));
  INV_X1    g468(.A(new_n572), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n649), .A2(new_n444), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n605), .A2(new_n614), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT109), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT109), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n605), .A2(new_n614), .A3(new_n674), .A4(new_n671), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n673), .A2(new_n313), .A3(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n649), .A2(new_n444), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n515), .B(new_n677), .C1(new_n612), .C2(new_n613), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT51), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(KEYINPUT110), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n414), .A2(new_n515), .A3(new_n677), .A4(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n681), .A2(new_n572), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n313), .A2(new_n488), .ZN(new_n685));
  OAI22_X1  g484(.A1(new_n676), .A2(new_n488), .B1(new_n684), .B2(new_n685), .ZN(G1336gat));
  INV_X1    g485(.A(KEYINPUT52), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n687), .B(G92gat), .C1(new_n672), .C2(new_n410), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n410), .A2(G92gat), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  OAI221_X1 g489(.A(new_n688), .B1(KEYINPUT111), .B2(new_n687), .C1(new_n684), .C2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n673), .A2(new_n364), .A3(new_n675), .ZN(new_n692));
  AND4_X1   g491(.A1(new_n572), .A2(new_n681), .A3(new_n683), .A4(new_n689), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT111), .ZN(new_n694));
  AOI22_X1  g493(.A1(new_n692), .A2(G92gat), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n691), .B1(new_n695), .B2(new_n687), .ZN(G1337gat));
  AND3_X1   g495(.A1(new_n673), .A2(new_n587), .A3(new_n675), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT112), .B(G99gat), .Z(new_n698));
  NAND2_X1  g497(.A1(new_n407), .A2(new_n698), .ZN(new_n699));
  OAI22_X1  g498(.A1(new_n697), .A2(new_n698), .B1(new_n684), .B2(new_n699), .ZN(G1338gat));
  INV_X1    g499(.A(KEYINPUT53), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n701), .B(G106gat), .C1(new_n672), .C2(new_n347), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n347), .A2(G106gat), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n681), .A2(new_n683), .A3(new_n572), .A4(new_n703), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n702), .B(new_n704), .C1(KEYINPUT113), .C2(new_n701), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n673), .A2(new_n375), .A3(new_n675), .ZN(new_n706));
  INV_X1    g505(.A(new_n704), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT113), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n706), .A2(G106gat), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n705), .B1(new_n709), .B2(new_n701), .ZN(G1339gat));
  NAND2_X1  g509(.A1(new_n650), .A2(new_n670), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT54), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n712), .B(new_n549), .C1(new_n559), .C2(new_n561), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n568), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(KEYINPUT115), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT115), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n713), .A2(new_n716), .A3(new_n568), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT114), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n560), .A2(new_n563), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT54), .B1(new_n559), .B2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT10), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n428), .A2(new_n429), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n492), .A2(new_n550), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n724), .A2(new_n553), .A3(new_n494), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n497), .A2(new_n552), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n723), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n722), .B1(new_n729), .B2(new_n557), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n563), .B1(new_n730), .B2(new_n560), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n719), .B1(new_n721), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n720), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n712), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n562), .A2(new_n734), .A3(KEYINPUT114), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT55), .B1(new_n718), .B2(new_n736), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n721), .A2(new_n731), .A3(new_n719), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT114), .B1(new_n562), .B2(new_n734), .ZN(new_n739));
  OAI21_X1  g538(.A(KEYINPUT55), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n713), .A2(new_n716), .A3(new_n568), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n716), .B1(new_n713), .B2(new_n568), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n570), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT116), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT55), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n746), .B1(new_n732), .B2(new_n735), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n569), .B1(new_n718), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT116), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n737), .B1(new_n745), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n536), .A2(new_n537), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n530), .A2(new_n524), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n542), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n751), .A2(new_n648), .A3(new_n515), .A4(new_n754), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n648), .A2(new_n572), .A3(new_n754), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n756), .B1(new_n751), .B2(new_n649), .ZN(new_n757));
  OAI211_X1 g556(.A(KEYINPUT117), .B(new_n755), .C1(new_n757), .C2(new_n515), .ZN(new_n758));
  INV_X1    g557(.A(new_n444), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n648), .A2(new_n572), .A3(new_n754), .ZN(new_n761));
  INV_X1    g560(.A(new_n737), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n718), .A2(new_n747), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n749), .B1(new_n763), .B2(new_n570), .ZN(new_n764));
  AOI211_X1 g563(.A(KEYINPUT116), .B(new_n569), .C1(new_n718), .C2(new_n747), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n761), .B1(new_n766), .B2(new_n548), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n516), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT117), .B1(new_n768), .B2(new_n755), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n711), .B1(new_n760), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n313), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n771), .A2(new_n364), .A3(new_n408), .ZN(new_n772));
  INV_X1    g571(.A(G113gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(new_n773), .A3(new_n649), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n751), .A2(new_n649), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n515), .B1(new_n776), .B2(new_n761), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n515), .A2(new_n648), .A3(new_n754), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n766), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n775), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n780), .A2(new_n759), .A3(new_n758), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n375), .B1(new_n781), .B2(new_n711), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n410), .A2(new_n313), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n783), .A2(new_n401), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(G113gat), .B1(new_n785), .B2(new_n548), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n774), .A2(new_n786), .ZN(new_n787));
  XOR2_X1   g586(.A(new_n787), .B(KEYINPUT118), .Z(G1340gat));
  AOI21_X1  g587(.A(G120gat), .B1(new_n772), .B2(new_n572), .ZN(new_n789));
  INV_X1    g588(.A(G120gat), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n785), .A2(new_n790), .A3(new_n670), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n789), .A2(new_n791), .ZN(G1341gat));
  NAND3_X1  g591(.A1(new_n772), .A2(new_n440), .A3(new_n444), .ZN(new_n793));
  OAI21_X1  g592(.A(G127gat), .B1(new_n785), .B2(new_n759), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(G1342gat));
  NAND2_X1  g594(.A1(new_n410), .A2(new_n515), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n408), .A2(new_n796), .A3(G134gat), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n770), .A2(new_n313), .A3(new_n797), .ZN(new_n798));
  XOR2_X1   g597(.A(new_n798), .B(KEYINPUT119), .Z(new_n799));
  OR2_X1    g598(.A1(new_n799), .A2(KEYINPUT56), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(KEYINPUT56), .ZN(new_n801));
  OAI21_X1  g600(.A(G134gat), .B1(new_n785), .B2(new_n516), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(G1343gat));
  NOR2_X1   g602(.A1(new_n587), .A2(new_n783), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT57), .B1(new_n770), .B2(new_n375), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n375), .A2(KEYINPUT57), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n762), .B(new_n748), .C1(new_n546), .C2(new_n547), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n515), .B1(new_n807), .B2(new_n761), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n759), .B1(new_n808), .B2(new_n779), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n806), .B1(new_n809), .B2(new_n711), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n804), .B1(new_n805), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(G141gat), .B1(new_n811), .B2(new_n548), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n771), .A2(KEYINPUT121), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT121), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n770), .A2(new_n815), .A3(new_n313), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n587), .A2(new_n347), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n814), .A2(new_n410), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n548), .A2(G141gat), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n812), .B(new_n813), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n811), .A2(KEYINPUT120), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n823), .B(new_n804), .C1(new_n805), .C2(new_n810), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n822), .A2(new_n649), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n821), .B1(new_n825), .B2(G141gat), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n820), .B1(new_n826), .B2(new_n813), .ZN(G1344gat));
  NAND3_X1  g626(.A1(new_n822), .A2(new_n572), .A3(new_n824), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(G148gat), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT122), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n804), .A2(new_n572), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n806), .B1(new_n781), .B2(new_n711), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n809), .A2(new_n711), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT57), .B1(new_n836), .B2(new_n375), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n834), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  AOI211_X1 g637(.A(new_n832), .B(new_n829), .C1(new_n838), .C2(G148gat), .ZN(new_n839));
  INV_X1    g638(.A(new_n806), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n837), .B1(new_n770), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(G148gat), .B1(new_n841), .B2(new_n833), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT122), .B1(new_n842), .B2(KEYINPUT59), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n831), .A2(new_n844), .ZN(new_n845));
  OR3_X1    g644(.A1(new_n818), .A2(G148gat), .A3(new_n670), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1345gat));
  NOR2_X1   g646(.A1(new_n818), .A2(new_n759), .ZN(new_n848));
  AOI21_X1  g647(.A(G155gat), .B1(new_n848), .B2(KEYINPUT123), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT123), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(new_n818), .B2(new_n759), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n822), .A2(new_n824), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n759), .A2(new_n268), .ZN(new_n854));
  AOI22_X1  g653(.A1(new_n849), .A2(new_n851), .B1(new_n853), .B2(new_n854), .ZN(G1346gat));
  OAI21_X1  g654(.A(G162gat), .B1(new_n852), .B2(new_n516), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n796), .A2(G162gat), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n814), .A2(new_n816), .A3(new_n817), .A4(new_n857), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT124), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n856), .A2(new_n859), .ZN(G1347gat));
  NAND2_X1  g659(.A1(new_n364), .A2(new_n312), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n664), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n782), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(G169gat), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n863), .A2(new_n864), .A3(new_n548), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n408), .A2(new_n861), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n770), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(G169gat), .B1(new_n867), .B2(new_n649), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n865), .A2(new_n868), .ZN(G1348gat));
  OAI21_X1  g668(.A(G176gat), .B1(new_n863), .B2(new_n670), .ZN(new_n870));
  INV_X1    g669(.A(new_n867), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n670), .A2(G176gat), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(G1349gat));
  OAI21_X1  g672(.A(G183gat), .B1(new_n863), .B2(new_n759), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT125), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n867), .A2(new_n206), .A3(new_n444), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g677(.A1(new_n867), .A2(new_n207), .A3(new_n515), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n782), .A2(new_n515), .A3(new_n862), .ZN(new_n880));
  XNOR2_X1  g679(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n880), .A2(G190gat), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n880), .B2(G190gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n879), .B1(new_n882), .B2(new_n883), .ZN(G1351gat));
  NOR2_X1   g683(.A1(new_n587), .A2(new_n861), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n770), .A2(new_n375), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(G197gat), .B1(new_n886), .B2(new_n649), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n841), .A2(new_n587), .A3(new_n861), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n649), .A2(G197gat), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(G1352gat));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n572), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G204gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n886), .A2(new_n251), .A3(new_n572), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n893), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT127), .B1(new_n893), .B2(KEYINPUT62), .ZN(new_n895));
  OAI221_X1 g694(.A(new_n892), .B1(KEYINPUT62), .B2(new_n893), .C1(new_n894), .C2(new_n895), .ZN(G1353gat));
  NAND3_X1  g695(.A1(new_n886), .A2(new_n248), .A3(new_n444), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n888), .A2(new_n444), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n898), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT63), .B1(new_n898), .B2(G211gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(G1354gat));
  AOI21_X1  g700(.A(G218gat), .B1(new_n886), .B2(new_n515), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n516), .A2(new_n247), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n888), .B2(new_n903), .ZN(G1355gat));
endmodule


