

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U549 ( .A1(n655), .A2(n654), .ZN(n669) );
  NOR2_X1 U550 ( .A1(n671), .A2(n667), .ZN(n646) );
  NAND2_X1 U551 ( .A1(n685), .A2(n588), .ZN(n658) );
  XNOR2_X1 U552 ( .A(n645), .B(KEYINPUT94), .ZN(n657) );
  BUF_X1 U553 ( .A(n657), .Z(n682) );
  INV_X1 U554 ( .A(n910), .ZN(n717) );
  NAND2_X1 U555 ( .A1(n718), .A2(n717), .ZN(n719) );
  AND2_X1 U556 ( .A1(n525), .A2(n524), .ZN(G164) );
  INV_X1 U557 ( .A(G2105), .ZN(n515) );
  NOR2_X1 U558 ( .A1(G2104), .A2(n515), .ZN(n880) );
  NAND2_X1 U559 ( .A1(G126), .A2(n880), .ZN(n517) );
  AND2_X1 U560 ( .A1(n515), .A2(G2104), .ZN(n885) );
  NAND2_X1 U561 ( .A1(G102), .A2(n885), .ZN(n516) );
  NAND2_X1 U562 ( .A1(n517), .A2(n516), .ZN(n521) );
  NAND2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  XNOR2_X1 U564 ( .A(n518), .B(KEYINPUT65), .ZN(n878) );
  NAND2_X1 U565 ( .A1(n878), .A2(G114), .ZN(n519) );
  XNOR2_X1 U566 ( .A(n519), .B(KEYINPUT87), .ZN(n520) );
  NOR2_X1 U567 ( .A1(n521), .A2(n520), .ZN(n525) );
  NOR2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XOR2_X2 U569 ( .A(KEYINPUT17), .B(n522), .Z(n884) );
  NAND2_X1 U570 ( .A1(G138), .A2(n884), .ZN(n523) );
  XNOR2_X1 U571 ( .A(n523), .B(KEYINPUT88), .ZN(n524) );
  INV_X1 U572 ( .A(G651), .ZN(n529) );
  NOR2_X1 U573 ( .A1(G543), .A2(n529), .ZN(n526) );
  XOR2_X1 U574 ( .A(KEYINPUT1), .B(n526), .Z(n793) );
  NAND2_X1 U575 ( .A1(G64), .A2(n793), .ZN(n528) );
  XOR2_X1 U576 ( .A(G543), .B(KEYINPUT0), .Z(n566) );
  NOR2_X2 U577 ( .A1(G651), .A2(n566), .ZN(n794) );
  NAND2_X1 U578 ( .A1(G52), .A2(n794), .ZN(n527) );
  NAND2_X1 U579 ( .A1(n528), .A2(n527), .ZN(n536) );
  NOR2_X1 U580 ( .A1(n566), .A2(n529), .ZN(n790) );
  NAND2_X1 U581 ( .A1(n790), .A2(G77), .ZN(n530) );
  XNOR2_X1 U582 ( .A(n530), .B(KEYINPUT68), .ZN(n532) );
  NOR2_X1 U583 ( .A1(G651), .A2(G543), .ZN(n789) );
  NAND2_X1 U584 ( .A1(G90), .A2(n789), .ZN(n531) );
  NAND2_X1 U585 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U586 ( .A(KEYINPUT69), .B(n533), .ZN(n534) );
  XNOR2_X1 U587 ( .A(KEYINPUT9), .B(n534), .ZN(n535) );
  NOR2_X1 U588 ( .A1(n536), .A2(n535), .ZN(G171) );
  NAND2_X1 U589 ( .A1(n884), .A2(G137), .ZN(n539) );
  NAND2_X1 U590 ( .A1(G101), .A2(n885), .ZN(n537) );
  XOR2_X1 U591 ( .A(KEYINPUT23), .B(n537), .Z(n538) );
  NAND2_X1 U592 ( .A1(n539), .A2(n538), .ZN(n543) );
  NAND2_X1 U593 ( .A1(G125), .A2(n880), .ZN(n541) );
  NAND2_X1 U594 ( .A1(G113), .A2(n878), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U596 ( .A1(n543), .A2(n542), .ZN(G160) );
  NAND2_X1 U597 ( .A1(G89), .A2(n789), .ZN(n544) );
  XNOR2_X1 U598 ( .A(n544), .B(KEYINPUT4), .ZN(n545) );
  XNOR2_X1 U599 ( .A(n545), .B(KEYINPUT76), .ZN(n547) );
  NAND2_X1 U600 ( .A1(G76), .A2(n790), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U602 ( .A(KEYINPUT5), .B(n548), .ZN(n556) );
  NAND2_X1 U603 ( .A1(G51), .A2(n794), .ZN(n551) );
  NAND2_X1 U604 ( .A1(n793), .A2(G63), .ZN(n549) );
  XOR2_X1 U605 ( .A(KEYINPUT77), .B(n549), .Z(n550) );
  NAND2_X1 U606 ( .A1(n551), .A2(n550), .ZN(n554) );
  XNOR2_X1 U607 ( .A(KEYINPUT78), .B(KEYINPUT79), .ZN(n552) );
  XNOR2_X1 U608 ( .A(n552), .B(KEYINPUT6), .ZN(n553) );
  XNOR2_X1 U609 ( .A(n554), .B(n553), .ZN(n555) );
  NAND2_X1 U610 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U611 ( .A(KEYINPUT7), .B(n557), .ZN(G168) );
  XOR2_X1 U612 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U613 ( .A1(G88), .A2(n789), .ZN(n559) );
  NAND2_X1 U614 ( .A1(G75), .A2(n790), .ZN(n558) );
  NAND2_X1 U615 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U616 ( .A1(G62), .A2(n793), .ZN(n561) );
  NAND2_X1 U617 ( .A1(G50), .A2(n794), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U619 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U620 ( .A(KEYINPUT84), .B(n564), .Z(G303) );
  NAND2_X1 U621 ( .A1(G49), .A2(n794), .ZN(n565) );
  XNOR2_X1 U622 ( .A(n565), .B(KEYINPUT82), .ZN(n571) );
  NAND2_X1 U623 ( .A1(G87), .A2(n566), .ZN(n568) );
  NAND2_X1 U624 ( .A1(G74), .A2(G651), .ZN(n567) );
  NAND2_X1 U625 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U626 ( .A1(n793), .A2(n569), .ZN(n570) );
  NAND2_X1 U627 ( .A1(n571), .A2(n570), .ZN(G288) );
  NAND2_X1 U628 ( .A1(n794), .A2(G48), .ZN(n578) );
  NAND2_X1 U629 ( .A1(G61), .A2(n793), .ZN(n573) );
  NAND2_X1 U630 ( .A1(G86), .A2(n789), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U632 ( .A1(n790), .A2(G73), .ZN(n574) );
  XOR2_X1 U633 ( .A(KEYINPUT2), .B(n574), .Z(n575) );
  NOR2_X1 U634 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U635 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U636 ( .A(KEYINPUT83), .B(n579), .Z(G305) );
  INV_X1 U637 ( .A(G303), .ZN(G166) );
  NAND2_X1 U638 ( .A1(n793), .A2(G60), .ZN(n580) );
  XNOR2_X1 U639 ( .A(n580), .B(KEYINPUT66), .ZN(n582) );
  NAND2_X1 U640 ( .A1(G47), .A2(n794), .ZN(n581) );
  NAND2_X1 U641 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U642 ( .A(KEYINPUT67), .B(n583), .ZN(n587) );
  NAND2_X1 U643 ( .A1(G85), .A2(n789), .ZN(n585) );
  NAND2_X1 U644 ( .A1(G72), .A2(n790), .ZN(n584) );
  AND2_X1 U645 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U646 ( .A1(n587), .A2(n586), .ZN(G290) );
  NOR2_X1 U647 ( .A1(G164), .A2(G1384), .ZN(n685) );
  NAND2_X1 U648 ( .A1(G160), .A2(G40), .ZN(n684) );
  INV_X1 U649 ( .A(n684), .ZN(n588) );
  XNOR2_X1 U650 ( .A(G2078), .B(KEYINPUT25), .ZN(n941) );
  NOR2_X1 U651 ( .A1(n658), .A2(n941), .ZN(n590) );
  INV_X1 U652 ( .A(n658), .ZN(n632) );
  INV_X1 U653 ( .A(G1961), .ZN(n965) );
  NOR2_X1 U654 ( .A1(n632), .A2(n965), .ZN(n589) );
  NOR2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n650) );
  AND2_X1 U656 ( .A1(G171), .A2(n650), .ZN(n591) );
  XNOR2_X1 U657 ( .A(KEYINPUT95), .B(n591), .ZN(n644) );
  XNOR2_X1 U658 ( .A(KEYINPUT99), .B(KEYINPUT29), .ZN(n642) );
  NAND2_X1 U659 ( .A1(n789), .A2(G81), .ZN(n592) );
  XNOR2_X1 U660 ( .A(n592), .B(KEYINPUT12), .ZN(n594) );
  NAND2_X1 U661 ( .A1(G68), .A2(n790), .ZN(n593) );
  NAND2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n596) );
  XOR2_X1 U663 ( .A(KEYINPUT13), .B(KEYINPUT72), .Z(n595) );
  XNOR2_X1 U664 ( .A(n596), .B(n595), .ZN(n599) );
  NAND2_X1 U665 ( .A1(n793), .A2(G56), .ZN(n597) );
  XOR2_X1 U666 ( .A(KEYINPUT14), .B(n597), .Z(n598) );
  NOR2_X1 U667 ( .A1(n599), .A2(n598), .ZN(n601) );
  NAND2_X1 U668 ( .A1(n794), .A2(G43), .ZN(n600) );
  NAND2_X1 U669 ( .A1(n601), .A2(n600), .ZN(n920) );
  NAND2_X1 U670 ( .A1(n658), .A2(G1341), .ZN(n605) );
  XNOR2_X1 U671 ( .A(G1996), .B(KEYINPUT97), .ZN(n935) );
  NOR2_X1 U672 ( .A1(n658), .A2(n935), .ZN(n603) );
  XOR2_X1 U673 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n602) );
  XNOR2_X1 U674 ( .A(n603), .B(n602), .ZN(n604) );
  NAND2_X1 U675 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U676 ( .A1(n920), .A2(n606), .ZN(n618) );
  NAND2_X1 U677 ( .A1(n794), .A2(G54), .ZN(n607) );
  XOR2_X1 U678 ( .A(KEYINPUT73), .B(n607), .Z(n609) );
  NAND2_X1 U679 ( .A1(n790), .A2(G79), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U681 ( .A(KEYINPUT74), .B(n610), .ZN(n614) );
  NAND2_X1 U682 ( .A1(G66), .A2(n793), .ZN(n612) );
  NAND2_X1 U683 ( .A1(G92), .A2(n789), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U685 ( .A1(n614), .A2(n613), .ZN(n616) );
  XNOR2_X1 U686 ( .A(KEYINPUT75), .B(KEYINPUT15), .ZN(n615) );
  XNOR2_X1 U687 ( .A(n616), .B(n615), .ZN(n908) );
  NOR2_X1 U688 ( .A1(n618), .A2(n908), .ZN(n617) );
  XOR2_X1 U689 ( .A(n617), .B(KEYINPUT98), .Z(n624) );
  NAND2_X1 U690 ( .A1(n618), .A2(n908), .ZN(n622) );
  NOR2_X1 U691 ( .A1(n632), .A2(G1348), .ZN(n620) );
  NOR2_X1 U692 ( .A1(G2067), .A2(n658), .ZN(n619) );
  NOR2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U694 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U695 ( .A1(n624), .A2(n623), .ZN(n636) );
  NAND2_X1 U696 ( .A1(G65), .A2(n793), .ZN(n626) );
  NAND2_X1 U697 ( .A1(G53), .A2(n794), .ZN(n625) );
  NAND2_X1 U698 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U699 ( .A1(G91), .A2(n789), .ZN(n628) );
  NAND2_X1 U700 ( .A1(G78), .A2(n790), .ZN(n627) );
  NAND2_X1 U701 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U702 ( .A1(n630), .A2(n629), .ZN(n801) );
  NAND2_X1 U703 ( .A1(n632), .A2(G2072), .ZN(n631) );
  XNOR2_X1 U704 ( .A(n631), .B(KEYINPUT27), .ZN(n634) );
  XOR2_X1 U705 ( .A(G1956), .B(KEYINPUT96), .Z(n956) );
  NOR2_X1 U706 ( .A1(n632), .A2(n956), .ZN(n633) );
  NOR2_X1 U707 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U708 ( .A1(n801), .A2(n637), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n640) );
  NOR2_X1 U710 ( .A1(n801), .A2(n637), .ZN(n638) );
  XOR2_X1 U711 ( .A(n638), .B(KEYINPUT28), .Z(n639) );
  NAND2_X1 U712 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n642), .B(n641), .ZN(n643) );
  AND2_X1 U714 ( .A1(n644), .A2(n643), .ZN(n655) );
  NAND2_X1 U715 ( .A1(n658), .A2(G8), .ZN(n645) );
  NOR2_X1 U716 ( .A1(n657), .A2(G1966), .ZN(n671) );
  NOR2_X1 U717 ( .A1(G2084), .A2(n658), .ZN(n667) );
  XNOR2_X1 U718 ( .A(n646), .B(KEYINPUT100), .ZN(n647) );
  NAND2_X1 U719 ( .A1(n647), .A2(G8), .ZN(n648) );
  XNOR2_X1 U720 ( .A(KEYINPUT30), .B(n648), .ZN(n649) );
  NOR2_X1 U721 ( .A1(G168), .A2(n649), .ZN(n652) );
  NOR2_X1 U722 ( .A1(G171), .A2(n650), .ZN(n651) );
  NOR2_X1 U723 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U724 ( .A(KEYINPUT31), .B(n653), .ZN(n654) );
  AND2_X1 U725 ( .A1(G286), .A2(G8), .ZN(n656) );
  NAND2_X1 U726 ( .A1(n669), .A2(n656), .ZN(n665) );
  INV_X1 U727 ( .A(G8), .ZN(n663) );
  NOR2_X1 U728 ( .A1(n682), .A2(G1971), .ZN(n660) );
  NOR2_X1 U729 ( .A1(G2090), .A2(n658), .ZN(n659) );
  NOR2_X1 U730 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U731 ( .A1(G303), .A2(n661), .ZN(n662) );
  OR2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n664) );
  AND2_X1 U733 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U734 ( .A(n666), .B(KEYINPUT32), .ZN(n673) );
  NAND2_X1 U735 ( .A1(G8), .A2(n667), .ZN(n668) );
  NAND2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n670) );
  OR2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U738 ( .A1(n673), .A2(n672), .ZN(n723) );
  NOR2_X1 U739 ( .A1(G288), .A2(G1976), .ZN(n674) );
  XOR2_X1 U740 ( .A(n674), .B(KEYINPUT101), .Z(n681) );
  NOR2_X1 U741 ( .A1(G303), .A2(G1971), .ZN(n675) );
  NOR2_X1 U742 ( .A1(n681), .A2(n675), .ZN(n924) );
  NAND2_X1 U743 ( .A1(n723), .A2(n924), .ZN(n676) );
  XNOR2_X1 U744 ( .A(n676), .B(KEYINPUT102), .ZN(n679) );
  NAND2_X1 U745 ( .A1(G1976), .A2(G288), .ZN(n915) );
  INV_X1 U746 ( .A(n915), .ZN(n677) );
  NOR2_X1 U747 ( .A1(n682), .A2(n677), .ZN(n678) );
  AND2_X1 U748 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U749 ( .A1(n680), .A2(KEYINPUT33), .ZN(n720) );
  AND2_X1 U750 ( .A1(n681), .A2(KEYINPUT33), .ZN(n683) );
  INV_X1 U751 ( .A(n682), .ZN(n727) );
  NAND2_X1 U752 ( .A1(n683), .A2(n727), .ZN(n716) );
  NOR2_X1 U753 ( .A1(n685), .A2(n684), .ZN(n748) );
  NAND2_X1 U754 ( .A1(n885), .A2(G104), .ZN(n686) );
  XNOR2_X1 U755 ( .A(n686), .B(KEYINPUT90), .ZN(n688) );
  NAND2_X1 U756 ( .A1(G140), .A2(n884), .ZN(n687) );
  NAND2_X1 U757 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U758 ( .A(KEYINPUT34), .B(n689), .ZN(n695) );
  NAND2_X1 U759 ( .A1(n880), .A2(G128), .ZN(n690) );
  XOR2_X1 U760 ( .A(KEYINPUT91), .B(n690), .Z(n692) );
  NAND2_X1 U761 ( .A1(n878), .A2(G116), .ZN(n691) );
  NAND2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U763 ( .A(n693), .B(KEYINPUT35), .Z(n694) );
  NOR2_X1 U764 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U765 ( .A(KEYINPUT36), .B(n696), .Z(n697) );
  XOR2_X1 U766 ( .A(KEYINPUT92), .B(n697), .Z(n893) );
  XNOR2_X1 U767 ( .A(G2067), .B(KEYINPUT37), .ZN(n745) );
  NOR2_X1 U768 ( .A1(n893), .A2(n745), .ZN(n1004) );
  NAND2_X1 U769 ( .A1(n748), .A2(n1004), .ZN(n743) );
  NAND2_X1 U770 ( .A1(G141), .A2(n884), .ZN(n699) );
  NAND2_X1 U771 ( .A1(G129), .A2(n880), .ZN(n698) );
  NAND2_X1 U772 ( .A1(n699), .A2(n698), .ZN(n702) );
  NAND2_X1 U773 ( .A1(n885), .A2(G105), .ZN(n700) );
  XOR2_X1 U774 ( .A(KEYINPUT38), .B(n700), .Z(n701) );
  NOR2_X1 U775 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U776 ( .A1(n878), .A2(G117), .ZN(n703) );
  NAND2_X1 U777 ( .A1(n704), .A2(n703), .ZN(n874) );
  AND2_X1 U778 ( .A1(n874), .A2(G1996), .ZN(n713) );
  NAND2_X1 U779 ( .A1(G131), .A2(n884), .ZN(n706) );
  NAND2_X1 U780 ( .A1(G95), .A2(n885), .ZN(n705) );
  NAND2_X1 U781 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U782 ( .A1(G119), .A2(n880), .ZN(n707) );
  XNOR2_X1 U783 ( .A(KEYINPUT93), .B(n707), .ZN(n708) );
  NOR2_X1 U784 ( .A1(n709), .A2(n708), .ZN(n711) );
  NAND2_X1 U785 ( .A1(n878), .A2(G107), .ZN(n710) );
  NAND2_X1 U786 ( .A1(n711), .A2(n710), .ZN(n875) );
  AND2_X1 U787 ( .A1(n875), .A2(G1991), .ZN(n712) );
  NOR2_X1 U788 ( .A1(n713), .A2(n712), .ZN(n988) );
  INV_X1 U789 ( .A(n748), .ZN(n714) );
  NOR2_X1 U790 ( .A1(n988), .A2(n714), .ZN(n740) );
  INV_X1 U791 ( .A(n740), .ZN(n715) );
  AND2_X1 U792 ( .A1(n743), .A2(n715), .ZN(n732) );
  AND2_X1 U793 ( .A1(n716), .A2(n732), .ZN(n718) );
  XNOR2_X1 U794 ( .A(G1981), .B(G305), .ZN(n910) );
  NOR2_X1 U795 ( .A1(n720), .A2(n719), .ZN(n734) );
  NOR2_X1 U796 ( .A1(G1981), .A2(G305), .ZN(n721) );
  XNOR2_X1 U797 ( .A(n721), .B(KEYINPUT24), .ZN(n722) );
  NAND2_X1 U798 ( .A1(n722), .A2(n727), .ZN(n730) );
  INV_X1 U799 ( .A(n723), .ZN(n726) );
  NAND2_X1 U800 ( .A1(G166), .A2(G8), .ZN(n724) );
  NOR2_X1 U801 ( .A1(G2090), .A2(n724), .ZN(n725) );
  NOR2_X1 U802 ( .A1(n726), .A2(n725), .ZN(n728) );
  OR2_X1 U803 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U804 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U805 ( .A1(n732), .A2(n731), .ZN(n733) );
  OR2_X1 U806 ( .A1(n734), .A2(n733), .ZN(n737) );
  XNOR2_X1 U807 ( .A(G1986), .B(G290), .ZN(n926) );
  NAND2_X1 U808 ( .A1(n926), .A2(n748), .ZN(n735) );
  XOR2_X1 U809 ( .A(KEYINPUT89), .B(n735), .Z(n736) );
  NAND2_X1 U810 ( .A1(n737), .A2(n736), .ZN(n750) );
  NOR2_X1 U811 ( .A1(G1996), .A2(n874), .ZN(n996) );
  NOR2_X1 U812 ( .A1(G1986), .A2(G290), .ZN(n738) );
  NOR2_X1 U813 ( .A1(G1991), .A2(n875), .ZN(n983) );
  NOR2_X1 U814 ( .A1(n738), .A2(n983), .ZN(n739) );
  NOR2_X1 U815 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U816 ( .A1(n996), .A2(n741), .ZN(n742) );
  XNOR2_X1 U817 ( .A(n742), .B(KEYINPUT39), .ZN(n744) );
  NAND2_X1 U818 ( .A1(n744), .A2(n743), .ZN(n746) );
  NAND2_X1 U819 ( .A1(n893), .A2(n745), .ZN(n987) );
  NAND2_X1 U820 ( .A1(n746), .A2(n987), .ZN(n747) );
  NAND2_X1 U821 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U822 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U823 ( .A(n751), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U824 ( .A(G2443), .B(KEYINPUT105), .Z(n753) );
  XNOR2_X1 U825 ( .A(G2451), .B(G2427), .ZN(n752) );
  XNOR2_X1 U826 ( .A(n753), .B(n752), .ZN(n754) );
  XOR2_X1 U827 ( .A(n754), .B(G2430), .Z(n756) );
  XNOR2_X1 U828 ( .A(G1348), .B(G1341), .ZN(n755) );
  XNOR2_X1 U829 ( .A(n756), .B(n755), .ZN(n760) );
  XOR2_X1 U830 ( .A(G2435), .B(KEYINPUT104), .Z(n758) );
  XNOR2_X1 U831 ( .A(G2438), .B(G2454), .ZN(n757) );
  XNOR2_X1 U832 ( .A(n758), .B(n757), .ZN(n759) );
  XOR2_X1 U833 ( .A(n760), .B(n759), .Z(n762) );
  XNOR2_X1 U834 ( .A(G2446), .B(KEYINPUT103), .ZN(n761) );
  XNOR2_X1 U835 ( .A(n762), .B(n761), .ZN(n763) );
  AND2_X1 U836 ( .A1(n763), .A2(G14), .ZN(G401) );
  INV_X1 U837 ( .A(n801), .ZN(G299) );
  INV_X1 U838 ( .A(G57), .ZN(G237) );
  INV_X1 U839 ( .A(G82), .ZN(G220) );
  NAND2_X1 U840 ( .A1(G94), .A2(G452), .ZN(n764) );
  XOR2_X1 U841 ( .A(KEYINPUT70), .B(n764), .Z(G173) );
  NAND2_X1 U842 ( .A1(G7), .A2(G661), .ZN(n765) );
  XNOR2_X1 U843 ( .A(n765), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U844 ( .A(G223), .ZN(n823) );
  NAND2_X1 U845 ( .A1(n823), .A2(G567), .ZN(n766) );
  XOR2_X1 U846 ( .A(KEYINPUT11), .B(n766), .Z(G234) );
  INV_X1 U847 ( .A(G860), .ZN(n771) );
  OR2_X1 U848 ( .A1(n920), .A2(n771), .ZN(G153) );
  INV_X1 U849 ( .A(G171), .ZN(G301) );
  NAND2_X1 U850 ( .A1(G868), .A2(G301), .ZN(n768) );
  OR2_X1 U851 ( .A1(n908), .A2(G868), .ZN(n767) );
  NAND2_X1 U852 ( .A1(n768), .A2(n767), .ZN(G284) );
  INV_X1 U853 ( .A(G868), .ZN(n806) );
  NOR2_X1 U854 ( .A1(G286), .A2(n806), .ZN(n770) );
  NOR2_X1 U855 ( .A1(G868), .A2(G299), .ZN(n769) );
  NOR2_X1 U856 ( .A1(n770), .A2(n769), .ZN(G297) );
  NAND2_X1 U857 ( .A1(n771), .A2(G559), .ZN(n772) );
  NAND2_X1 U858 ( .A1(n772), .A2(n908), .ZN(n773) );
  XNOR2_X1 U859 ( .A(n773), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U860 ( .A1(G868), .A2(n920), .ZN(n774) );
  XNOR2_X1 U861 ( .A(KEYINPUT80), .B(n774), .ZN(n777) );
  NAND2_X1 U862 ( .A1(G868), .A2(n908), .ZN(n775) );
  NOR2_X1 U863 ( .A1(G559), .A2(n775), .ZN(n776) );
  NOR2_X1 U864 ( .A1(n777), .A2(n776), .ZN(G282) );
  NAND2_X1 U865 ( .A1(n880), .A2(G123), .ZN(n778) );
  XNOR2_X1 U866 ( .A(n778), .B(KEYINPUT18), .ZN(n780) );
  NAND2_X1 U867 ( .A1(G99), .A2(n885), .ZN(n779) );
  NAND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n784) );
  NAND2_X1 U869 ( .A1(G135), .A2(n884), .ZN(n782) );
  NAND2_X1 U870 ( .A1(G111), .A2(n878), .ZN(n781) );
  NAND2_X1 U871 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n982) );
  XNOR2_X1 U873 ( .A(n982), .B(G2096), .ZN(n786) );
  INV_X1 U874 ( .A(G2100), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n786), .A2(n785), .ZN(G156) );
  NAND2_X1 U876 ( .A1(G559), .A2(n908), .ZN(n787) );
  XNOR2_X1 U877 ( .A(n787), .B(n920), .ZN(n830) );
  XNOR2_X1 U878 ( .A(G303), .B(G305), .ZN(n788) );
  XNOR2_X1 U879 ( .A(n788), .B(G288), .ZN(n800) );
  NAND2_X1 U880 ( .A1(G93), .A2(n789), .ZN(n792) );
  NAND2_X1 U881 ( .A1(G80), .A2(n790), .ZN(n791) );
  NAND2_X1 U882 ( .A1(n792), .A2(n791), .ZN(n798) );
  NAND2_X1 U883 ( .A1(G67), .A2(n793), .ZN(n796) );
  NAND2_X1 U884 ( .A1(G55), .A2(n794), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U886 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U887 ( .A(KEYINPUT81), .B(n799), .ZN(n831) );
  XNOR2_X1 U888 ( .A(n800), .B(n831), .ZN(n803) );
  XNOR2_X1 U889 ( .A(n801), .B(KEYINPUT19), .ZN(n802) );
  XNOR2_X1 U890 ( .A(n803), .B(n802), .ZN(n804) );
  XNOR2_X1 U891 ( .A(n804), .B(G290), .ZN(n896) );
  XNOR2_X1 U892 ( .A(n830), .B(n896), .ZN(n805) );
  NAND2_X1 U893 ( .A1(n805), .A2(G868), .ZN(n808) );
  NAND2_X1 U894 ( .A1(n806), .A2(n831), .ZN(n807) );
  NAND2_X1 U895 ( .A1(n808), .A2(n807), .ZN(G295) );
  XOR2_X1 U896 ( .A(KEYINPUT85), .B(KEYINPUT21), .Z(n812) );
  NAND2_X1 U897 ( .A1(G2078), .A2(G2084), .ZN(n809) );
  XOR2_X1 U898 ( .A(KEYINPUT20), .B(n809), .Z(n810) );
  NAND2_X1 U899 ( .A1(n810), .A2(G2090), .ZN(n811) );
  XNOR2_X1 U900 ( .A(n812), .B(n811), .ZN(n813) );
  NAND2_X1 U901 ( .A1(G2072), .A2(n813), .ZN(G158) );
  XNOR2_X1 U902 ( .A(KEYINPUT86), .B(G44), .ZN(n814) );
  XNOR2_X1 U903 ( .A(n814), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U904 ( .A(KEYINPUT71), .B(G132), .ZN(G219) );
  NOR2_X1 U905 ( .A1(G220), .A2(G219), .ZN(n815) );
  XOR2_X1 U906 ( .A(KEYINPUT22), .B(n815), .Z(n816) );
  NOR2_X1 U907 ( .A1(G218), .A2(n816), .ZN(n817) );
  NAND2_X1 U908 ( .A1(G96), .A2(n817), .ZN(n828) );
  NAND2_X1 U909 ( .A1(G2106), .A2(n828), .ZN(n821) );
  NAND2_X1 U910 ( .A1(G69), .A2(G120), .ZN(n818) );
  NOR2_X1 U911 ( .A1(G237), .A2(n818), .ZN(n819) );
  NAND2_X1 U912 ( .A1(G108), .A2(n819), .ZN(n829) );
  NAND2_X1 U913 ( .A1(G567), .A2(n829), .ZN(n820) );
  NAND2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n852) );
  NAND2_X1 U915 ( .A1(G483), .A2(G661), .ZN(n822) );
  NOR2_X1 U916 ( .A1(n852), .A2(n822), .ZN(n827) );
  NAND2_X1 U917 ( .A1(n827), .A2(G36), .ZN(G176) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n823), .ZN(G217) );
  NAND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n824) );
  XOR2_X1 U920 ( .A(KEYINPUT106), .B(n824), .Z(n825) );
  NAND2_X1 U921 ( .A1(G661), .A2(n825), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n826) );
  NAND2_X1 U923 ( .A1(n827), .A2(n826), .ZN(G188) );
  NOR2_X1 U924 ( .A1(n829), .A2(n828), .ZN(G325) );
  XNOR2_X1 U925 ( .A(KEYINPUT107), .B(G325), .ZN(G261) );
  INV_X1 U927 ( .A(G120), .ZN(G236) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  INV_X1 U929 ( .A(G69), .ZN(G235) );
  NOR2_X1 U930 ( .A1(n830), .A2(G860), .ZN(n832) );
  XOR2_X1 U931 ( .A(n832), .B(n831), .Z(G145) );
  XNOR2_X1 U932 ( .A(G1996), .B(G2474), .ZN(n842) );
  XOR2_X1 U933 ( .A(G1976), .B(G1961), .Z(n834) );
  XNOR2_X1 U934 ( .A(G1991), .B(G1956), .ZN(n833) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U936 ( .A(G1971), .B(G1966), .Z(n836) );
  XNOR2_X1 U937 ( .A(G1986), .B(G1981), .ZN(n835) );
  XNOR2_X1 U938 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U939 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U940 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(G229) );
  XOR2_X1 U943 ( .A(G2678), .B(G2084), .Z(n844) );
  XNOR2_X1 U944 ( .A(G2072), .B(G2078), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U946 ( .A(n845), .B(G2100), .Z(n847) );
  XNOR2_X1 U947 ( .A(G2067), .B(G2090), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U949 ( .A(G2096), .B(KEYINPUT109), .Z(n849) );
  XNOR2_X1 U950 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U952 ( .A(n851), .B(n850), .Z(G227) );
  XOR2_X1 U953 ( .A(KEYINPUT108), .B(n852), .Z(G319) );
  NAND2_X1 U954 ( .A1(G136), .A2(n884), .ZN(n854) );
  NAND2_X1 U955 ( .A1(G100), .A2(n885), .ZN(n853) );
  NAND2_X1 U956 ( .A1(n854), .A2(n853), .ZN(n860) );
  NAND2_X1 U957 ( .A1(G124), .A2(n880), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n855), .B(KEYINPUT44), .ZN(n858) );
  NAND2_X1 U959 ( .A1(G112), .A2(n878), .ZN(n856) );
  XOR2_X1 U960 ( .A(KEYINPUT111), .B(n856), .Z(n857) );
  NAND2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U962 ( .A1(n860), .A2(n859), .ZN(G162) );
  XOR2_X1 U963 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n862) );
  XNOR2_X1 U964 ( .A(n982), .B(KEYINPUT114), .ZN(n861) );
  XNOR2_X1 U965 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U966 ( .A(n863), .B(G162), .Z(n865) );
  XNOR2_X1 U967 ( .A(G164), .B(G160), .ZN(n864) );
  XNOR2_X1 U968 ( .A(n865), .B(n864), .ZN(n873) );
  NAND2_X1 U969 ( .A1(G139), .A2(n884), .ZN(n867) );
  NAND2_X1 U970 ( .A1(G103), .A2(n885), .ZN(n866) );
  NAND2_X1 U971 ( .A1(n867), .A2(n866), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G127), .A2(n880), .ZN(n869) );
  NAND2_X1 U973 ( .A1(G115), .A2(n878), .ZN(n868) );
  NAND2_X1 U974 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U975 ( .A(KEYINPUT47), .B(n870), .Z(n871) );
  NOR2_X1 U976 ( .A1(n872), .A2(n871), .ZN(n991) );
  XOR2_X1 U977 ( .A(n873), .B(n991), .Z(n877) );
  XNOR2_X1 U978 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U979 ( .A(n877), .B(n876), .ZN(n892) );
  NAND2_X1 U980 ( .A1(n878), .A2(G118), .ZN(n879) );
  XNOR2_X1 U981 ( .A(n879), .B(KEYINPUT112), .ZN(n882) );
  NAND2_X1 U982 ( .A1(G130), .A2(n880), .ZN(n881) );
  NAND2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U984 ( .A(KEYINPUT113), .B(n883), .Z(n890) );
  NAND2_X1 U985 ( .A1(G142), .A2(n884), .ZN(n887) );
  NAND2_X1 U986 ( .A1(G106), .A2(n885), .ZN(n886) );
  NAND2_X1 U987 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U988 ( .A(n888), .B(KEYINPUT45), .Z(n889) );
  NOR2_X1 U989 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U990 ( .A(n892), .B(n891), .Z(n894) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U992 ( .A1(G37), .A2(n895), .ZN(G395) );
  XNOR2_X1 U993 ( .A(n896), .B(KEYINPUT115), .ZN(n898) );
  XNOR2_X1 U994 ( .A(n920), .B(G171), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n898), .B(n897), .ZN(n900) );
  XNOR2_X1 U996 ( .A(G286), .B(n908), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U998 ( .A1(G37), .A2(n901), .ZN(G397) );
  NOR2_X1 U999 ( .A1(G229), .A2(G227), .ZN(n902) );
  XOR2_X1 U1000 ( .A(KEYINPUT49), .B(n902), .Z(n903) );
  NAND2_X1 U1001 ( .A1(n903), .A2(G319), .ZN(n904) );
  NOR2_X1 U1002 ( .A1(G401), .A2(n904), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(KEYINPUT116), .B(n905), .ZN(n907) );
  NOR2_X1 U1004 ( .A1(G395), .A2(G397), .ZN(n906) );
  NAND2_X1 U1005 ( .A1(n907), .A2(n906), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1008 ( .A(KEYINPUT56), .B(G16), .ZN(n930) );
  XOR2_X1 U1009 ( .A(G1348), .B(n908), .Z(n913) );
  XOR2_X1 U1010 ( .A(G1966), .B(G168), .Z(n909) );
  NOR2_X1 U1011 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1012 ( .A(KEYINPUT57), .B(n911), .ZN(n912) );
  NOR2_X1 U1013 ( .A1(n913), .A2(n912), .ZN(n928) );
  XNOR2_X1 U1014 ( .A(G171), .B(G1961), .ZN(n919) );
  NAND2_X1 U1015 ( .A1(G303), .A2(G1971), .ZN(n914) );
  NAND2_X1 U1016 ( .A1(n915), .A2(n914), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(G1956), .B(G299), .ZN(n916) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(G1341), .B(n920), .ZN(n921) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1025 ( .A1(n930), .A2(n929), .ZN(n1014) );
  XNOR2_X1 U1026 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n1006) );
  XNOR2_X1 U1027 ( .A(n1006), .B(KEYINPUT123), .ZN(n952) );
  XNOR2_X1 U1028 ( .A(G2090), .B(G35), .ZN(n946) );
  XNOR2_X1 U1029 ( .A(G2067), .B(G26), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(G33), .B(G2072), .ZN(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n940) );
  XOR2_X1 U1032 ( .A(G1991), .B(G25), .Z(n933) );
  NAND2_X1 U1033 ( .A1(n933), .A2(G28), .ZN(n934) );
  XNOR2_X1 U1034 ( .A(n934), .B(KEYINPUT120), .ZN(n938) );
  XNOR2_X1 U1035 ( .A(n935), .B(G32), .ZN(n936) );
  XNOR2_X1 U1036 ( .A(KEYINPUT121), .B(n936), .ZN(n937) );
  NOR2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n943) );
  XOR2_X1 U1039 ( .A(G27), .B(n941), .Z(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(KEYINPUT53), .B(n944), .ZN(n945) );
  NOR2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n950) );
  XOR2_X1 U1043 ( .A(G34), .B(KEYINPUT122), .Z(n948) );
  XNOR2_X1 U1044 ( .A(G2084), .B(KEYINPUT54), .ZN(n947) );
  XNOR2_X1 U1045 ( .A(n948), .B(n947), .ZN(n949) );
  NAND2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(n952), .B(n951), .ZN(n953) );
  OR2_X1 U1048 ( .A1(G29), .A2(n953), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(G11), .A2(n954), .ZN(n1012) );
  XOR2_X1 U1050 ( .A(G1348), .B(KEYINPUT59), .Z(n955) );
  XNOR2_X1 U1051 ( .A(G4), .B(n955), .ZN(n963) );
  XOR2_X1 U1052 ( .A(G1981), .B(G6), .Z(n958) );
  XNOR2_X1 U1053 ( .A(n956), .B(G20), .ZN(n957) );
  NAND2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(G19), .B(G1341), .ZN(n959) );
  NOR2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1057 ( .A(KEYINPUT124), .B(n961), .Z(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(KEYINPUT60), .B(n964), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(n965), .B(G5), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n978) );
  XOR2_X1 U1062 ( .A(G1966), .B(G21), .Z(n976) );
  XOR2_X1 U1063 ( .A(G1971), .B(G22), .Z(n970) );
  XOR2_X1 U1064 ( .A(G24), .B(KEYINPUT126), .Z(n968) );
  XNOR2_X1 U1065 ( .A(n968), .B(G1986), .ZN(n969) );
  NAND2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n973) );
  XOR2_X1 U1067 ( .A(KEYINPUT125), .B(G1976), .Z(n971) );
  XNOR2_X1 U1068 ( .A(G23), .B(n971), .ZN(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(n974), .B(KEYINPUT58), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1073 ( .A(KEYINPUT61), .B(n979), .Z(n980) );
  NOR2_X1 U1074 ( .A1(G16), .A2(n980), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(KEYINPUT127), .B(n981), .ZN(n1010) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n986) );
  XOR2_X1 U1077 ( .A(G160), .B(G2084), .Z(n984) );
  XNOR2_X1 U1078 ( .A(KEYINPUT117), .B(n984), .ZN(n985) );
  NAND2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n990) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n1002) );
  XOR2_X1 U1082 ( .A(G2072), .B(n991), .Z(n993) );
  XOR2_X1 U1083 ( .A(G164), .B(G2078), .Z(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1085 ( .A(KEYINPUT50), .B(n994), .Z(n1000) );
  XOR2_X1 U1086 ( .A(G2090), .B(G162), .Z(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1088 ( .A(KEYINPUT118), .B(n997), .Z(n998) );
  XOR2_X1 U1089 ( .A(KEYINPUT51), .B(n998), .Z(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(KEYINPUT52), .B(n1005), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(G29), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1098 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1099 ( .A(KEYINPUT62), .B(n1015), .Z(G311) );
  INV_X1 U1100 ( .A(G311), .ZN(G150) );
endmodule

