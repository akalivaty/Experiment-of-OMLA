//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1222, new_n1223, new_n1224, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT65), .Z(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT66), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n208), .B1(new_n210), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT1), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n208), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT0), .Z(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n203), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n216), .B(new_n219), .C1(new_n222), .C2(new_n224), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G87), .B(G97), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT68), .ZN(new_n235));
  XOR2_X1   g0035(.A(G107), .B(G116), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G68), .B(G77), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n201), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT67), .B(G50), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n237), .B(new_n241), .Z(G351));
  NAND3_X1  g0042(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(new_n220), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT8), .B(G58), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n221), .A2(G33), .ZN(new_n246));
  INV_X1    g0046(.A(G150), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  OAI22_X1  g0049(.A1(new_n245), .A2(new_n246), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n203), .A2(G50), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(new_n221), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n244), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G13), .ZN(new_n254));
  NOR3_X1   g0054(.A1(new_n254), .A2(new_n221), .A3(G1), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(new_n244), .ZN(new_n256));
  INV_X1    g0056(.A(G50), .ZN(new_n257));
  OAI21_X1  g0057(.A(KEYINPUT71), .B1(new_n221), .B2(G1), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT71), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(new_n260), .A3(G20), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n257), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n256), .A2(new_n262), .B1(new_n257), .B2(new_n255), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n253), .A2(new_n263), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n264), .A2(KEYINPUT9), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(KEYINPUT9), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT74), .ZN(new_n268));
  AOI21_X1  g0068(.A(KEYINPUT10), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n265), .A2(KEYINPUT74), .A3(new_n266), .ZN(new_n270));
  AND2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G33), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT70), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n272), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT70), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(G222), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G77), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(G223), .ZN(new_n286));
  OAI221_X1 g0086(.A(new_n283), .B1(new_n284), .B2(new_n281), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  AND2_X1   g0087(.A1(G1), .A2(G13), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G41), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G274), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(new_n288), .B2(new_n289), .ZN(new_n294));
  INV_X1    g0094(.A(G41), .ZN(new_n295));
  INV_X1    g0095(.A(G45), .ZN(new_n296));
  AOI21_X1  g0096(.A(G1), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n297), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n290), .ZN(new_n300));
  INV_X1    g0100(.A(G226), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT69), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n292), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G200), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n292), .A2(G190), .A3(new_n303), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(new_n306), .A3(new_n267), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n271), .A2(new_n307), .B1(new_n308), .B2(KEYINPUT10), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n304), .A2(new_n310), .B1(new_n253), .B2(new_n263), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(G179), .B2(new_n304), .ZN(new_n312));
  OAI22_X1  g0112(.A1(new_n245), .A2(new_n249), .B1(new_n221), .B2(new_n284), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT15), .B(G87), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(new_n246), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n244), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n258), .A2(new_n261), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n256), .A2(G77), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n255), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n316), .B(new_n318), .C1(G77), .C2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G244), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n298), .B1(new_n300), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n281), .A2(G232), .A3(new_n282), .ZN(new_n323));
  AND3_X1   g0123(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n279), .B1(new_n277), .B2(new_n278), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G107), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT72), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT72), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G107), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G238), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n323), .B(new_n332), .C1(new_n285), .C2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n322), .B1(new_n334), .B2(new_n291), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n320), .B1(new_n336), .B2(G200), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n335), .A2(KEYINPUT73), .A3(G190), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT73), .B1(new_n335), .B2(G190), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n336), .A2(G179), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n320), .B1(new_n335), .B2(G169), .ZN(new_n342));
  OR2_X1    g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n312), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n309), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G190), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT75), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n294), .A2(new_n347), .A3(new_n297), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n347), .B1(new_n294), .B2(new_n297), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n348), .A2(new_n349), .B1(new_n333), .B2(new_n300), .ZN(new_n350));
  OAI211_X1 g0150(.A(G226), .B(new_n282), .C1(new_n324), .C2(new_n325), .ZN(new_n351));
  OAI211_X1 g0151(.A(G232), .B(G1698), .C1(new_n324), .C2(new_n325), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G33), .A2(G97), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n350), .B1(new_n354), .B2(new_n291), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT13), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n346), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT76), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT13), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  AOI211_X1 g0159(.A(KEYINPUT76), .B(new_n350), .C1(new_n354), .C2(new_n291), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n355), .A2(new_n356), .ZN(new_n362));
  AOI211_X1 g0162(.A(KEYINPUT13), .B(new_n350), .C1(new_n354), .C2(new_n291), .ZN(new_n363));
  OAI21_X1  g0163(.A(G200), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n248), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n284), .B2(new_n246), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n244), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT11), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n255), .A2(new_n202), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n370), .B(KEYINPUT12), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n366), .A2(KEYINPUT11), .A3(new_n244), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n256), .A2(G68), .A3(new_n317), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n369), .A2(new_n371), .A3(new_n372), .A4(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n361), .A2(new_n364), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT77), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n361), .A2(new_n364), .A3(KEYINPUT77), .A4(new_n375), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n345), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n245), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n256), .A2(new_n382), .A3(new_n317), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n245), .A2(new_n255), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g0185(.A(new_n385), .B(KEYINPUT80), .ZN(new_n386));
  XNOR2_X1  g0186(.A(G58), .B(G68), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(G20), .B1(G159), .B2(new_n248), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n272), .A2(KEYINPUT78), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT78), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT3), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(new_n391), .A3(G33), .ZN(new_n392));
  AOI21_X1  g0192(.A(G20), .B1(new_n392), .B2(new_n277), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n202), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n273), .B1(new_n396), .B2(G33), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT7), .B1(new_n397), .B2(G20), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n395), .A2(KEYINPUT79), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT79), .B1(new_n395), .B2(new_n398), .ZN(new_n400));
  OAI211_X1 g0200(.A(KEYINPUT16), .B(new_n388), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n244), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n276), .A2(new_n221), .A3(new_n280), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n278), .B1(new_n396), .B2(G33), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n394), .A2(G20), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n403), .A2(new_n394), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n388), .B1(new_n406), .B2(new_n202), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT16), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n402), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n386), .B1(new_n401), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT82), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G87), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n412), .B(KEYINPUT81), .ZN(new_n413));
  NOR2_X1   g0213(.A1(G223), .A2(G1698), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n301), .B2(G1698), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n413), .B1(new_n397), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n411), .B1(new_n416), .B2(new_n290), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n392), .A3(new_n277), .ZN(new_n418));
  INV_X1    g0218(.A(new_n413), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(KEYINPUT82), .A3(new_n291), .ZN(new_n421));
  INV_X1    g0221(.A(G232), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n298), .B1(new_n300), .B2(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(G179), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n417), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT83), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n416), .A2(new_n290), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n310), .B1(new_n428), .B2(new_n423), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n417), .A2(KEYINPUT83), .A3(new_n421), .A4(new_n424), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n427), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n410), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n432), .B(KEYINPUT18), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n423), .A2(G190), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n417), .A2(new_n421), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(G200), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n428), .B2(new_n423), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n410), .A2(new_n438), .ZN(new_n439));
  AND2_X1   g0239(.A1(KEYINPUT84), .A2(KEYINPUT17), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(KEYINPUT84), .A2(KEYINPUT17), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n439), .B1(new_n442), .B2(new_n440), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n433), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT85), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n359), .A2(new_n360), .ZN(new_n448));
  INV_X1    g0248(.A(G179), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n363), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n354), .A2(new_n291), .ZN(new_n452));
  INV_X1    g0252(.A(new_n350), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT13), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n355), .A2(new_n356), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(KEYINPUT14), .B1(new_n457), .B2(G169), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT14), .ZN(new_n459));
  AOI211_X1 g0259(.A(new_n459), .B(new_n310), .C1(new_n455), .C2(new_n456), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n451), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n374), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n381), .A2(new_n446), .A3(new_n447), .A4(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n345), .A2(new_n462), .A3(new_n380), .ZN(new_n464));
  OAI21_X1  g0264(.A(KEYINPUT85), .B1(new_n464), .B2(new_n445), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(G250), .A2(G1698), .ZN(new_n467));
  INV_X1    g0267(.A(G257), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n467), .B1(new_n468), .B2(G1698), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n469), .A2(new_n392), .A3(new_n277), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G294), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n290), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  XNOR2_X1  g0273(.A(KEYINPUT5), .B(G41), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n296), .A2(G1), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n290), .ZN(new_n477));
  INV_X1    g0277(.A(G264), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n294), .A2(new_n475), .A3(new_n474), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n473), .A2(new_n480), .A3(new_n449), .A4(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n481), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n472), .A2(new_n479), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n482), .B1(new_n484), .B2(G169), .ZN(new_n485));
  OAI21_X1  g0285(.A(KEYINPUT23), .B1(new_n331), .B2(new_n221), .ZN(new_n486));
  INV_X1    g0286(.A(G116), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n246), .A2(new_n487), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n221), .A2(KEYINPUT23), .A3(G107), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(G87), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n492), .A2(KEYINPUT22), .A3(G20), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n281), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n392), .A2(new_n221), .A3(G87), .A4(new_n277), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT22), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n491), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT24), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n281), .A2(new_n493), .B1(new_n495), .B2(KEYINPUT22), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n500), .A2(KEYINPUT24), .A3(new_n491), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n244), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n260), .A2(G33), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n256), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n504), .A2(new_n327), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n254), .A2(G1), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(G20), .A3(new_n327), .ZN(new_n507));
  XNOR2_X1  g0307(.A(new_n507), .B(KEYINPUT25), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n485), .B1(new_n502), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n497), .A2(new_n498), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT24), .B1(new_n500), .B2(new_n491), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n402), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n509), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n472), .A2(new_n479), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n481), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT90), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n518), .A3(new_n436), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT90), .B1(new_n484), .B2(G200), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n484), .A2(new_n346), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n510), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n256), .A2(G116), .A3(new_n503), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n255), .A2(new_n487), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n243), .A2(new_n220), .B1(G20), .B2(new_n487), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G283), .ZN(new_n527));
  INV_X1    g0327(.A(G97), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n527), .B(new_n221), .C1(G33), .C2(new_n528), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n526), .A2(KEYINPUT20), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT20), .B1(new_n526), .B2(new_n529), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n524), .B(new_n525), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  XOR2_X1   g0332(.A(KEYINPUT88), .B(G303), .Z(new_n533));
  NAND3_X1  g0333(.A1(new_n276), .A2(new_n280), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(G257), .A2(G1698), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n478), .B2(G1698), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(new_n392), .A3(new_n277), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n290), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(G270), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n481), .B1(new_n477), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n532), .B(G169), .C1(new_n538), .C2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(KEYINPUT21), .B1(new_n542), .B2(KEYINPUT89), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n538), .A2(new_n540), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n544), .A2(G179), .A3(new_n532), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT89), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT21), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n541), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n543), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n544), .A2(new_n436), .ZN(new_n550));
  AOI211_X1 g0350(.A(new_n532), .B(new_n550), .C1(G190), .C2(new_n544), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n314), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(new_n319), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n504), .A2(new_n314), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n397), .A2(new_n221), .A3(G68), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n246), .B2(new_n528), .ZN(new_n558));
  OR2_X1    g0358(.A1(new_n558), .A2(KEYINPUT87), .ZN(new_n559));
  XNOR2_X1  g0359(.A(KEYINPUT72), .B(G107), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(new_n492), .A3(new_n528), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n221), .B1(new_n353), .B2(new_n557), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n558), .A2(KEYINPUT87), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n556), .A2(new_n559), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  AOI211_X1 g0365(.A(new_n554), .B(new_n555), .C1(new_n565), .C2(new_n244), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(G238), .A2(G1698), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n568), .B1(new_n321), .B2(G1698), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(new_n392), .A3(new_n277), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G33), .A2(G116), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n290), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n290), .B(G250), .C1(G1), .C2(new_n296), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n294), .A2(new_n475), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n449), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n310), .B1(new_n572), .B2(new_n575), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n504), .A2(new_n492), .ZN(new_n581));
  AOI211_X1 g0381(.A(new_n554), .B(new_n581), .C1(new_n565), .C2(new_n244), .ZN(new_n582));
  INV_X1    g0382(.A(new_n575), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n570), .A2(new_n571), .ZN(new_n584));
  OAI211_X1 g0384(.A(G190), .B(new_n583), .C1(new_n584), .C2(new_n290), .ZN(new_n585));
  OAI21_X1  g0385(.A(G200), .B1(new_n572), .B2(new_n575), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n567), .A2(new_n580), .B1(new_n582), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n481), .B1(new_n477), .B2(new_n468), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n321), .A2(G1698), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n392), .A2(new_n277), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT4), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n282), .A2(KEYINPUT4), .A3(G244), .ZN(new_n594));
  INV_X1    g0394(.A(G250), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n594), .B1(new_n595), .B2(new_n282), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n324), .B2(new_n325), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n593), .A2(new_n527), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n589), .B1(new_n598), .B2(new_n291), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G190), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n255), .A2(new_n528), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n504), .B2(new_n528), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n327), .A2(KEYINPUT6), .A3(G97), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n528), .A2(new_n327), .ZN(new_n604));
  NOR2_X1   g0404(.A1(G97), .A2(G107), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n603), .B1(new_n606), .B2(KEYINPUT6), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n607), .A2(G20), .B1(G77), .B2(new_n248), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n406), .B2(new_n560), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n602), .B1(new_n609), .B2(new_n244), .ZN(new_n610));
  OAI21_X1  g0410(.A(G200), .B1(new_n599), .B2(KEYINPUT86), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT86), .ZN(new_n612));
  AOI211_X1 g0412(.A(new_n612), .B(new_n589), .C1(new_n598), .C2(new_n291), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n600), .B(new_n610), .C1(new_n611), .C2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n609), .A2(new_n244), .ZN(new_n615));
  INV_X1    g0415(.A(new_n602), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n598), .A2(new_n291), .ZN(new_n618));
  INV_X1    g0418(.A(new_n589), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n310), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n599), .A2(new_n449), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n617), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n588), .A2(new_n614), .A3(new_n623), .ZN(new_n624));
  AND4_X1   g0424(.A1(new_n466), .A2(new_n523), .A3(new_n552), .A4(new_n624), .ZN(G372));
  NOR2_X1   g0425(.A1(new_n566), .A2(new_n579), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n617), .A2(new_n621), .A3(new_n622), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n627), .A2(new_n588), .A3(KEYINPUT26), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n565), .A2(new_n244), .ZN(new_n630));
  INV_X1    g0430(.A(new_n554), .ZN(new_n631));
  INV_X1    g0431(.A(new_n581), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n585), .A2(new_n586), .ZN(new_n634));
  OAI22_X1  g0434(.A1(new_n566), .A2(new_n579), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n629), .B1(new_n623), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n626), .B1(new_n628), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n614), .A2(new_n623), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n515), .A2(new_n522), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n639), .B(new_n588), .C1(new_n549), .C2(new_n510), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n637), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n466), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n312), .ZN(new_n643));
  INV_X1    g0443(.A(new_n444), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n341), .A2(new_n342), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n461), .A2(new_n374), .B1(new_n376), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n433), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT91), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n309), .B(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n643), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n642), .A2(new_n650), .ZN(G369));
  NAND2_X1  g0451(.A1(new_n506), .A2(new_n221), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(G213), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(G343), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n657), .A2(new_n532), .ZN(new_n658));
  MUX2_X1   g0458(.A(new_n552), .B(new_n549), .S(new_n658), .Z(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  INV_X1    g0460(.A(new_n657), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n523), .B1(new_n515), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n517), .A2(new_n310), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n482), .B(new_n663), .C1(new_n513), .C2(new_n514), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n662), .B1(new_n664), .B2(new_n661), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n549), .A2(new_n661), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n668), .A2(new_n523), .B1(new_n510), .B2(new_n661), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n666), .A2(new_n669), .ZN(G399));
  INV_X1    g0470(.A(new_n217), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G41), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n224), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n561), .A2(G116), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G1), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n673), .B1(new_n672), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n641), .A2(new_n661), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT29), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n614), .A2(new_n623), .A3(KEYINPUT93), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(KEYINPUT93), .B1(new_n614), .B2(new_n623), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n640), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n628), .A2(new_n636), .ZN(new_n684));
  INV_X1    g0484(.A(new_n626), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n661), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT29), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n679), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n599), .A2(new_n516), .A3(new_n576), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n544), .A2(G179), .ZN(new_n692));
  OAI21_X1  g0492(.A(KEYINPUT92), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT30), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT30), .ZN(new_n695));
  OAI211_X1 g0495(.A(KEYINPUT92), .B(new_n695), .C1(new_n691), .C2(new_n692), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n544), .A2(new_n576), .A3(G179), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(new_n517), .A3(new_n620), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n694), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n657), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT31), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n624), .A2(new_n523), .A3(new_n552), .A4(new_n661), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n699), .A2(KEYINPUT31), .A3(new_n657), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(G330), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n690), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n677), .B1(new_n711), .B2(G1), .ZN(G364));
  NOR2_X1   g0512(.A1(new_n659), .A2(G330), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n254), .A2(G20), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n260), .B1(new_n714), .B2(G45), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n672), .A2(new_n716), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n660), .A2(new_n713), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT94), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n221), .A2(G179), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G190), .A2(G200), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G159), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT32), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n346), .A2(G179), .A3(G200), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n221), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n720), .A2(G190), .A3(G200), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n727), .A2(new_n528), .B1(new_n728), .B2(new_n492), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n221), .A2(new_n449), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n732), .A2(new_n346), .A3(G200), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n732), .A2(new_n436), .A3(G190), .ZN(new_n734));
  AOI22_X1  g0534(.A1(G58), .A2(new_n733), .B1(new_n734), .B2(G68), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n731), .A2(new_n721), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n735), .B1(new_n284), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n731), .A2(G190), .A3(G200), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(KEYINPUT96), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n738), .A2(KEYINPUT96), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n257), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n720), .A2(new_n346), .A3(G200), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n327), .ZN(new_n745));
  NOR4_X1   g0545(.A1(new_n737), .A2(new_n743), .A3(new_n326), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(KEYINPUT33), .B(G317), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n734), .A2(new_n747), .B1(G329), .B2(new_n723), .ZN(new_n748));
  INV_X1    g0548(.A(G311), .ZN(new_n749));
  INV_X1    g0549(.A(G322), .ZN(new_n750));
  INV_X1    g0550(.A(new_n733), .ZN(new_n751));
  OAI221_X1 g0551(.A(new_n748), .B1(new_n749), .B2(new_n736), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n742), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n752), .B1(G326), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G294), .ZN(new_n755));
  INV_X1    g0555(.A(G283), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n727), .A2(new_n755), .B1(new_n744), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n728), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n281), .B(new_n757), .C1(G303), .C2(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n730), .A2(new_n746), .B1(new_n754), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n220), .B1(G20), .B2(new_n310), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n717), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n761), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n671), .A2(new_n397), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n770), .B1(new_n296), .B2(new_n224), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n241), .A2(G45), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT95), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n217), .A2(new_n281), .A3(G355), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(G116), .B2(new_n217), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n771), .A2(new_n772), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n775), .A2(new_n773), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n768), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n763), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n766), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(new_n659), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n719), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT97), .ZN(G396));
  NOR2_X1   g0583(.A1(new_n343), .A2(new_n657), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n320), .A2(new_n657), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n645), .B1(new_n340), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n678), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n784), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n641), .A2(new_n661), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n717), .B1(new_n790), .B2(new_n709), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n709), .B2(new_n790), .ZN(new_n792));
  INV_X1    g0592(.A(new_n736), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n734), .A2(G150), .B1(G159), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G143), .ZN(new_n795));
  INV_X1    g0595(.A(G137), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n794), .B1(new_n795), .B2(new_n751), .C1(new_n742), .C2(new_n796), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT34), .Z(new_n798));
  INV_X1    g0598(.A(G132), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n397), .B1(new_n799), .B2(new_n722), .ZN(new_n800));
  INV_X1    g0600(.A(new_n744), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n758), .A2(G50), .B1(new_n801), .B2(G68), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n201), .B2(new_n727), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n798), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n758), .A2(G107), .ZN(new_n805));
  XOR2_X1   g0605(.A(KEYINPUT98), .B(G283), .Z(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n734), .A2(new_n807), .B1(new_n793), .B2(G116), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(KEYINPUT99), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n751), .A2(new_n755), .B1(new_n722), .B2(new_n749), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n809), .A2(new_n810), .A3(new_n281), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n753), .A2(G303), .B1(KEYINPUT99), .B2(new_n808), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n744), .A2(new_n492), .ZN(new_n813));
  INV_X1    g0613(.A(new_n727), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n813), .B1(G97), .B2(new_n814), .ZN(new_n815));
  AND4_X1   g0615(.A1(new_n805), .A2(new_n811), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n761), .B1(new_n804), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n717), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n761), .A2(new_n764), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n818), .B1(new_n284), .B2(new_n819), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n817), .B(new_n820), .C1(new_n788), .C2(new_n765), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n792), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G384));
  OR2_X1    g0623(.A1(new_n607), .A2(KEYINPUT35), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n607), .A2(KEYINPUT35), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n824), .A2(G116), .A3(new_n222), .A4(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT36), .Z(new_n827));
  OAI211_X1 g0627(.A(new_n224), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n257), .A2(G68), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n260), .B(G13), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n705), .A2(new_n788), .ZN(new_n832));
  OAI21_X1  g0632(.A(G169), .B1(new_n362), .B2(new_n363), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n459), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n457), .A2(KEYINPUT14), .A3(G169), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n834), .A2(new_n835), .B1(new_n448), .B2(new_n450), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n374), .B1(new_n457), .B2(G200), .ZN(new_n837));
  AOI21_X1  g0637(.A(KEYINPUT77), .B1(new_n837), .B2(new_n361), .ZN(new_n838));
  INV_X1    g0638(.A(new_n379), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n374), .A2(new_n657), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n841), .B(KEYINPUT100), .Z(new_n844));
  OAI211_X1 g0644(.A(new_n376), .B(new_n844), .C1(new_n836), .C2(new_n375), .ZN(new_n845));
  AOI21_X1  g0645(.A(KEYINPUT101), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n841), .B1(new_n380), .B2(new_n836), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT101), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n376), .A2(new_n844), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n461), .B2(new_n374), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n832), .B1(new_n846), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT104), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT40), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n401), .A2(new_n409), .ZN(new_n856));
  INV_X1    g0656(.A(new_n386), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n431), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n655), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n860), .A2(new_n862), .A3(new_n863), .A4(new_n439), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT102), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI221_X4 g0666(.A(new_n386), .B1(new_n437), .B2(new_n435), .C1(new_n401), .C2(new_n409), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n432), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n868), .A2(KEYINPUT102), .A3(new_n863), .A4(new_n862), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n385), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n401), .A2(new_n244), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n392), .A2(new_n277), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n873), .A2(new_n394), .A3(new_n221), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n398), .A2(G68), .A3(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT79), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n395), .A2(KEYINPUT79), .A3(new_n398), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT16), .B1(new_n879), .B2(new_n388), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n871), .B1(new_n872), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n861), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n859), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(new_n883), .A3(new_n439), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n870), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n882), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n445), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n886), .A2(KEYINPUT38), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n863), .B1(new_n868), .B2(new_n862), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n866), .B2(new_n869), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n862), .B1(new_n433), .B2(new_n444), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n890), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n855), .B1(new_n889), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n705), .A2(new_n788), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n848), .B1(new_n847), .B2(new_n850), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n461), .B1(new_n378), .B2(new_n379), .ZN(new_n898));
  OAI211_X1 g0698(.A(KEYINPUT101), .B(new_n845), .C1(new_n898), .C2(new_n841), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n896), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(KEYINPUT104), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n854), .A2(new_n895), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT38), .B1(new_n886), .B2(new_n888), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n866), .A2(new_n869), .B1(KEYINPUT37), .B2(new_n884), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n882), .B1(new_n433), .B2(new_n444), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n904), .A2(new_n905), .A3(new_n890), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n900), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n855), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n466), .A2(new_n705), .ZN(new_n911));
  OAI21_X1  g0711(.A(G330), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n910), .B2(new_n911), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n466), .A2(new_n689), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n650), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT103), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n462), .A2(new_n657), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n890), .B1(new_n904), .B2(new_n905), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n889), .A2(new_n918), .A3(KEYINPUT39), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n889), .A2(new_n894), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n917), .B(new_n919), .C1(new_n920), .C2(KEYINPUT39), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n897), .A2(new_n899), .ZN(new_n922));
  INV_X1    g0722(.A(new_n784), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n789), .A2(new_n923), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n889), .A2(new_n918), .ZN(new_n926));
  INV_X1    g0726(.A(new_n433), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n925), .A2(new_n926), .B1(new_n927), .B2(new_n655), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n921), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n916), .B(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n913), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n913), .A2(new_n930), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT105), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n931), .B1(new_n260), .B2(new_n714), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n932), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n935), .A2(KEYINPUT105), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n831), .B1(new_n934), .B2(new_n936), .ZN(G367));
  INV_X1    g0737(.A(KEYINPUT93), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n638), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n939), .B(new_n680), .C1(new_n610), .C2(new_n661), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n627), .A2(new_n657), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(new_n523), .A3(new_n668), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n943), .A2(KEYINPUT42), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n623), .B1(new_n940), .B2(new_n664), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n943), .A2(KEYINPUT42), .B1(new_n661), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n947), .A2(KEYINPUT106), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n633), .A2(new_n657), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n588), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n685), .B2(new_n949), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n947), .A2(KEYINPUT106), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n948), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n951), .B(KEYINPUT43), .Z(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(new_n948), .B2(new_n953), .ZN(new_n957));
  OAI21_X1  g0757(.A(KEYINPUT107), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT107), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n948), .A2(new_n953), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n959), .B(new_n954), .C1(new_n960), .C2(new_n956), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n942), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n666), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n958), .B(new_n961), .C1(new_n666), .C2(new_n963), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n672), .B(KEYINPUT41), .Z(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n668), .A2(new_n523), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n665), .B2(new_n668), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(new_n660), .Z(new_n971));
  NOR2_X1   g0771(.A1(new_n710), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n942), .A2(new_n669), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT45), .Z(new_n974));
  NOR2_X1   g0774(.A1(new_n942), .A2(new_n669), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT44), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n974), .A2(new_n666), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n666), .B1(new_n974), .B2(new_n976), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  AND3_X1   g0779(.A1(new_n972), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n968), .B1(new_n980), .B2(new_n710), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n715), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n965), .A2(new_n966), .A3(new_n982), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n767), .B1(new_n217), .B2(new_n314), .C1(new_n770), .C2(new_n232), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n984), .A2(new_n717), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n728), .A2(new_n487), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n742), .A2(new_n749), .B1(KEYINPUT46), .B2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(KEYINPUT108), .B(G317), .Z(new_n988));
  AOI22_X1  g0788(.A1(new_n733), .A2(new_n533), .B1(new_n723), .B2(new_n988), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n734), .A2(G294), .B1(new_n807), .B2(new_n793), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n986), .A2(KEYINPUT46), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n873), .B1(new_n528), .B2(new_n744), .C1(new_n560), .C2(new_n727), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n987), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G50), .A2(new_n793), .B1(new_n723), .B2(G137), .ZN(new_n995));
  INV_X1    g0795(.A(G159), .ZN(new_n996));
  INV_X1    g0796(.A(new_n734), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n995), .B1(new_n996), .B2(new_n997), .C1(new_n742), .C2(new_n795), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n281), .B1(new_n201), .B2(new_n728), .C1(new_n284), .C2(new_n744), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n727), .A2(new_n202), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G150), .B2(new_n733), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT109), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n994), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT47), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n985), .B1(new_n1005), .B2(new_n762), .C1(new_n780), .C2(new_n951), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n983), .A2(new_n1006), .ZN(G387));
  OAI21_X1  g0807(.A(new_n769), .B1(new_n229), .B2(new_n296), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n217), .A2(new_n281), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1008), .B1(new_n674), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n245), .A2(G50), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT50), .ZN(new_n1012));
  AOI21_X1  g0812(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(new_n674), .A3(new_n1013), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n1010), .A2(new_n1014), .B1(new_n327), .B2(new_n671), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n717), .B1(new_n1015), .B2(new_n768), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n751), .A2(new_n257), .B1(new_n736), .B2(new_n202), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n997), .A2(new_n245), .B1(new_n722), .B2(new_n247), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n753), .A2(G159), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n873), .B1(G97), .B2(new_n801), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n814), .A2(new_n553), .B1(new_n758), .B2(G77), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n397), .B1(G326), .B2(new_n723), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n988), .A2(new_n733), .B1(new_n734), .B2(G311), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n793), .A2(new_n533), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(new_n742), .C2(new_n750), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT48), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n814), .A2(new_n807), .B1(new_n758), .B2(G294), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT49), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1024), .B1(new_n487), .B2(new_n744), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1023), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1016), .B1(new_n1036), .B2(new_n761), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n665), .B2(new_n780), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n710), .A2(new_n971), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n672), .B1(new_n710), .B2(new_n971), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1038), .B1(new_n715), .B2(new_n971), .C1(new_n1039), .C2(new_n1040), .ZN(G393));
  AND2_X1   g0841(.A1(new_n979), .A2(new_n977), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1042), .A2(new_n972), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n972), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1043), .A2(new_n672), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1042), .A2(new_n716), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n237), .A2(new_n770), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n768), .B1(new_n671), .B2(G97), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n818), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n742), .A2(new_n247), .B1(new_n996), .B2(new_n751), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT111), .Z(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT110), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1053), .A2(KEYINPUT51), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n727), .A2(new_n284), .B1(new_n728), .B2(new_n202), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1055), .A2(new_n873), .A3(new_n813), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n382), .A2(new_n793), .B1(new_n723), .B2(G143), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n257), .C2(new_n997), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n1053), .B2(KEYINPUT51), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n753), .A2(G317), .B1(G311), .B2(new_n733), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT52), .Z(new_n1061));
  AOI22_X1  g0861(.A1(new_n734), .A2(new_n533), .B1(G322), .B2(new_n723), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n755), .B2(new_n736), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n727), .A2(new_n487), .B1(new_n806), .B2(new_n728), .ZN(new_n1064));
  NOR4_X1   g0864(.A1(new_n1063), .A2(new_n281), .A3(new_n745), .A4(new_n1064), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1054), .A2(new_n1059), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1050), .B1(new_n942), .B2(new_n780), .C1(new_n1066), .C2(new_n762), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1045), .A2(new_n1046), .A3(new_n1067), .ZN(G390));
  AND3_X1   g0868(.A1(new_n889), .A2(new_n918), .A3(KEYINPUT39), .ZN(new_n1069));
  AOI21_X1  g0869(.A(KEYINPUT39), .B1(new_n889), .B2(new_n894), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n1069), .A2(new_n1070), .B1(new_n925), .B2(new_n917), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n917), .B1(new_n889), .B2(new_n894), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT113), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT112), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n664), .A2(new_n548), .A3(new_n545), .A4(new_n543), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n635), .B1(new_n515), .B2(new_n522), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n939), .A2(new_n1075), .A3(new_n1076), .A4(new_n680), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n657), .B(new_n786), .C1(new_n1077), .C2(new_n637), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1074), .B1(new_n1078), .B2(new_n784), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n786), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n661), .B(new_n1080), .C1(new_n683), .C2(new_n686), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(KEYINPUT112), .A3(new_n923), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1079), .A2(new_n922), .A3(new_n1082), .ZN(new_n1083));
  AND3_X1   g0883(.A1(new_n1072), .A2(new_n1073), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1073), .B1(new_n1072), .B2(new_n1083), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1071), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n896), .A2(new_n707), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n922), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1071), .B(new_n1088), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1087), .A2(new_n922), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1094), .A2(new_n1095), .A3(new_n1088), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n924), .B1(new_n1089), .B2(new_n1093), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n466), .A2(new_n708), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n914), .A2(new_n1099), .A3(new_n650), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT114), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1100), .B1(new_n1097), .B2(new_n1096), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(KEYINPUT114), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1092), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1090), .A2(new_n1091), .A3(new_n1105), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1107), .A2(new_n672), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1090), .A2(new_n716), .A3(new_n1091), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n764), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n819), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n717), .B1(new_n382), .B2(new_n1112), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT115), .Z(new_n1114));
  INV_X1    g0914(.A(G125), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n997), .A2(new_n796), .B1(new_n722), .B2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT54), .B(G143), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n751), .A2(new_n799), .B1(new_n736), .B2(new_n1117), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1116), .B(new_n1118), .C1(G128), .C2(new_n753), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n728), .A2(new_n247), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT53), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n281), .B1(new_n257), .B2(new_n744), .C1(new_n996), .C2(new_n727), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1119), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT116), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n281), .B1(G87), .B2(new_n758), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n751), .A2(new_n487), .B1(new_n736), .B2(new_n528), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n997), .A2(new_n560), .B1(new_n722), .B2(new_n755), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n753), .A2(G283), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n814), .A2(G77), .B1(new_n801), .B2(G68), .ZN(new_n1133));
  AND4_X1   g0933(.A1(new_n1128), .A2(new_n1131), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  NOR3_X1   g0934(.A1(new_n1126), .A2(new_n1127), .A3(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1111), .B(new_n1114), .C1(new_n762), .C2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1109), .A2(new_n1110), .A3(new_n1136), .ZN(G378));
  INV_X1    g0937(.A(KEYINPUT119), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n929), .B(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n902), .A2(new_n908), .A3(G330), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(KEYINPUT118), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n649), .A2(new_n312), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n264), .A2(new_n861), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1142), .B(new_n1143), .ZN(new_n1144));
  XOR2_X1   g0944(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1145));
  XOR2_X1   g0945(.A(new_n1144), .B(new_n1145), .Z(new_n1146));
  INV_X1    g0946(.A(KEYINPUT118), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n902), .A2(new_n908), .A3(new_n1147), .A4(G330), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1141), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1144), .B(new_n1145), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n909), .A2(new_n1150), .A3(new_n1147), .A4(G330), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1139), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1152), .B1(new_n1153), .B2(new_n929), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1108), .A2(new_n1101), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT57), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT57), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n1108), .B2(new_n1101), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1149), .A2(new_n929), .A3(new_n1151), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n929), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n672), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n1156), .A2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n717), .B1(G50), .B2(new_n1112), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n257), .B1(G33), .B2(G41), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n873), .B2(new_n295), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n751), .A2(new_n327), .B1(new_n314), .B2(new_n736), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n997), .A2(new_n528), .B1(new_n722), .B2(new_n756), .ZN(new_n1168));
  NOR4_X1   g0968(.A1(new_n1167), .A2(new_n1168), .A3(G41), .A4(new_n397), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n744), .A2(new_n201), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1170), .B(new_n1001), .C1(G77), .C2(new_n758), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(new_n487), .C2(new_n742), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT58), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1166), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(G128), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n1175), .A2(new_n751), .B1(new_n997), .B2(new_n799), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G137), .B2(new_n793), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1117), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n814), .A2(G150), .B1(new_n758), .B2(new_n1178), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1177), .B(new_n1179), .C1(new_n1115), .C2(new_n742), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(KEYINPUT59), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n801), .A2(G159), .ZN(new_n1182));
  AOI211_X1 g0982(.A(G33), .B(G41), .C1(new_n723), .C2(G124), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1180), .A2(KEYINPUT59), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1174), .B1(new_n1173), .B2(new_n1172), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1164), .B1(new_n1186), .B2(new_n761), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n1146), .B2(new_n765), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT117), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n1154), .B2(new_n716), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1163), .A2(new_n1190), .ZN(G375));
  NAND3_X1  g0991(.A1(new_n1100), .A2(new_n1097), .A3(new_n1096), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1104), .A2(new_n1106), .A3(new_n968), .A4(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT120), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n897), .A2(new_n899), .A3(new_n764), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n796), .A2(new_n751), .B1(new_n997), .B2(new_n1117), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n201), .A2(new_n744), .B1(new_n728), .B2(new_n996), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n397), .B1(new_n1175), .B2(new_n722), .C1(new_n247), .C2(new_n736), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(G50), .C2(new_n814), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT122), .Z(new_n1200));
  AOI211_X1 g1000(.A(new_n1196), .B(new_n1200), .C1(G132), .C2(new_n753), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n734), .A2(G116), .B1(new_n331), .B2(new_n793), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n733), .A2(G283), .B1(G303), .B2(new_n723), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(new_n742), .C2(new_n755), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n326), .B1(new_n284), .B2(new_n744), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n727), .A2(new_n314), .B1(new_n728), .B2(new_n528), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n761), .B1(new_n1201), .B2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n717), .B1(G68), .B2(new_n1112), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT121), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT123), .Z(new_n1212));
  AOI22_X1  g1012(.A1(new_n1098), .A2(new_n716), .B1(new_n1195), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1194), .A2(new_n1213), .ZN(G381));
  INV_X1    g1014(.A(G375), .ZN(new_n1215));
  INV_X1    g1015(.A(G378), .ZN(new_n1216));
  INV_X1    g1016(.A(G390), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1217), .A2(new_n1006), .A3(new_n983), .ZN(new_n1218));
  OR2_X1    g1018(.A1(G393), .A2(G396), .ZN(new_n1219));
  NOR4_X1   g1019(.A1(new_n1218), .A2(G381), .A3(G384), .A4(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1215), .A2(new_n1216), .A3(new_n1220), .ZN(G407));
  NAND2_X1  g1021(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1222));
  OAI211_X1 g1022(.A(G407), .B(G213), .C1(new_n1222), .C2(G343), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT124), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1223), .B(new_n1224), .ZN(G409));
  NAND2_X1  g1025(.A1(G387), .A2(G390), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT126), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1226), .A2(new_n1227), .A3(new_n1218), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT127), .ZN(new_n1229));
  XOR2_X1   g1029(.A(G393), .B(G396), .Z(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1228), .A2(new_n1229), .A3(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1226), .A2(KEYINPUT127), .A3(new_n1218), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1231), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G378), .B(new_n1190), .C1(new_n1156), .C2(new_n1162), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1139), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n968), .B(new_n1155), .C1(new_n1238), .C2(new_n1160), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n716), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n1188), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1216), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1237), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n656), .A2(G213), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT60), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1192), .B1(new_n1105), .B2(new_n1245), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1100), .A2(new_n1096), .A3(new_n1097), .A4(KEYINPUT60), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1246), .A2(new_n672), .A3(new_n1247), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1248), .A2(G384), .A3(new_n1213), .ZN(new_n1249));
  AOI21_X1  g1049(.A(G384), .B1(new_n1248), .B2(new_n1213), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1243), .A2(new_n1244), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT125), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT125), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1243), .A2(new_n1254), .A3(new_n1244), .A4(new_n1251), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT62), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n656), .A2(G213), .A3(G2897), .ZN(new_n1258));
  XOR2_X1   g1058(.A(new_n1251), .B(new_n1258), .Z(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT61), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1252), .A2(KEYINPUT62), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1236), .B1(new_n1256), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT63), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1253), .A2(new_n1264), .A3(new_n1255), .ZN(new_n1265));
  OR2_X1    g1065(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1266));
  OR2_X1    g1066(.A1(new_n1252), .A2(new_n1264), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1265), .A2(new_n1266), .A3(new_n1260), .A4(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1263), .A2(new_n1268), .ZN(G405));
  NAND2_X1  g1069(.A1(G375), .A2(new_n1216), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1237), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1251), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1270), .B(new_n1237), .C1(new_n1250), .C2(new_n1249), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n1272), .A2(new_n1236), .A3(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1236), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(G402));
endmodule


