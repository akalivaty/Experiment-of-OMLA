

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744;

  XNOR2_X2 U372 ( .A(n542), .B(n410), .ZN(n409) );
  XNOR2_X2 U373 ( .A(n508), .B(n507), .ZN(n636) );
  XNOR2_X2 U374 ( .A(n441), .B(n440), .ZN(n520) );
  XNOR2_X2 U375 ( .A(KEYINPUT41), .B(n551), .ZN(n666) );
  XNOR2_X2 U376 ( .A(n480), .B(G469), .ZN(n534) );
  XNOR2_X1 U377 ( .A(n400), .B(KEYINPUT35), .ZN(n742) );
  XNOR2_X1 U378 ( .A(n613), .B(n612), .ZN(n614) );
  NOR2_X1 U379 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U380 ( .A1(n404), .A2(n350), .ZN(n548) );
  NOR2_X1 U381 ( .A1(n581), .A2(n742), .ZN(n363) );
  NAND2_X1 U382 ( .A1(n395), .A2(n394), .ZN(n400) );
  NAND2_X1 U383 ( .A1(n385), .A2(n509), .ZN(n569) );
  XNOR2_X1 U384 ( .A(n384), .B(KEYINPUT32), .ZN(n570) );
  NAND2_X1 U385 ( .A1(n418), .A2(n642), .ZN(n593) );
  XNOR2_X1 U386 ( .A(n554), .B(n553), .ZN(n740) );
  XNOR2_X1 U387 ( .A(n419), .B(n451), .ZN(n578) );
  XNOR2_X1 U388 ( .A(n525), .B(KEYINPUT65), .ZN(n573) );
  AND2_X1 U389 ( .A1(n532), .A2(n640), .ZN(n533) );
  XNOR2_X1 U390 ( .A(n539), .B(KEYINPUT104), .ZN(n389) );
  XNOR2_X1 U391 ( .A(n515), .B(KEYINPUT103), .ZN(n557) );
  NAND2_X1 U392 ( .A1(n371), .A2(n489), .ZN(n508) );
  XNOR2_X1 U393 ( .A(G478), .B(n468), .ZN(n537) );
  XNOR2_X1 U394 ( .A(n388), .B(n387), .ZN(n497) );
  INV_X2 U395 ( .A(G953), .ZN(n732) );
  AND2_X1 U396 ( .A1(n555), .A2(n518), .ZN(n655) );
  XNOR2_X1 U397 ( .A(n548), .B(n547), .ZN(n562) );
  BUF_X1 U398 ( .A(n617), .Z(n349) );
  XNOR2_X1 U399 ( .A(n361), .B(KEYINPUT45), .ZN(n617) );
  XNOR2_X2 U400 ( .A(n370), .B(n369), .ZN(n418) );
  NOR2_X2 U401 ( .A1(n534), .A2(n573), .ZN(n587) );
  NOR2_X1 U402 ( .A1(n535), .A2(n534), .ZN(n552) );
  NAND2_X1 U403 ( .A1(n683), .A2(n389), .ZN(n386) );
  NAND2_X1 U404 ( .A1(n536), .A2(n450), .ZN(n419) );
  NOR2_X1 U405 ( .A1(n537), .A2(n538), .ZN(n515) );
  INV_X1 U406 ( .A(KEYINPUT78), .ZN(n410) );
  INV_X1 U407 ( .A(KEYINPUT19), .ZN(n366) );
  NAND2_X1 U408 ( .A1(n569), .A2(n570), .ZN(n571) );
  XNOR2_X1 U409 ( .A(G119), .B(G128), .ZN(n491) );
  INV_X1 U410 ( .A(KEYINPUT8), .ZN(n387) );
  NAND2_X1 U411 ( .A1(n732), .A2(G234), .ZN(n388) );
  XNOR2_X1 U412 ( .A(G146), .B(G125), .ZN(n452) );
  XNOR2_X1 U413 ( .A(n506), .B(KEYINPUT25), .ZN(n507) );
  XNOR2_X1 U414 ( .A(n462), .B(n392), .ZN(n391) );
  XNOR2_X1 U415 ( .A(n463), .B(KEYINPUT7), .ZN(n392) );
  XNOR2_X1 U416 ( .A(n403), .B(G116), .ZN(n465) );
  XNOR2_X1 U417 ( .A(KEYINPUT98), .B(KEYINPUT12), .ZN(n378) );
  XNOR2_X1 U418 ( .A(G131), .B(G143), .ZN(n456) );
  XNOR2_X1 U419 ( .A(G113), .B(G104), .ZN(n453) );
  XOR2_X1 U420 ( .A(G140), .B(G122), .Z(n454) );
  XNOR2_X1 U421 ( .A(n380), .B(KEYINPUT11), .ZN(n379) );
  NAND2_X1 U422 ( .A1(n483), .A2(G214), .ZN(n380) );
  INV_X1 U423 ( .A(KEYINPUT22), .ZN(n369) );
  NAND2_X1 U424 ( .A1(n578), .A2(n352), .ZN(n370) );
  INV_X1 U425 ( .A(n520), .ZN(n367) );
  AND2_X1 U426 ( .A1(n412), .A2(n587), .ZN(n556) );
  AND2_X1 U427 ( .A1(n529), .A2(n528), .ZN(n412) );
  OR2_X1 U428 ( .A1(G902), .A2(n711), .ZN(n468) );
  XNOR2_X1 U429 ( .A(n383), .B(n381), .ZN(n538) );
  XNOR2_X1 U430 ( .A(n459), .B(n382), .ZN(n381) );
  OR2_X1 U431 ( .A1(n705), .A2(G902), .ZN(n383) );
  INV_X1 U432 ( .A(G475), .ZN(n382) );
  NAND2_X1 U433 ( .A1(n406), .A2(n543), .ZN(n405) );
  XNOR2_X1 U434 ( .A(G146), .B(G137), .ZN(n481) );
  XOR2_X1 U435 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n482) );
  XNOR2_X1 U436 ( .A(n560), .B(n374), .ZN(n561) );
  XNOR2_X1 U437 ( .A(n559), .B(KEYINPUT64), .ZN(n374) );
  XNOR2_X1 U438 ( .A(n416), .B(n415), .ZN(n487) );
  XNOR2_X1 U439 ( .A(G116), .B(G113), .ZN(n415) );
  XNOR2_X1 U440 ( .A(n421), .B(G119), .ZN(n416) );
  XNOR2_X1 U441 ( .A(G101), .B(KEYINPUT3), .ZN(n421) );
  XNOR2_X1 U442 ( .A(G134), .B(G107), .ZN(n460) );
  NOR2_X1 U443 ( .A1(G953), .A2(G237), .ZN(n483) );
  XNOR2_X1 U444 ( .A(n474), .B(n473), .ZN(n486) );
  XNOR2_X1 U445 ( .A(G131), .B(G134), .ZN(n473) );
  XNOR2_X1 U446 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n428) );
  NAND2_X1 U447 ( .A1(G234), .A2(G237), .ZN(n444) );
  INV_X1 U448 ( .A(G237), .ZN(n436) );
  NAND2_X1 U449 ( .A1(n353), .A2(n364), .ZN(n536) );
  NAND2_X1 U450 ( .A1(n367), .A2(n356), .ZN(n364) );
  NAND2_X1 U451 ( .A1(n651), .A2(KEYINPUT19), .ZN(n368) );
  XNOR2_X1 U452 ( .A(G107), .B(G104), .ZN(n425) );
  XNOR2_X1 U453 ( .A(n487), .B(n422), .ZN(n724) );
  XNOR2_X1 U454 ( .A(KEYINPUT16), .B(G122), .ZN(n422) );
  INV_X1 U455 ( .A(KEYINPUT80), .ZN(n498) );
  XNOR2_X1 U456 ( .A(KEYINPUT94), .B(KEYINPUT24), .ZN(n493) );
  XOR2_X1 U457 ( .A(G137), .B(G140), .Z(n502) );
  XNOR2_X1 U458 ( .A(n475), .B(KEYINPUT73), .ZN(n477) );
  XNOR2_X1 U459 ( .A(n486), .B(n402), .ZN(n730) );
  INV_X1 U460 ( .A(n502), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n373), .B(n372), .ZN(n564) );
  INV_X1 U462 ( .A(KEYINPUT39), .ZN(n372) );
  AND2_X1 U463 ( .A1(n397), .A2(n580), .ZN(n396) );
  NAND2_X1 U464 ( .A1(n398), .A2(KEYINPUT34), .ZN(n397) );
  XNOR2_X1 U465 ( .A(n466), .B(n390), .ZN(n711) );
  XNOR2_X1 U466 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U467 ( .A(n467), .B(n391), .ZN(n390) );
  XNOR2_X1 U468 ( .A(n379), .B(n377), .ZN(n457) );
  XNOR2_X1 U469 ( .A(n456), .B(n378), .ZN(n377) );
  XNOR2_X1 U470 ( .A(n730), .B(n401), .ZN(n702) );
  XNOR2_X1 U471 ( .A(n478), .B(n479), .ZN(n401) );
  XNOR2_X1 U472 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U473 ( .A(G101), .B(G146), .ZN(n476) );
  AND2_X1 U474 ( .A1(n606), .A2(G953), .ZN(n717) );
  AND2_X1 U475 ( .A1(n375), .A2(n522), .ZN(n697) );
  XNOR2_X1 U476 ( .A(n376), .B(n545), .ZN(n375) );
  XNOR2_X1 U477 ( .A(n557), .B(KEYINPUT107), .ZN(n688) );
  AND2_X1 U478 ( .A1(n580), .A2(n367), .ZN(n411) );
  XNOR2_X1 U479 ( .A(n593), .B(n417), .ZN(n385) );
  INV_X1 U480 ( .A(KEYINPUT106), .ZN(n417) );
  AND2_X1 U481 ( .A1(n409), .A2(n360), .ZN(n350) );
  BUF_X1 U482 ( .A(n578), .Z(n583) );
  INV_X1 U483 ( .A(n583), .ZN(n398) );
  OR2_X1 U484 ( .A1(n386), .A2(KEYINPUT47), .ZN(n351) );
  AND2_X1 U485 ( .A1(n653), .A2(n472), .ZN(n352) );
  AND2_X1 U486 ( .A1(n365), .A2(n368), .ZN(n353) );
  AND2_X1 U487 ( .A1(n367), .A2(n518), .ZN(n354) );
  AND2_X1 U488 ( .A1(n546), .A2(n405), .ZN(n355) );
  AND2_X1 U489 ( .A1(n518), .A2(n366), .ZN(n356) );
  NOR2_X1 U490 ( .A1(n527), .A2(n635), .ZN(n357) );
  AND2_X1 U491 ( .A1(n516), .A2(n354), .ZN(n358) );
  BUF_X1 U492 ( .A(n520), .Z(n550) );
  AND2_X1 U493 ( .A1(n524), .A2(n523), .ZN(n359) );
  AND2_X1 U494 ( .A1(n351), .A2(KEYINPUT69), .ZN(n360) );
  AND2_X1 U495 ( .A1(n556), .A2(n411), .ZN(n531) );
  NAND2_X1 U496 ( .A1(n362), .A2(n596), .ZN(n361) );
  XNOR2_X1 U497 ( .A(n363), .B(KEYINPUT44), .ZN(n362) );
  NAND2_X1 U498 ( .A1(n520), .A2(KEYINPUT19), .ZN(n365) );
  NAND2_X1 U499 ( .A1(n418), .A2(n359), .ZN(n384) );
  NAND2_X1 U500 ( .A1(n617), .A2(n628), .ZN(n625) );
  INV_X1 U501 ( .A(n714), .ZN(n371) );
  XNOR2_X1 U502 ( .A(n504), .B(n503), .ZN(n714) );
  NOR2_X1 U503 ( .A1(n582), .A2(n591), .ZN(n577) );
  XNOR2_X1 U504 ( .A(n575), .B(KEYINPUT71), .ZN(n582) );
  NAND2_X1 U505 ( .A1(n556), .A2(n555), .ZN(n373) );
  NAND2_X1 U506 ( .A1(n688), .A2(n516), .ZN(n544) );
  NAND2_X1 U507 ( .A1(n688), .A2(n358), .ZN(n376) );
  NAND2_X1 U508 ( .A1(n386), .A2(KEYINPUT47), .ZN(n540) );
  NAND2_X1 U509 ( .A1(n497), .A2(G221), .ZN(n499) );
  INV_X1 U510 ( .A(n636), .ZN(n590) );
  AND2_X1 U511 ( .A1(n636), .A2(n357), .ZN(n532) );
  NAND2_X1 U512 ( .A1(n389), .A2(n655), .ZN(n656) );
  NAND2_X1 U513 ( .A1(n589), .A2(n389), .ZN(n595) );
  XNOR2_X1 U514 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U515 ( .A(n501), .B(n500), .ZN(n504) );
  AND2_X1 U516 ( .A1(n536), .A2(n552), .ZN(n683) );
  AND2_X2 U517 ( .A1(n710), .A2(G472), .ZN(n613) );
  NOR2_X2 U518 ( .A1(n614), .A2(n717), .ZN(n616) );
  AND2_X1 U519 ( .A1(n393), .A2(n396), .ZN(n395) );
  NAND2_X1 U520 ( .A1(n665), .A2(n399), .ZN(n393) );
  OR2_X1 U521 ( .A1(n665), .A2(n579), .ZN(n394) );
  AND2_X1 U522 ( .A1(n583), .A2(n579), .ZN(n399) );
  XNOR2_X2 U523 ( .A(n403), .B(n424), .ZN(n474) );
  XNOR2_X2 U524 ( .A(n423), .B(G143), .ZN(n403) );
  NAND2_X1 U525 ( .A1(n407), .A2(n355), .ZN(n404) );
  INV_X1 U526 ( .A(n351), .ZN(n406) );
  NAND2_X1 U527 ( .A1(n408), .A2(n543), .ZN(n407) );
  INV_X1 U528 ( .A(n409), .ZN(n408) );
  XNOR2_X2 U529 ( .A(n413), .B(n490), .ZN(n586) );
  NAND2_X1 U530 ( .A1(n611), .A2(n489), .ZN(n413) );
  XNOR2_X1 U531 ( .A(n486), .B(n414), .ZN(n611) );
  XNOR2_X1 U532 ( .A(n488), .B(n485), .ZN(n414) );
  AND2_X1 U533 ( .A1(n483), .A2(G210), .ZN(n420) );
  INV_X1 U534 ( .A(KEYINPUT69), .ZN(n543) );
  INV_X1 U535 ( .A(KEYINPUT66), .ZN(n547) );
  XNOR2_X1 U536 ( .A(n484), .B(n420), .ZN(n485) );
  INV_X1 U537 ( .A(KEYINPUT33), .ZN(n576) );
  INV_X1 U538 ( .A(n527), .ZN(n528) );
  INV_X1 U539 ( .A(KEYINPUT102), .ZN(n464) );
  INV_X1 U540 ( .A(n688), .ZN(n691) );
  XNOR2_X2 U541 ( .A(G128), .B(KEYINPUT75), .ZN(n423) );
  INV_X1 U542 ( .A(KEYINPUT4), .ZN(n424) );
  XNOR2_X1 U543 ( .A(n724), .B(n474), .ZN(n433) );
  XNOR2_X1 U544 ( .A(n425), .B(G110), .ZN(n722) );
  INV_X1 U545 ( .A(KEYINPUT68), .ZN(n426) );
  XNOR2_X1 U546 ( .A(n722), .B(n426), .ZN(n479) );
  NAND2_X1 U547 ( .A1(n732), .A2(G224), .ZN(n427) );
  XNOR2_X1 U548 ( .A(n427), .B(KEYINPUT90), .ZN(n429) );
  XNOR2_X1 U549 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U550 ( .A(n452), .B(n430), .ZN(n431) );
  XNOR2_X1 U551 ( .A(n479), .B(n431), .ZN(n432) );
  XNOR2_X1 U552 ( .A(n433), .B(n432), .ZN(n600) );
  XNOR2_X1 U553 ( .A(G902), .B(KEYINPUT89), .ZN(n435) );
  INV_X1 U554 ( .A(KEYINPUT15), .ZN(n434) );
  XNOR2_X1 U555 ( .A(n435), .B(n434), .ZN(n597) );
  NAND2_X1 U556 ( .A1(n600), .A2(n597), .ZN(n441) );
  INV_X1 U557 ( .A(G902), .ZN(n489) );
  NAND2_X1 U558 ( .A1(n489), .A2(n436), .ZN(n442) );
  NAND2_X1 U559 ( .A1(n442), .A2(G210), .ZN(n439) );
  INV_X1 U560 ( .A(KEYINPUT76), .ZN(n437) );
  XNOR2_X1 U561 ( .A(n437), .B(KEYINPUT91), .ZN(n438) );
  XNOR2_X1 U562 ( .A(n439), .B(n438), .ZN(n440) );
  NAND2_X1 U563 ( .A1(n442), .A2(G214), .ZN(n443) );
  XNOR2_X1 U564 ( .A(n443), .B(KEYINPUT92), .ZN(n518) );
  INV_X1 U565 ( .A(n518), .ZN(n651) );
  XNOR2_X1 U566 ( .A(n444), .B(KEYINPUT14), .ZN(n446) );
  NAND2_X1 U567 ( .A1(G952), .A2(n446), .ZN(n663) );
  NOR2_X1 U568 ( .A1(n663), .A2(G953), .ZN(n513) );
  INV_X1 U569 ( .A(n513), .ZN(n449) );
  AND2_X1 U570 ( .A1(G953), .A2(G902), .ZN(n445) );
  NAND2_X1 U571 ( .A1(n446), .A2(n445), .ZN(n510) );
  NOR2_X1 U572 ( .A1(G898), .A2(n510), .ZN(n447) );
  XNOR2_X1 U573 ( .A(n447), .B(KEYINPUT93), .ZN(n448) );
  NAND2_X1 U574 ( .A1(n449), .A2(n448), .ZN(n450) );
  INV_X1 U575 ( .A(KEYINPUT0), .ZN(n451) );
  XNOR2_X1 U576 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n459) );
  XNOR2_X1 U577 ( .A(KEYINPUT10), .B(n452), .ZN(n729) );
  XNOR2_X1 U578 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U579 ( .A(n729), .B(n455), .ZN(n458) );
  XNOR2_X1 U580 ( .A(n458), .B(n457), .ZN(n705) );
  XOR2_X1 U581 ( .A(KEYINPUT101), .B(G122), .Z(n461) );
  XNOR2_X1 U582 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U583 ( .A(KEYINPUT100), .B(KEYINPUT9), .ZN(n463) );
  NAND2_X1 U584 ( .A1(n497), .A2(G217), .ZN(n467) );
  INV_X1 U585 ( .A(n537), .ZN(n530) );
  AND2_X1 U586 ( .A1(n538), .A2(n530), .ZN(n653) );
  XOR2_X1 U587 ( .A(KEYINPUT20), .B(KEYINPUT95), .Z(n470) );
  NAND2_X1 U588 ( .A1(G234), .A2(n597), .ZN(n469) );
  XNOR2_X1 U589 ( .A(n470), .B(n469), .ZN(n505) );
  NAND2_X1 U590 ( .A1(n505), .A2(G221), .ZN(n471) );
  XNOR2_X1 U591 ( .A(n471), .B(KEYINPUT21), .ZN(n635) );
  INV_X1 U592 ( .A(n635), .ZN(n472) );
  AND2_X1 U593 ( .A1(G227), .A2(n732), .ZN(n475) );
  NOR2_X1 U594 ( .A1(n702), .A2(G902), .ZN(n480) );
  XNOR2_X1 U595 ( .A(n534), .B(KEYINPUT1), .ZN(n574) );
  INV_X1 U596 ( .A(n574), .ZN(n522) );
  XNOR2_X1 U597 ( .A(n482), .B(n481), .ZN(n484) );
  INV_X1 U598 ( .A(n487), .ZN(n488) );
  INV_X1 U599 ( .A(G472), .ZN(n490) );
  INV_X1 U600 ( .A(n586), .ZN(n640) );
  XOR2_X1 U601 ( .A(KEYINPUT23), .B(G110), .Z(n492) );
  XNOR2_X1 U602 ( .A(n492), .B(n491), .ZN(n496) );
  XOR2_X1 U603 ( .A(KEYINPUT72), .B(KEYINPUT67), .Z(n494) );
  XNOR2_X1 U604 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U605 ( .A(n496), .B(n495), .Z(n501) );
  XNOR2_X1 U606 ( .A(n502), .B(n729), .ZN(n503) );
  NAND2_X1 U607 ( .A1(n505), .A2(G217), .ZN(n506) );
  NOR2_X1 U608 ( .A1(n640), .A2(n590), .ZN(n509) );
  XNOR2_X1 U609 ( .A(n569), .B(G110), .ZN(G12) );
  XNOR2_X1 U610 ( .A(n586), .B(KEYINPUT6), .ZN(n572) );
  XNOR2_X1 U611 ( .A(KEYINPUT108), .B(n510), .ZN(n511) );
  NOR2_X1 U612 ( .A1(G900), .A2(n511), .ZN(n512) );
  NOR2_X1 U613 ( .A1(n513), .A2(n512), .ZN(n527) );
  NAND2_X1 U614 ( .A1(n572), .A2(n532), .ZN(n514) );
  XNOR2_X1 U615 ( .A(KEYINPUT109), .B(n514), .ZN(n516) );
  NOR2_X1 U616 ( .A1(n522), .A2(n544), .ZN(n517) );
  NAND2_X1 U617 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U618 ( .A(KEYINPUT43), .B(n519), .ZN(n521) );
  AND2_X1 U619 ( .A1(n521), .A2(n550), .ZN(n566) );
  XOR2_X1 U620 ( .A(n566), .B(G140), .Z(G42) );
  INV_X1 U621 ( .A(n522), .ZN(n642) );
  NOR2_X1 U622 ( .A1(n642), .A2(n590), .ZN(n524) );
  XOR2_X1 U623 ( .A(KEYINPUT74), .B(n572), .Z(n523) );
  XNOR2_X1 U624 ( .A(n570), .B(G119), .ZN(G21) );
  NOR2_X1 U625 ( .A1(n636), .A2(n635), .ZN(n525) );
  NOR2_X1 U626 ( .A1(n651), .A2(n586), .ZN(n526) );
  XNOR2_X1 U627 ( .A(KEYINPUT30), .B(n526), .ZN(n529) );
  NOR2_X1 U628 ( .A1(n538), .A2(n530), .ZN(n580) );
  XOR2_X1 U629 ( .A(G143), .B(n531), .Z(G45) );
  XNOR2_X1 U630 ( .A(n531), .B(KEYINPUT79), .ZN(n541) );
  XOR2_X1 U631 ( .A(KEYINPUT28), .B(n533), .Z(n535) );
  NAND2_X1 U632 ( .A1(n538), .A2(n537), .ZN(n694) );
  NAND2_X1 U633 ( .A1(n694), .A2(n557), .ZN(n539) );
  NAND2_X1 U634 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U635 ( .A(KEYINPUT87), .B(KEYINPUT36), .ZN(n545) );
  INV_X1 U636 ( .A(n697), .ZN(n546) );
  XOR2_X1 U637 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n554) );
  XNOR2_X1 U638 ( .A(KEYINPUT70), .B(KEYINPUT38), .ZN(n549) );
  XNOR2_X1 U639 ( .A(n550), .B(n549), .ZN(n555) );
  INV_X1 U640 ( .A(n555), .ZN(n652) );
  NAND2_X1 U641 ( .A1(n653), .A2(n655), .ZN(n551) );
  NAND2_X1 U642 ( .A1(n552), .A2(n666), .ZN(n553) );
  NOR2_X1 U643 ( .A1(n564), .A2(n557), .ZN(n558) );
  XNOR2_X1 U644 ( .A(KEYINPUT40), .B(n558), .ZN(n744) );
  NOR2_X1 U645 ( .A1(n740), .A2(n744), .ZN(n560) );
  XNOR2_X1 U646 ( .A(KEYINPUT46), .B(KEYINPUT85), .ZN(n559) );
  XNOR2_X1 U647 ( .A(n563), .B(KEYINPUT48), .ZN(n568) );
  OR2_X1 U648 ( .A1(n694), .A2(n564), .ZN(n565) );
  XNOR2_X1 U649 ( .A(n565), .B(KEYINPUT111), .ZN(n739) );
  NOR2_X1 U650 ( .A1(n739), .A2(n566), .ZN(n567) );
  AND2_X2 U651 ( .A1(n568), .A2(n567), .ZN(n628) );
  XNOR2_X1 U652 ( .A(n571), .B(KEYINPUT86), .ZN(n581) );
  INV_X1 U653 ( .A(n572), .ZN(n591) );
  NOR2_X1 U654 ( .A1(n573), .A2(n574), .ZN(n575) );
  XNOR2_X1 U655 ( .A(n577), .B(n576), .ZN(n665) );
  INV_X1 U656 ( .A(KEYINPUT34), .ZN(n579) );
  NOR2_X1 U657 ( .A1(n582), .A2(n586), .ZN(n647) );
  NAND2_X1 U658 ( .A1(n647), .A2(n583), .ZN(n584) );
  XNOR2_X1 U659 ( .A(n584), .B(KEYINPUT97), .ZN(n585) );
  XNOR2_X1 U660 ( .A(KEYINPUT31), .B(n585), .ZN(n693) );
  NAND2_X1 U661 ( .A1(n587), .A2(n586), .ZN(n588) );
  OR2_X1 U662 ( .A1(n588), .A2(n398), .ZN(n680) );
  NAND2_X1 U663 ( .A1(n693), .A2(n680), .ZN(n589) );
  NAND2_X1 U664 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U666 ( .A(n594), .B(KEYINPUT105), .ZN(n743) );
  AND2_X1 U667 ( .A1(n595), .A2(n743), .ZN(n596) );
  XNOR2_X1 U668 ( .A(n625), .B(KEYINPUT2), .ZN(n599) );
  INV_X1 U669 ( .A(n597), .ZN(n598) );
  AND2_X2 U670 ( .A1(n599), .A2(n598), .ZN(n710) );
  NAND2_X1 U671 ( .A1(n710), .A2(G210), .ZN(n605) );
  XOR2_X1 U672 ( .A(KEYINPUT54), .B(KEYINPUT124), .Z(n602) );
  XNOR2_X1 U673 ( .A(KEYINPUT77), .B(KEYINPUT55), .ZN(n601) );
  XNOR2_X1 U674 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U675 ( .A(n600), .B(n603), .ZN(n604) );
  XNOR2_X1 U676 ( .A(n605), .B(n604), .ZN(n607) );
  INV_X1 U677 ( .A(G952), .ZN(n606) );
  NOR2_X2 U678 ( .A1(n607), .A2(n717), .ZN(n610) );
  XNOR2_X1 U679 ( .A(KEYINPUT125), .B(KEYINPUT56), .ZN(n608) );
  XOR2_X1 U680 ( .A(n608), .B(KEYINPUT84), .Z(n609) );
  XNOR2_X1 U681 ( .A(n610), .B(n609), .ZN(G51) );
  XNOR2_X1 U682 ( .A(n611), .B(KEYINPUT62), .ZN(n612) );
  XOR2_X1 U683 ( .A(KEYINPUT88), .B(KEYINPUT63), .Z(n615) );
  XNOR2_X1 U684 ( .A(n616), .B(n615), .ZN(G57) );
  NOR2_X1 U685 ( .A1(n349), .A2(KEYINPUT81), .ZN(n622) );
  INV_X1 U686 ( .A(n628), .ZN(n618) );
  NAND2_X1 U687 ( .A1(n618), .A2(KEYINPUT82), .ZN(n620) );
  INV_X1 U688 ( .A(KEYINPUT2), .ZN(n619) );
  NAND2_X1 U689 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U690 ( .A1(n622), .A2(n621), .ZN(n627) );
  NAND2_X1 U691 ( .A1(KEYINPUT2), .A2(KEYINPUT82), .ZN(n623) );
  NOR2_X1 U692 ( .A1(n623), .A2(KEYINPUT81), .ZN(n624) );
  AND2_X1 U693 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U694 ( .A1(n627), .A2(n626), .ZN(n633) );
  NAND2_X1 U695 ( .A1(n349), .A2(KEYINPUT81), .ZN(n631) );
  INV_X1 U696 ( .A(KEYINPUT82), .ZN(n629) );
  NAND2_X1 U697 ( .A1(n628), .A2(n629), .ZN(n630) );
  NAND2_X1 U698 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U699 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U700 ( .A(n634), .B(KEYINPUT83), .ZN(n672) );
  XOR2_X1 U701 ( .A(KEYINPUT52), .B(KEYINPUT121), .Z(n662) );
  NAND2_X1 U702 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U703 ( .A(n637), .B(KEYINPUT49), .ZN(n638) );
  XNOR2_X1 U704 ( .A(n638), .B(KEYINPUT118), .ZN(n639) );
  NOR2_X1 U705 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U706 ( .A(KEYINPUT119), .B(n641), .ZN(n645) );
  NAND2_X1 U707 ( .A1(n642), .A2(n573), .ZN(n643) );
  XOR2_X1 U708 ( .A(KEYINPUT50), .B(n643), .Z(n644) );
  NOR2_X1 U709 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U710 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U711 ( .A(KEYINPUT51), .B(n648), .ZN(n649) );
  NAND2_X1 U712 ( .A1(n649), .A2(n666), .ZN(n650) );
  XNOR2_X1 U713 ( .A(n650), .B(KEYINPUT120), .ZN(n660) );
  NAND2_X1 U714 ( .A1(n652), .A2(n651), .ZN(n654) );
  NAND2_X1 U715 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U716 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U717 ( .A1(n665), .A2(n658), .ZN(n659) );
  NAND2_X1 U718 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U719 ( .A(n662), .B(n661), .Z(n664) );
  NOR2_X1 U720 ( .A1(n664), .A2(n663), .ZN(n670) );
  NAND2_X1 U721 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U722 ( .A(n667), .B(KEYINPUT122), .ZN(n668) );
  NAND2_X1 U723 ( .A1(n668), .A2(n732), .ZN(n669) );
  NOR2_X1 U724 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U725 ( .A1(n672), .A2(n671), .ZN(n674) );
  XNOR2_X1 U726 ( .A(KEYINPUT123), .B(KEYINPUT53), .ZN(n673) );
  XNOR2_X1 U727 ( .A(n674), .B(n673), .ZN(G75) );
  NOR2_X1 U728 ( .A1(n691), .A2(n680), .ZN(n676) );
  XNOR2_X1 U729 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n675) );
  XNOR2_X1 U730 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U731 ( .A(G104), .B(n677), .ZN(G6) );
  XOR2_X1 U732 ( .A(KEYINPUT26), .B(KEYINPUT114), .Z(n679) );
  XNOR2_X1 U733 ( .A(G107), .B(KEYINPUT27), .ZN(n678) );
  XNOR2_X1 U734 ( .A(n679), .B(n678), .ZN(n682) );
  NOR2_X1 U735 ( .A1(n694), .A2(n680), .ZN(n681) );
  XOR2_X1 U736 ( .A(n682), .B(n681), .Z(G9) );
  XOR2_X1 U737 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n686) );
  BUF_X1 U738 ( .A(n683), .Z(n689) );
  INV_X1 U739 ( .A(n694), .ZN(n684) );
  NAND2_X1 U740 ( .A1(n689), .A2(n684), .ZN(n685) );
  XNOR2_X1 U741 ( .A(n686), .B(n685), .ZN(n687) );
  XOR2_X1 U742 ( .A(G128), .B(n687), .Z(G30) );
  NAND2_X1 U743 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U744 ( .A(n690), .B(G146), .ZN(G48) );
  NOR2_X1 U745 ( .A1(n691), .A2(n693), .ZN(n692) );
  XOR2_X1 U746 ( .A(G113), .B(n692), .Z(G15) );
  NOR2_X1 U747 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U748 ( .A(KEYINPUT116), .B(n695), .Z(n696) );
  XNOR2_X1 U749 ( .A(G116), .B(n696), .ZN(G18) );
  XOR2_X1 U750 ( .A(KEYINPUT117), .B(KEYINPUT37), .Z(n699) );
  XNOR2_X1 U751 ( .A(G125), .B(n697), .ZN(n698) );
  XNOR2_X1 U752 ( .A(n699), .B(n698), .ZN(G27) );
  NAND2_X1 U753 ( .A1(n710), .A2(G469), .ZN(n701) );
  XOR2_X1 U754 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n700) );
  XNOR2_X1 U755 ( .A(n701), .B(n700), .ZN(n703) );
  XNOR2_X1 U756 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U757 ( .A1(n704), .A2(n717), .ZN(G54) );
  NAND2_X1 U758 ( .A1(n710), .A2(G475), .ZN(n707) );
  XOR2_X1 U759 ( .A(n705), .B(KEYINPUT59), .Z(n706) );
  XNOR2_X1 U760 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X2 U761 ( .A1(n708), .A2(n717), .ZN(n709) );
  XNOR2_X1 U762 ( .A(n709), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U763 ( .A1(n710), .A2(G478), .ZN(n712) );
  XNOR2_X1 U764 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U765 ( .A1(n717), .A2(n713), .ZN(G63) );
  NAND2_X1 U766 ( .A1(n710), .A2(G217), .ZN(n715) );
  XNOR2_X1 U767 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U768 ( .A1(n717), .A2(n716), .ZN(G66) );
  NAND2_X1 U769 ( .A1(n349), .A2(n732), .ZN(n721) );
  NAND2_X1 U770 ( .A1(G953), .A2(G224), .ZN(n718) );
  XNOR2_X1 U771 ( .A(KEYINPUT61), .B(n718), .ZN(n719) );
  NAND2_X1 U772 ( .A1(n719), .A2(G898), .ZN(n720) );
  NAND2_X1 U773 ( .A1(n721), .A2(n720), .ZN(n728) );
  XNOR2_X1 U774 ( .A(n722), .B(KEYINPUT126), .ZN(n723) );
  XNOR2_X1 U775 ( .A(n724), .B(n723), .ZN(n726) );
  NOR2_X1 U776 ( .A1(G898), .A2(n732), .ZN(n725) );
  NOR2_X1 U777 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U778 ( .A(n728), .B(n727), .ZN(G69) );
  XNOR2_X1 U779 ( .A(n730), .B(n729), .ZN(n734) );
  INV_X1 U780 ( .A(n734), .ZN(n731) );
  XOR2_X1 U781 ( .A(n731), .B(n628), .Z(n733) );
  NAND2_X1 U782 ( .A1(n733), .A2(n732), .ZN(n738) );
  XOR2_X1 U783 ( .A(G227), .B(n734), .Z(n735) );
  NAND2_X1 U784 ( .A1(n735), .A2(G900), .ZN(n736) );
  NAND2_X1 U785 ( .A1(n736), .A2(G953), .ZN(n737) );
  NAND2_X1 U786 ( .A1(n738), .A2(n737), .ZN(G72) );
  XOR2_X1 U787 ( .A(G134), .B(n739), .Z(G36) );
  XNOR2_X1 U788 ( .A(G137), .B(n740), .ZN(n741) );
  XNOR2_X1 U789 ( .A(n741), .B(KEYINPUT127), .ZN(G39) );
  XOR2_X1 U790 ( .A(n742), .B(G122), .Z(G24) );
  XNOR2_X1 U791 ( .A(G101), .B(n743), .ZN(G3) );
  XOR2_X1 U792 ( .A(G131), .B(n744), .Z(G33) );
endmodule

