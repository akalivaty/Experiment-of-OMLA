//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G116), .ZN(new_n209));
  INV_X1    g0009(.A(G270), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G68), .A2(G238), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G107), .A2(G264), .ZN(new_n214));
  AND3_X1   g0014(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(KEYINPUT67), .B(G77), .Z(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n206), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n202), .A2(G50), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR3_X1   g0029(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(KEYINPUT65), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n231), .B1(new_n206), .B2(G13), .ZN(new_n232));
  INV_X1    g0032(.A(G13), .ZN(new_n233));
  NAND4_X1  g0033(.A1(new_n233), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n235), .B(G250), .C1(G257), .C2(G264), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT66), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT0), .ZN(new_n238));
  NOR3_X1   g0038(.A1(new_n226), .A2(new_n230), .A3(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n210), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT68), .B(G264), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XNOR2_X1  g0043(.A(G238), .B(G244), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n219), .ZN(new_n245));
  XOR2_X1   g0045(.A(KEYINPUT2), .B(G226), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n243), .B(new_n247), .Z(G358));
  XOR2_X1   g0048(.A(G50), .B(G58), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT69), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G68), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G87), .B(G97), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G107), .B(G116), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n253), .B(new_n254), .Z(new_n255));
  XOR2_X1   g0055(.A(new_n252), .B(new_n255), .Z(G351));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n258));
  INV_X1    g0058(.A(G274), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G97), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n266), .B1(G232), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G226), .A2(G1698), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n261), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n229), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n260), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT13), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  INV_X1    g0077(.A(G45), .ZN(new_n278));
  AOI21_X1  g0078(.A(G1), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT70), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n258), .A2(KEYINPUT70), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(new_n273), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT73), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n281), .A2(new_n273), .A3(new_n282), .A4(KEYINPUT73), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(G238), .A3(new_n286), .ZN(new_n287));
  AND3_X1   g0087(.A1(new_n275), .A2(new_n276), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n276), .B1(new_n275), .B2(new_n287), .ZN(new_n289));
  OAI21_X1  g0089(.A(G169), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT14), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n288), .A2(new_n289), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G179), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT14), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n294), .B(G169), .C1(new_n288), .C2(new_n289), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n291), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n263), .A2(G20), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n297), .A2(G77), .B1(new_n298), .B2(G50), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(new_n228), .B2(G68), .ZN(new_n300));
  NAND3_X1  g0100(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(KEYINPUT71), .A3(new_n229), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(KEYINPUT71), .B1(new_n301), .B2(new_n229), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT11), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n301), .A2(new_n229), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n228), .A2(G1), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n306), .A2(new_n307), .B1(G68), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n300), .A2(new_n305), .A3(KEYINPUT11), .ZN(new_n312));
  INV_X1    g0112(.A(G68), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n257), .A2(new_n313), .A3(G13), .A4(G20), .ZN(new_n314));
  OAI21_X1  g0114(.A(KEYINPUT12), .B1(new_n314), .B2(KEYINPUT74), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(KEYINPUT74), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n315), .B(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n311), .A2(new_n312), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT75), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT75), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n311), .A2(new_n320), .A3(new_n312), .A4(new_n317), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n296), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(G200), .B1(new_n288), .B2(new_n289), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n292), .A2(G190), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT76), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n296), .A2(new_n323), .B1(new_n326), .B2(new_n327), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT76), .ZN(new_n333));
  INV_X1    g0133(.A(new_n298), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT8), .B(G58), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n222), .A2(new_n228), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XOR2_X1   g0136(.A(KEYINPUT15), .B(G87), .Z(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n297), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n308), .B1(new_n336), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n310), .A2(G77), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n341), .B(new_n342), .C1(new_n221), .C2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n260), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n283), .B2(new_n223), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT72), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n266), .A2(G238), .A3(G1698), .ZN(new_n349));
  INV_X1    g0149(.A(G107), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n266), .A2(new_n267), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n349), .B1(new_n350), .B2(new_n266), .C1(new_n351), .C2(new_n219), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n274), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n346), .A2(new_n347), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n348), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n344), .B1(new_n355), .B2(G200), .ZN(new_n356));
  INV_X1    g0156(.A(G190), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n356), .B1(new_n357), .B2(new_n355), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n331), .A2(new_n333), .A3(new_n358), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n283), .A2(new_n217), .ZN(new_n360));
  NOR2_X1   g0160(.A1(G222), .A2(G1698), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n267), .A2(G223), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n266), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(new_n274), .C1(new_n221), .C2(new_n266), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n360), .A2(new_n345), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G169), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n305), .A2(new_n309), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G50), .ZN(new_n369));
  INV_X1    g0169(.A(new_n343), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n216), .ZN(new_n371));
  INV_X1    g0171(.A(G150), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n335), .A2(new_n339), .B1(new_n372), .B2(new_n334), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n228), .B1(new_n201), .B2(new_n216), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n305), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n369), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n367), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G179), .ZN(new_n378));
  INV_X1    g0178(.A(new_n365), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(G190), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT9), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n365), .A2(G200), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n369), .A2(KEYINPUT9), .A3(new_n371), .A4(new_n375), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n381), .A2(new_n383), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  OR2_X1    g0186(.A1(new_n386), .A2(KEYINPUT10), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(KEYINPUT10), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n380), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n355), .A2(new_n366), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n390), .B(new_n344), .C1(G179), .C2(new_n355), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g0192(.A1(KEYINPUT3), .A2(G33), .ZN(new_n393));
  NOR2_X1   g0193(.A1(KEYINPUT3), .A2(G33), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT7), .B1(new_n395), .B2(new_n228), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  NOR4_X1   g0197(.A1(new_n393), .A2(new_n394), .A3(new_n397), .A4(G20), .ZN(new_n398));
  OAI21_X1  g0198(.A(G68), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n298), .A2(G159), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G58), .A2(G68), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n202), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G20), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n399), .A2(new_n400), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT16), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n399), .A2(KEYINPUT16), .A3(new_n400), .A4(new_n403), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n406), .A2(new_n308), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n335), .A2(new_n343), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n368), .B2(new_n335), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n410), .A2(KEYINPUT77), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(KEYINPUT77), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n408), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n345), .B1(new_n283), .B2(new_n219), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n217), .A2(G1698), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n266), .B(new_n415), .C1(G223), .C2(G1698), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G87), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n273), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G179), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n366), .B2(new_n419), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n413), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(KEYINPUT78), .A2(KEYINPUT18), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT78), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT18), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n422), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n408), .A2(new_n411), .A3(new_n412), .ZN(new_n428));
  INV_X1    g0228(.A(new_n419), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(new_n357), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(G200), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n428), .A2(KEYINPUT17), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT17), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n408), .A2(new_n432), .A3(new_n411), .A4(new_n412), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n434), .B1(new_n435), .B2(new_n430), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n413), .A2(new_n424), .A3(new_n425), .A4(new_n421), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n427), .A2(new_n433), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n392), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n359), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(G244), .B(new_n267), .C1(new_n393), .C2(new_n394), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT80), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n443), .A2(KEYINPUT4), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n266), .A2(G244), .A3(new_n267), .A4(new_n444), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n266), .A2(G250), .A3(G1698), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G283), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n274), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n278), .A2(G1), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n277), .A2(KEYINPUT5), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT5), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G41), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(new_n259), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n457), .A2(new_n273), .A3(G257), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n452), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT81), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n446), .A2(new_n447), .A3(new_n450), .A4(new_n449), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n460), .B1(new_n465), .B2(new_n274), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(KEYINPUT81), .A3(new_n459), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n464), .A2(new_n366), .A3(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n370), .A2(G97), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n343), .B1(G1), .B2(new_n263), .ZN(new_n471));
  INV_X1    g0271(.A(new_n304), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n471), .B1(new_n472), .B2(new_n302), .ZN(new_n473));
  INV_X1    g0273(.A(G97), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT79), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n309), .A2(G13), .B1(new_n257), .B2(G33), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n303), .B2(new_n304), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n469), .B1(new_n478), .B2(G97), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT79), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT6), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n483), .A2(new_n474), .A3(G107), .ZN(new_n484));
  XNOR2_X1  g0284(.A(G97), .B(G107), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G77), .ZN(new_n487));
  OAI22_X1  g0287(.A1(new_n486), .A2(new_n228), .B1(new_n487), .B2(new_n334), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n397), .B1(new_n266), .B2(G20), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n395), .A2(KEYINPUT7), .A3(new_n228), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n350), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n308), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  AOI211_X1 g0292(.A(new_n458), .B(new_n460), .C1(new_n465), .C2(new_n274), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n482), .A2(new_n492), .B1(new_n493), .B2(new_n378), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n468), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n257), .A2(new_n350), .A3(G13), .A4(G20), .ZN(new_n496));
  XOR2_X1   g0296(.A(new_n496), .B(KEYINPUT25), .Z(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n228), .B(G87), .C1(new_n393), .C2(new_n394), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT22), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT22), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n266), .A2(new_n501), .A3(new_n228), .A4(G87), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n297), .A2(G116), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT23), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n505), .A2(new_n228), .A3(G107), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT23), .B1(new_n350), .B2(G20), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  AND4_X1   g0309(.A1(KEYINPUT24), .A2(new_n503), .A3(new_n504), .A4(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n508), .B1(new_n500), .B2(new_n502), .ZN(new_n511));
  AOI21_X1  g0311(.A(KEYINPUT24), .B1(new_n511), .B2(new_n504), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n498), .B1(new_n513), .B2(new_n308), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n266), .A2(G257), .A3(G1698), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G294), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n515), .B(new_n516), .C1(new_n351), .C2(new_n208), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n274), .ZN(new_n518));
  XNOR2_X1  g0318(.A(KEYINPUT5), .B(G41), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(new_n453), .B1(new_n271), .B2(new_n272), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G264), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n518), .A2(new_n459), .A3(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(new_n357), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n473), .A2(G107), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n522), .A2(G200), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n514), .A2(new_n524), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT19), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n297), .A2(new_n528), .A3(G97), .ZN(new_n529));
  NOR2_X1   g0329(.A1(G97), .A2(G107), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n530), .A2(new_n207), .B1(new_n261), .B2(new_n228), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n529), .B1(new_n531), .B2(new_n528), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n228), .B(G68), .C1(new_n393), .C2(new_n394), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT82), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT82), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n266), .A2(new_n535), .A3(new_n228), .A4(G68), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n532), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n537), .A2(new_n308), .B1(new_n370), .B2(new_n338), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n257), .A2(G45), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(new_n259), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n272), .ZN(new_n542));
  OAI211_X1 g0342(.A(G250), .B(new_n539), .C1(new_n542), .C2(new_n229), .ZN(new_n543));
  INV_X1    g0343(.A(G238), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n267), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n223), .A2(G1698), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n545), .B(new_n546), .C1(new_n393), .C2(new_n394), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G116), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n541), .B(new_n543), .C1(new_n549), .C2(new_n273), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G200), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n273), .B1(new_n547), .B2(new_n548), .ZN(new_n552));
  INV_X1    g0352(.A(new_n543), .ZN(new_n553));
  NOR3_X1   g0353(.A1(new_n552), .A2(new_n553), .A3(new_n540), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G190), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n473), .A2(G87), .ZN(new_n556));
  AND4_X1   g0356(.A1(new_n538), .A2(new_n551), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n537), .A2(new_n308), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n338), .A2(new_n370), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n473), .A2(new_n337), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT83), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT83), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n538), .A2(new_n563), .A3(new_n560), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n554), .A2(G169), .ZN(new_n566));
  NOR4_X1   g0366(.A1(new_n552), .A2(new_n553), .A3(G179), .A4(new_n540), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n557), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  AND4_X1   g0369(.A1(KEYINPUT81), .A2(new_n452), .A3(new_n459), .A4(new_n461), .ZN(new_n570));
  AOI21_X1  g0370(.A(KEYINPUT81), .B1(new_n466), .B2(new_n459), .ZN(new_n571));
  OAI21_X1  g0371(.A(G190), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n479), .A2(new_n480), .ZN(new_n573));
  AOI211_X1 g0373(.A(KEYINPUT79), .B(new_n469), .C1(new_n478), .C2(G97), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n492), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(G200), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n466), .B2(new_n459), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n572), .A2(new_n578), .ZN(new_n579));
  AND4_X1   g0379(.A1(new_n495), .A2(new_n527), .A3(new_n569), .A4(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n301), .A2(new_n229), .B1(G20), .B2(new_n209), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n450), .B(new_n228), .C1(G33), .C2(new_n474), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT20), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n584), .A2(KEYINPUT85), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n585), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n581), .A2(new_n587), .A3(new_n582), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n586), .A2(new_n588), .B1(KEYINPUT85), .B2(new_n584), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n477), .A2(G116), .ZN(new_n590));
  OAI22_X1  g0390(.A1(new_n590), .A2(new_n308), .B1(G116), .B2(new_n343), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n589), .A2(KEYINPUT86), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT86), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n584), .A2(KEYINPUT85), .ZN(new_n594));
  INV_X1    g0394(.A(new_n588), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n587), .B1(new_n581), .B2(new_n582), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n471), .A2(new_n209), .ZN(new_n598));
  INV_X1    g0398(.A(new_n308), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n598), .A2(new_n599), .B1(new_n209), .B2(new_n370), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n593), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n592), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(G257), .B(new_n267), .C1(new_n393), .C2(new_n394), .ZN(new_n603));
  OAI211_X1 g0403(.A(G264), .B(G1698), .C1(new_n393), .C2(new_n394), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n264), .A2(G303), .A3(new_n265), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n274), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n520), .A2(G270), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(new_n459), .A3(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT84), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n606), .A2(new_n274), .B1(new_n520), .B2(G270), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(KEYINPUT84), .A3(new_n459), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n614), .A2(KEYINPUT21), .A3(G169), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n609), .A2(new_n378), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n602), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT21), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n609), .A2(new_n610), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT84), .B1(new_n612), .B2(new_n459), .ZN(new_n621));
  OAI21_X1  g0421(.A(G169), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n619), .B1(new_n622), .B2(new_n602), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(KEYINPUT87), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT86), .B1(new_n589), .B2(new_n591), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n597), .A2(new_n593), .A3(new_n600), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n627), .A2(new_n614), .A3(G169), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT87), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(new_n629), .A3(new_n619), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n618), .B1(new_n624), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n614), .A2(G200), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n632), .B(new_n602), .C1(new_n357), .C2(new_n614), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n503), .A2(new_n504), .A3(new_n509), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT24), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n511), .A2(KEYINPUT24), .A3(new_n504), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(new_n308), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n638), .A2(new_n525), .A3(new_n497), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n522), .A2(new_n366), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n518), .A2(new_n521), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(new_n378), .A3(new_n459), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT88), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n639), .A2(KEYINPUT88), .A3(new_n640), .A4(new_n642), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n580), .A2(new_n631), .A3(new_n633), .A4(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n441), .A2(new_n648), .ZN(G372));
  NAND2_X1  g0449(.A1(new_n324), .A2(new_n391), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n433), .A2(new_n436), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n650), .A2(new_n328), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g0453(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n413), .A2(KEYINPUT90), .A3(new_n421), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT90), .B1(new_n413), .B2(new_n421), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT90), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n422), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n661), .A2(new_n656), .A3(new_n654), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n653), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n387), .A2(new_n388), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n380), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT89), .B1(new_n550), .B2(new_n366), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n667), .B1(new_n562), .B2(new_n564), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT89), .B1(new_n566), .B2(new_n567), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n557), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n670), .A2(new_n527), .A3(new_n495), .A4(new_n579), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n631), .B2(new_n643), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n565), .A2(new_n568), .ZN(new_n673));
  INV_X1    g0473(.A(new_n557), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n673), .A2(new_n468), .A3(new_n674), .A4(new_n494), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT26), .ZN(new_n676));
  INV_X1    g0476(.A(new_n495), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT26), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(new_n670), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n667), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n561), .A2(KEYINPUT83), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n563), .B1(new_n538), .B2(new_n560), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n680), .B(new_n669), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n676), .A2(new_n679), .A3(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n672), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n666), .B1(new_n441), .B2(new_n685), .ZN(G369));
  AND2_X1   g0486(.A1(new_n645), .A2(new_n646), .ZN(new_n687));
  INV_X1    g0487(.A(new_n526), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n639), .A2(new_n688), .A3(new_n523), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n233), .A2(G1), .A3(G20), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT92), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT27), .ZN(new_n693));
  OR3_X1    g0493(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(G213), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n695), .B1(new_n691), .B2(new_n693), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n692), .B1(new_n691), .B2(new_n693), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n694), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT93), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(KEYINPUT93), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n702), .A2(G343), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n639), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT94), .Z(new_n705));
  NAND2_X1  g0505(.A1(new_n690), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n703), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(new_n643), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n615), .A2(new_n617), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n627), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n628), .A2(new_n629), .A3(new_n619), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n629), .B1(new_n628), .B2(new_n619), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n707), .A2(new_n602), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(G330), .A3(new_n633), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n710), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n631), .A2(new_n703), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n690), .A2(new_n705), .A3(new_n721), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n643), .A2(new_n703), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n720), .A2(new_n724), .ZN(G399));
  INV_X1    g0525(.A(new_n235), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G41), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR4_X1   g0528(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(G1), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n227), .B2(new_n728), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT28), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT29), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n570), .A2(new_n571), .A3(G169), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n575), .B1(G179), .B2(new_n462), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n357), .B1(new_n464), .B2(new_n467), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n482), .B(new_n492), .C1(new_n493), .C2(new_n576), .ZN(new_n737));
  OAI22_X1  g0537(.A1(new_n734), .A2(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n683), .A2(new_n674), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n738), .A2(new_n689), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n687), .B2(new_n715), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT26), .B1(new_n739), .B2(new_n495), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n683), .B1(new_n675), .B2(KEYINPUT26), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n733), .B1(new_n745), .B2(new_n707), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n707), .B1(new_n672), .B2(new_n684), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(KEYINPUT29), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT30), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n641), .B(new_n554), .C1(new_n570), .C2(new_n571), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n750), .B1(new_n751), .B2(new_n617), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n550), .B1(new_n464), .B2(new_n467), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n753), .A2(KEYINPUT30), .A3(new_n641), .A4(new_n616), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n493), .B1(new_n611), .B2(new_n613), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n755), .A2(new_n378), .A3(new_n522), .A4(new_n550), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n752), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n703), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT31), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n757), .A2(KEYINPUT31), .A3(new_n703), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n760), .B(new_n761), .C1(new_n648), .C2(new_n703), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G330), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n749), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n732), .B1(new_n765), .B2(G1), .ZN(G364));
  NOR2_X1   g0566(.A1(new_n233), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n257), .B1(new_n767), .B2(G45), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n727), .A2(new_n769), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n717), .A2(new_n633), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n770), .B1(new_n771), .B2(G330), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(G330), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT95), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n771), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n726), .A2(G116), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n271), .B1(new_n228), .B2(G169), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT96), .Z(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n777), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G355), .A2(new_n395), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n252), .A2(G45), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(G45), .B2(new_n227), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n785), .B1(new_n787), .B2(new_n395), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n780), .B(new_n784), .C1(new_n788), .C2(new_n726), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n378), .A2(new_n576), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT98), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n228), .A2(G190), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G329), .ZN(new_n795));
  INV_X1    g0595(.A(G326), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n228), .A2(new_n357), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n378), .A2(new_n576), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n795), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n798), .A2(new_n792), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(KEYINPUT33), .B(G317), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n378), .A2(G200), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n797), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G322), .ZN(new_n808));
  OAI21_X1  g0608(.A(G20), .B1(new_n791), .B2(new_n357), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G294), .ZN(new_n810));
  INV_X1    g0610(.A(G283), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n576), .A2(G179), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n792), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n805), .A2(new_n792), .ZN(new_n814));
  INV_X1    g0614(.A(G311), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n811), .A2(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n797), .A2(new_n812), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n266), .B(new_n816), .C1(G303), .C2(new_n818), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n804), .A2(new_n808), .A3(new_n810), .A4(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n799), .ZN(new_n821));
  INV_X1    g0621(.A(new_n814), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G50), .A2(new_n821), .B1(new_n822), .B2(new_n221), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n218), .B2(new_n806), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT97), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n809), .A2(G97), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n802), .A2(G68), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n794), .A2(G159), .ZN(new_n828));
  XNOR2_X1  g0628(.A(KEYINPUT99), .B(KEYINPUT32), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n828), .A2(new_n829), .B1(G87), .B2(new_n818), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n825), .A2(new_n826), .A3(new_n827), .A4(new_n830), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n266), .B1(new_n350), .B2(new_n813), .C1(new_n828), .C2(new_n829), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n820), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n783), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n789), .A2(new_n834), .A3(new_n770), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT100), .Z(new_n836));
  AOI22_X1  g0636(.A1(new_n772), .A2(new_n774), .B1(new_n779), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(G396));
  NOR2_X1   g0638(.A1(new_n391), .A2(new_n703), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n703), .A2(new_n344), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n358), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n839), .B1(new_n841), .B2(new_n391), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n747), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n707), .B(new_n842), .C1(new_n672), .C2(new_n684), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(G330), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n757), .A2(KEYINPUT31), .A3(new_n703), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT31), .B1(new_n757), .B2(new_n703), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n687), .A2(new_n715), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n851), .A2(new_n633), .A3(new_n580), .A4(new_n707), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n847), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n846), .B(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n727), .B2(new_n769), .ZN(new_n855));
  INV_X1    g0655(.A(new_n776), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n843), .A2(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(G143), .A2(new_n807), .B1(new_n802), .B2(G150), .ZN(new_n858));
  INV_X1    g0658(.A(G137), .ZN(new_n859));
  INV_X1    g0659(.A(G159), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n858), .B1(new_n859), .B2(new_n799), .C1(new_n860), .C2(new_n814), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT34), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n266), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n794), .A2(G132), .ZN(new_n865));
  INV_X1    g0665(.A(new_n813), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G50), .A2(new_n818), .B1(new_n866), .B2(G68), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n863), .B(new_n868), .C1(G58), .C2(new_n809), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n801), .A2(new_n811), .B1(new_n814), .B2(new_n209), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n266), .B(new_n870), .C1(G294), .C2(new_n807), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n794), .A2(G311), .ZN(new_n872));
  AOI22_X1  g0672(.A1(G107), .A2(new_n818), .B1(new_n866), .B2(G87), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n871), .A2(new_n826), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(G303), .B2(new_n821), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n783), .B1(new_n869), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n782), .A2(new_n776), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n877), .B(KEYINPUT101), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n487), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n857), .A2(new_n770), .A3(new_n876), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n855), .A2(new_n880), .ZN(G384));
  NAND2_X1  g0681(.A1(new_n440), .A2(new_n762), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n882), .B(KEYINPUT105), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n406), .A2(new_n305), .A3(new_n407), .ZN(new_n884));
  INV_X1    g0684(.A(new_n410), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n702), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n438), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n421), .B1(new_n884), .B2(new_n885), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n886), .B(new_n889), .C1(new_n430), .C2(new_n435), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  AND4_X1   g0691(.A1(new_n411), .A2(new_n408), .A3(new_n412), .A4(new_n432), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n431), .ZN(new_n893));
  XOR2_X1   g0693(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n413), .A2(new_n702), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n893), .A2(new_n422), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n888), .A2(KEYINPUT38), .A3(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT38), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n651), .B1(new_n659), .B2(new_n662), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n657), .A2(new_n658), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n892), .A2(new_n431), .B1(new_n413), .B2(new_n702), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n895), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n897), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n901), .A2(new_n896), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n899), .B1(new_n900), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n323), .A2(new_n703), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n329), .A2(new_n909), .B1(new_n324), .B2(new_n707), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n762), .A2(new_n842), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT40), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n843), .B1(new_n850), .B2(new_n852), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n888), .A2(new_n898), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n900), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n888), .A2(new_n898), .A3(KEYINPUT38), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT40), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n913), .A2(new_n917), .A3(new_n918), .A4(new_n910), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n912), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n883), .B(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(G330), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n324), .A2(new_n707), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n332), .B2(new_n908), .ZN(new_n924));
  INV_X1    g0724(.A(new_n839), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n924), .B1(new_n845), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n917), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n663), .A2(new_n702), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT104), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT39), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n657), .A2(new_n658), .A3(new_n655), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n654), .B1(new_n661), .B2(new_n656), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n652), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n896), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n661), .A2(new_n893), .A3(new_n656), .A4(new_n896), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n894), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n936), .A2(new_n937), .B1(new_n897), .B2(new_n939), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n933), .B(new_n916), .C1(new_n940), .C2(KEYINPUT38), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT38), .B1(new_n888), .B2(new_n898), .ZN(new_n942));
  OAI21_X1  g0742(.A(KEYINPUT39), .B1(new_n899), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n324), .A2(new_n703), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n927), .A2(KEYINPUT104), .A3(new_n929), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n932), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n440), .B1(new_n746), .B2(new_n748), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n949), .A2(new_n666), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n948), .B(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n922), .B(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n257), .B2(new_n767), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT35), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n228), .B(new_n229), .C1(new_n486), .C2(new_n954), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n955), .B(G116), .C1(new_n954), .C2(new_n486), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT36), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n202), .A2(G50), .A3(new_n401), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n222), .A2(new_n958), .B1(G50), .B2(new_n313), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n959), .A2(G1), .A3(new_n233), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT102), .Z(new_n961));
  NAND3_X1  g0761(.A1(new_n953), .A2(new_n957), .A3(new_n961), .ZN(G367));
  AOI21_X1  g0762(.A(new_n395), .B1(new_n821), .B2(G143), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n222), .B2(new_n813), .ZN(new_n964));
  INV_X1    g0764(.A(new_n809), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n965), .A2(new_n313), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(G58), .B2(new_n818), .ZN(new_n967));
  AOI22_X1  g0767(.A1(G159), .A2(new_n802), .B1(new_n822), .B2(G50), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n967), .B(new_n968), .C1(new_n372), .C2(new_n806), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n964), .B(new_n969), .C1(G137), .C2(new_n794), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n818), .A2(KEYINPUT46), .A3(G116), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n802), .A2(G294), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT46), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n817), .B2(new_n209), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT110), .ZN(new_n976));
  INV_X1    g0776(.A(G303), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n395), .B1(new_n814), .B2(new_n811), .C1(new_n977), .C2(new_n806), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n965), .A2(new_n350), .ZN(new_n979));
  INV_X1    g0779(.A(new_n794), .ZN(new_n980));
  INV_X1    g0780(.A(G317), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n799), .A2(new_n815), .ZN(new_n983));
  OR4_X1    g0783(.A1(new_n978), .A2(new_n979), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n976), .B(new_n984), .C1(G97), .C2(new_n866), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n970), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT47), .Z(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n783), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n707), .B1(new_n538), .B2(new_n556), .ZN(new_n989));
  INV_X1    g0789(.A(new_n683), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n739), .B2(new_n989), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n992), .A2(new_n778), .ZN(new_n993));
  INV_X1    g0793(.A(new_n243), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n235), .A2(new_n395), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n784), .B1(new_n235), .B2(new_n338), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n988), .A2(new_n770), .A3(new_n993), .A4(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n722), .A2(new_n723), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n677), .A2(new_n703), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n703), .A2(new_n575), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n1000), .A2(new_n579), .A3(new_n495), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n998), .A2(new_n1003), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n1004), .A2(KEYINPUT45), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1004), .A2(KEYINPUT45), .ZN(new_n1006));
  AOI21_X1  g0806(.A(KEYINPUT44), .B1(new_n998), .B2(new_n1003), .ZN(new_n1007));
  AND3_X1   g0807(.A1(new_n998), .A2(KEYINPUT44), .A3(new_n1003), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n1005), .A2(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1009), .A2(KEYINPUT109), .A3(new_n720), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1004), .B(KEYINPUT45), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1008), .A2(new_n1007), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n720), .A2(KEYINPUT109), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT109), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n719), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1010), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT108), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n722), .B1(new_n709), .B2(new_n721), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n719), .B1(new_n718), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n765), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n718), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n720), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(KEYINPUT108), .B1(new_n1023), .B2(new_n764), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n765), .B1(new_n1017), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n727), .B(KEYINPUT41), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n769), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n719), .A2(new_n1002), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT107), .Z(new_n1031));
  XNOR2_X1  g0831(.A(new_n1029), .B(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n722), .A2(new_n1003), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1034), .B(new_n1035), .Z(new_n1036));
  AOI21_X1  g0836(.A(new_n677), .B1(new_n687), .B2(new_n579), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1037), .A2(new_n703), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1033), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1032), .B(new_n1039), .Z(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n997), .B1(new_n1028), .B2(new_n1041), .ZN(G387));
  INV_X1    g0842(.A(KEYINPUT112), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n1025), .B2(new_n727), .ZN(new_n1044));
  AOI211_X1 g0844(.A(KEYINPUT112), .B(new_n728), .C1(new_n1021), .C2(new_n1024), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n765), .A2(new_n1020), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1020), .A2(new_n769), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n710), .A2(new_n777), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n266), .B1(new_n801), .B2(new_n335), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n794), .A2(G150), .B1(G97), .B2(new_n866), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n818), .A2(new_n221), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n822), .A2(G68), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n809), .A2(new_n337), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1051), .B(new_n1056), .C1(G159), .C2(new_n821), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n216), .B2(new_n806), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n809), .A2(G283), .B1(G294), .B2(new_n818), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT111), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G311), .A2(new_n802), .B1(new_n807), .B2(G317), .ZN(new_n1061));
  INV_X1    g0861(.A(G322), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1061), .B1(new_n977), .B2(new_n814), .C1(new_n1062), .C2(new_n799), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1060), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT49), .Z(new_n1068));
  OAI221_X1 g0868(.A(new_n395), .B1(new_n209), .B2(new_n813), .C1(new_n980), .C2(new_n796), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1058), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n783), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n726), .A2(G107), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n247), .A2(new_n278), .A3(new_n266), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n335), .A2(G50), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n278), .B1(new_n1075), .B2(KEYINPUT50), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT50), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1074), .A2(new_n1077), .B1(new_n313), .B2(new_n487), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n395), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1073), .B1(new_n729), .B2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n784), .B(new_n1072), .C1(new_n1080), .C2(new_n726), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1050), .A2(new_n770), .A3(new_n1071), .A4(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1049), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1048), .A2(new_n1084), .ZN(G393));
  NAND2_X1  g0885(.A1(new_n1003), .A2(new_n777), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n784), .B1(new_n474), .B2(new_n235), .C1(new_n255), .C2(new_n995), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(G283), .A2(new_n818), .B1(new_n866), .B2(G107), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n266), .B1(new_n822), .B2(G294), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT52), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n799), .A2(new_n981), .B1(new_n806), .B2(new_n815), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1088), .B(new_n1089), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1090), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n980), .B2(new_n1062), .C1(new_n209), .C2(new_n965), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1092), .B(new_n1094), .C1(G303), .C2(new_n802), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n799), .A2(new_n372), .B1(new_n806), .B2(new_n860), .ZN(new_n1096));
  XOR2_X1   g0896(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n1097));
  OR2_X1    g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n794), .A2(G143), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1098), .A2(new_n1099), .A3(new_n266), .A4(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G68), .A2(new_n818), .B1(new_n866), .B2(G87), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1102), .B1(new_n335), .B2(new_n814), .C1(new_n965), .C2(new_n487), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1101), .B(new_n1103), .C1(G50), .C2(new_n802), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n783), .B1(new_n1095), .B2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1086), .A2(new_n770), .A3(new_n1087), .A4(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n1017), .B2(new_n768), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1010), .A2(new_n1016), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1108), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n728), .B1(new_n1017), .B2(new_n1025), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1107), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(G390));
  AOI22_X1  g0912(.A1(new_n794), .A2(G294), .B1(G87), .B2(new_n818), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n350), .B2(new_n801), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n965), .A2(new_n487), .B1(new_n313), .B2(new_n813), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n806), .A2(new_n209), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n395), .B1(new_n814), .B2(new_n474), .C1(new_n811), .C2(new_n799), .ZN(new_n1117));
  NOR4_X1   g0917(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n809), .A2(G159), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n817), .A2(new_n372), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT53), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n807), .A2(G132), .ZN(new_n1123));
  XOR2_X1   g0923(.A(KEYINPUT54), .B(G143), .Z(new_n1124));
  AOI22_X1  g0924(.A1(G137), .A2(new_n802), .B1(new_n822), .B2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1119), .A2(new_n1122), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(G125), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n980), .A2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n813), .A2(new_n216), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n395), .B1(new_n821), .B2(G128), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n1121), .B2(new_n1120), .ZN(new_n1131));
  NOR4_X1   g0931(.A1(new_n1126), .A2(new_n1128), .A3(new_n1129), .A4(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n783), .B1(new_n1118), .B2(new_n1132), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n727), .B(new_n769), .C1(new_n878), .C2(new_n335), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT117), .Z(new_n1135));
  OAI211_X1 g0935(.A(new_n1133), .B(new_n1135), .C1(new_n944), .C2(new_n776), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT118), .Z(new_n1137));
  NOR2_X1   g0937(.A1(new_n926), .A2(new_n945), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n945), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n936), .A2(new_n937), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n939), .A2(new_n897), .ZN(new_n1141));
  AOI21_X1  g0941(.A(KEYINPUT38), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1139), .B1(new_n1142), .B2(new_n899), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n841), .A2(new_n391), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n745), .A2(new_n707), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n924), .B1(new_n1145), .B2(new_n925), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n944), .A2(new_n1138), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  AND4_X1   g0947(.A1(G330), .A2(new_n762), .A3(new_n842), .A4(new_n910), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n941), .B(new_n943), .C1(new_n945), .C2(new_n926), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n853), .A2(new_n842), .A3(new_n910), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(new_n1146), .C2(new_n1143), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1149), .A2(new_n769), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1137), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n440), .A2(G330), .A3(new_n762), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n949), .A2(new_n1156), .A3(new_n666), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n845), .A2(new_n925), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n910), .B1(new_n853), .B2(new_n842), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1158), .B1(new_n1159), .B2(new_n1148), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n924), .B1(new_n763), .B2(new_n843), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n631), .A2(new_n647), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n743), .B1(new_n1162), .B2(new_n740), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n703), .B1(new_n1163), .B2(new_n742), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n839), .B1(new_n1164), .B2(new_n1144), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1161), .A2(new_n1165), .A3(new_n1151), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1157), .B1(new_n1160), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1167), .A2(new_n1149), .A3(new_n1152), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n727), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(KEYINPUT114), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT114), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1168), .A2(new_n1171), .A3(new_n727), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(KEYINPUT115), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1167), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT115), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1149), .A2(new_n1152), .A3(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(KEYINPUT116), .B1(new_n1173), .B2(new_n1179), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n1168), .A2(new_n1171), .A3(new_n727), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1171), .B1(new_n1168), .B2(new_n727), .ZN(new_n1182));
  OAI211_X1 g0982(.A(KEYINPUT116), .B(new_n1179), .C1(new_n1181), .C2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1155), .B1(new_n1180), .B2(new_n1184), .ZN(G378));
  NAND2_X1  g0985(.A1(new_n702), .A2(new_n376), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n389), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n389), .A2(new_n1186), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1189), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n920), .B2(G330), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n847), .B(new_n1192), .C1(new_n912), .C2(new_n919), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n948), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  AND3_X1   g0996(.A1(new_n762), .A2(new_n842), .A3(new_n910), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n916), .B1(new_n940), .B2(KEYINPUT38), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n918), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n918), .B1(new_n899), .B2(new_n942), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n911), .A2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(G330), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n1192), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT104), .B1(new_n927), .B2(new_n929), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n931), .B(new_n928), .C1(new_n926), .C2(new_n917), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1139), .B1(new_n941), .B2(new_n943), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n920), .A2(G330), .A3(new_n1193), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1203), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1196), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1157), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1168), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT57), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1210), .A2(KEYINPUT57), .A3(new_n1212), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1215), .A2(new_n727), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1210), .A2(new_n769), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n980), .A2(new_n811), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n806), .A2(new_n350), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n802), .A2(G97), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n822), .A2(new_n337), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1053), .A2(new_n1221), .A3(new_n1222), .A4(new_n277), .ZN(new_n1223));
  NOR4_X1   g1023(.A1(new_n966), .A2(new_n1219), .A3(new_n1220), .A4(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n866), .A2(G58), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n821), .A2(G116), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1224), .A2(new_n395), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT58), .Z(new_n1228));
  OAI21_X1  g1028(.A(new_n216), .B1(new_n393), .B2(G41), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n809), .A2(G150), .B1(G128), .B2(new_n807), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1124), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n1231), .A2(new_n817), .B1(new_n1127), .B2(new_n799), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G132), .B2(new_n802), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1230), .B(new_n1233), .C1(new_n859), .C2(new_n814), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n866), .A2(G159), .ZN(new_n1236));
  AOI21_X1  g1036(.A(G41), .B1(new_n794), .B2(G124), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1235), .A2(new_n263), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1229), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n783), .B1(new_n1228), .B2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n770), .B1(new_n877), .B2(G50), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT119), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1241), .B(new_n1243), .C1(new_n1193), .C2(new_n776), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n1244), .B(KEYINPUT120), .Z(new_n1245));
  NAND2_X1  g1045(.A1(new_n1218), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1217), .A2(new_n1247), .ZN(G375));
  NAND3_X1  g1048(.A1(new_n1160), .A2(new_n1157), .A3(new_n1166), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1176), .A2(new_n1027), .A3(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n768), .B1(new_n1160), .B2(new_n1166), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(G294), .A2(new_n821), .B1(new_n802), .B2(G116), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT121), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n395), .B1(new_n813), .B2(new_n487), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1055), .B(new_n1252), .C1(new_n1253), .C2(new_n1254), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n794), .A2(G303), .B1(new_n1254), .B2(new_n1253), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n1256), .B1(new_n350), .B2(new_n814), .C1(new_n811), .C2(new_n806), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1255), .B(new_n1257), .C1(G97), .C2(new_n818), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n395), .B1(new_n821), .B2(G132), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n802), .A2(new_n1124), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n822), .A2(G150), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1259), .A2(new_n1225), .A3(new_n1260), .A4(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n794), .A2(G128), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n1263), .B1(new_n859), .B2(new_n806), .C1(new_n965), .C2(new_n216), .ZN(new_n1264));
  AOI211_X1 g1064(.A(new_n1262), .B(new_n1264), .C1(G159), .C2(new_n818), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n783), .B1(new_n1258), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n924), .A2(new_n856), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n878), .A2(new_n313), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1267), .A2(new_n770), .A3(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1251), .B1(new_n1266), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1250), .A2(new_n1270), .ZN(G381));
  AND3_X1   g1071(.A1(new_n1210), .A2(KEYINPUT57), .A3(new_n1212), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT57), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1246), .B1(new_n1274), .B2(new_n727), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1154), .B1(new_n1173), .B2(new_n1179), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(new_n1277), .A2(G384), .A3(G381), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1027), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(new_n1109), .B2(new_n765), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1040), .B1(new_n1280), .B2(new_n769), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(new_n997), .A3(new_n1111), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1048), .A2(new_n837), .A3(new_n1084), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1278), .A2(new_n1283), .A3(new_n1285), .ZN(G407));
  OAI211_X1 g1086(.A(G407), .B(G213), .C1(G343), .C2(new_n1277), .ZN(G409));
  NOR2_X1   g1087(.A1(new_n695), .A2(G343), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(G378), .A2(new_n1275), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1218), .B(new_n1244), .C1(new_n1213), .C2(new_n1279), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1276), .A2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1288), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1288), .A2(G2897), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT60), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n728), .B1(new_n1249), .B2(new_n1296), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1297), .B(new_n1176), .C1(new_n1296), .C2(new_n1249), .ZN(new_n1298));
  AOI21_X1  g1098(.A(G384), .B1(new_n1298), .B2(new_n1270), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT122), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1298), .A2(new_n1270), .A3(G384), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1300), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1301), .B1(new_n1300), .B2(new_n1302), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1295), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  OR2_X1    g1105(.A1(new_n1304), .A2(new_n1295), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(KEYINPUT123), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT123), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1305), .A2(new_n1306), .A3(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1293), .A2(new_n1308), .A3(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1179), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT116), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1154), .B1(new_n1314), .B2(new_n1183), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1291), .B1(new_n1315), .B2(G375), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1288), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1316), .A2(new_n1317), .A3(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT63), .ZN(new_n1321));
  AOI21_X1  g1121(.A(KEYINPUT61), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(G387), .A2(G390), .ZN(new_n1323));
  OAI21_X1  g1123(.A(G396), .B1(new_n1047), .B2(new_n1083), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1284), .A2(new_n1324), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1323), .A2(new_n1325), .A3(new_n1282), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1325), .B1(new_n1323), .B2(new_n1282), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1292), .A2(KEYINPUT63), .A3(new_n1319), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1311), .A2(new_n1322), .A3(new_n1328), .A4(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT124), .ZN(new_n1331));
  AND3_X1   g1131(.A1(new_n1320), .A2(new_n1331), .A3(KEYINPUT62), .ZN(new_n1332));
  AOI21_X1  g1132(.A(KEYINPUT62), .B1(new_n1320), .B2(new_n1331), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT61), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1334), .B1(new_n1292), .B2(new_n1307), .ZN(new_n1335));
  NOR3_X1   g1135(.A1(new_n1332), .A2(new_n1333), .A3(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1330), .B1(new_n1336), .B2(new_n1328), .ZN(G405));
  INV_X1    g1137(.A(KEYINPUT127), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1338), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1323), .A2(new_n1282), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1325), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1323), .A2(new_n1325), .A3(new_n1282), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1342), .A2(KEYINPUT127), .A3(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1339), .A2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(G375), .A2(new_n1276), .ZN(new_n1346));
  AND2_X1   g1146(.A1(new_n1289), .A2(new_n1346), .ZN(new_n1347));
  AOI21_X1  g1147(.A(KEYINPUT126), .B1(new_n1319), .B2(KEYINPUT125), .ZN(new_n1348));
  OR2_X1    g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  AND2_X1   g1149(.A1(new_n1319), .A2(KEYINPUT126), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1347), .B1(new_n1348), .B2(new_n1350), .ZN(new_n1351));
  AND3_X1   g1151(.A1(new_n1345), .A2(new_n1349), .A3(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1345), .B1(new_n1349), .B2(new_n1351), .ZN(new_n1353));
  NOR2_X1   g1153(.A1(new_n1352), .A2(new_n1353), .ZN(G402));
endmodule


