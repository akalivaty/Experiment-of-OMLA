//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G214), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G131), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n189), .B(G143), .ZN(new_n193));
  INV_X1    g007(.A(G131), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n192), .A2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(G125), .B(G140), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT16), .ZN(new_n198));
  INV_X1    g012(.A(G140), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G125), .ZN(new_n200));
  OR2_X1    g014(.A1(new_n200), .A2(KEYINPUT16), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n198), .A2(G146), .A3(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT90), .B1(new_n197), .B2(KEYINPUT78), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT19), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT78), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT90), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(new_n204), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n203), .A2(new_n204), .B1(new_n197), .B2(new_n207), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n196), .B(new_n202), .C1(G146), .C2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G125), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G140), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n200), .A2(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(G146), .B1(new_n212), .B2(new_n205), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n197), .A2(KEYINPUT78), .ZN(new_n214));
  AOI22_X1  g028(.A1(new_n213), .A2(new_n214), .B1(G146), .B2(new_n212), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT89), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT18), .A2(G131), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n193), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NOR3_X1   g034(.A1(new_n193), .A2(KEYINPUT88), .A3(new_n218), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT88), .ZN(new_n222));
  INV_X1    g036(.A(new_n218), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n222), .B1(new_n191), .B2(new_n223), .ZN(new_n224));
  OAI22_X1  g038(.A1(new_n221), .A2(new_n224), .B1(new_n215), .B2(new_n216), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n209), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G113), .B(G122), .ZN(new_n227));
  INV_X1    g041(.A(G104), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n227), .B(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  OR2_X1    g045(.A1(new_n215), .A2(new_n216), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT88), .B1(new_n193), .B2(new_n218), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n191), .A2(new_n222), .A3(new_n223), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n232), .A2(new_n217), .A3(new_n235), .A4(new_n219), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT91), .ZN(new_n237));
  INV_X1    g051(.A(new_n202), .ZN(new_n238));
  AOI21_X1  g052(.A(G146), .B1(new_n198), .B2(new_n201), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n239), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(KEYINPUT91), .A3(new_n202), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT17), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n192), .A2(new_n195), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n191), .A2(KEYINPUT17), .A3(G131), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n240), .A2(new_n242), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n236), .A2(new_n246), .A3(new_n229), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n231), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(G475), .A2(G902), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT92), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT20), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G902), .ZN(new_n254));
  INV_X1    g068(.A(new_n247), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n229), .B1(new_n236), .B2(new_n246), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G475), .ZN(new_n258));
  INV_X1    g072(.A(new_n249), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n259), .B1(new_n231), .B2(new_n247), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT92), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT20), .B1(new_n260), .B2(KEYINPUT92), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n253), .B(new_n258), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(G116), .B(G122), .ZN(new_n266));
  INV_X1    g080(.A(G107), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G122), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT14), .B1(new_n269), .B2(G116), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n270), .B(KEYINPUT94), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT14), .ZN(new_n272));
  INV_X1    g086(.A(G116), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n273), .A3(G122), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n274), .B1(new_n273), .B2(G122), .ZN(new_n275));
  OAI21_X1  g089(.A(G107), .B1(new_n271), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(G128), .B(G143), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n277), .B(KEYINPUT93), .ZN(new_n278));
  INV_X1    g092(.A(G134), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n278), .A2(new_n279), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n268), .B(new_n276), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n278), .A2(new_n279), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n266), .B(new_n267), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n277), .A2(KEYINPUT13), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n190), .A2(G128), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n285), .B(G134), .C1(KEYINPUT13), .C2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n283), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(KEYINPUT9), .B(G234), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n289), .B(KEYINPUT80), .ZN(new_n290));
  INV_X1    g104(.A(G217), .ZN(new_n291));
  NOR3_X1   g105(.A1(new_n290), .A2(new_n291), .A3(G953), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n282), .A2(new_n288), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n292), .B1(new_n282), .B2(new_n288), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n254), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT95), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n282), .A2(new_n288), .ZN(new_n299));
  INV_X1    g113(.A(new_n292), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n293), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(KEYINPUT95), .A3(new_n254), .ZN(new_n303));
  INV_X1    g117(.A(G478), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(KEYINPUT15), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n298), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT96), .ZN(new_n307));
  INV_X1    g121(.A(new_n296), .ZN(new_n308));
  INV_X1    g122(.A(new_n305), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n298), .A2(new_n303), .A3(new_n307), .A4(new_n305), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(G234), .A2(G237), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(G952), .A3(new_n188), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT21), .B(G898), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n314), .A2(G902), .A3(G953), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n265), .A2(new_n313), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT97), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT97), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n265), .A2(new_n313), .A3(new_n322), .A4(new_n319), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(G214), .B1(G237), .B2(G902), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(G110), .B(G122), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT85), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT83), .B1(new_n267), .B2(G104), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT83), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n228), .A3(G107), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n267), .A2(G104), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G101), .ZN(new_n335));
  INV_X1    g149(.A(G101), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n228), .A2(G107), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n267), .A2(KEYINPUT3), .A3(G104), .ZN(new_n338));
  AOI21_X1  g152(.A(KEYINPUT3), .B1(new_n267), .B2(G104), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n336), .B(new_n337), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT84), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT84), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n335), .A2(new_n343), .A3(new_n340), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G119), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G116), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n273), .A2(G119), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT5), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n347), .A2(KEYINPUT5), .ZN(new_n352));
  INV_X1    g166(.A(G113), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT2), .B(G113), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n351), .A2(new_n354), .B1(new_n350), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n329), .B1(new_n345), .B2(new_n357), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n335), .A2(new_n343), .A3(new_n340), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n343), .B1(new_n335), .B2(new_n340), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n329), .B(new_n357), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n350), .A2(new_n356), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n349), .A2(new_n355), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n368), .B1(new_n228), .B2(G107), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n267), .A2(KEYINPUT3), .A3(G104), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n369), .A2(new_n370), .B1(new_n228), .B2(G107), .ZN(new_n371));
  NOR3_X1   g185(.A1(new_n371), .A2(KEYINPUT4), .A3(new_n336), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(new_n371), .B2(new_n336), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n375), .B1(new_n371), .B2(new_n336), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(KEYINPUT81), .A3(G101), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n374), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n374), .A2(new_n376), .A3(new_n378), .A4(KEYINPUT82), .ZN(new_n382));
  AOI211_X1 g196(.A(new_n367), .B(new_n372), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n328), .B1(new_n363), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n382), .ZN(new_n385));
  INV_X1    g199(.A(new_n372), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n366), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT85), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n361), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n387), .A2(new_n390), .A3(new_n327), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n384), .A2(KEYINPUT6), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n393), .B(new_n328), .C1(new_n363), .C2(new_n383), .ZN(new_n394));
  INV_X1    g208(.A(G146), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G143), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n190), .A2(G146), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n396), .A2(new_n397), .A3(KEYINPUT0), .A4(G128), .ZN(new_n398));
  XNOR2_X1  g212(.A(G143), .B(G146), .ZN(new_n399));
  OR2_X1    g213(.A1(KEYINPUT0), .A2(G128), .ZN(new_n400));
  NAND2_X1  g214(.A1(KEYINPUT0), .A2(G128), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n398), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT86), .B1(new_n404), .B2(new_n210), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n396), .A2(new_n397), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n396), .A2(KEYINPUT1), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n407), .A3(G128), .ZN(new_n408));
  INV_X1    g222(.A(G128), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n396), .B(new_n397), .C1(KEYINPUT1), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n210), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT86), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n403), .A2(new_n413), .A3(G125), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n405), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G224), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(G953), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n415), .B(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n392), .A2(new_n394), .A3(new_n418), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n335), .A2(new_n340), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n388), .B1(new_n420), .B2(new_n357), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n327), .B(KEYINPUT8), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT7), .B1(new_n416), .B2(G953), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n415), .A2(new_n424), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n415), .A2(KEYINPUT87), .A3(new_n424), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT87), .B1(new_n415), .B2(new_n424), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n423), .B(new_n425), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(G902), .B1(new_n429), .B2(new_n391), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n419), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(G210), .B1(G237), .B2(G902), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n419), .A2(new_n430), .A3(new_n432), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n326), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G221), .ZN(new_n437));
  INV_X1    g251(.A(new_n290), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n437), .B1(new_n438), .B2(new_n254), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT66), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n398), .B(new_n441), .C1(new_n399), .C2(new_n402), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n406), .A2(new_n401), .A3(new_n400), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n441), .B1(new_n444), .B2(new_n398), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n385), .A2(new_n446), .A3(new_n386), .ZN(new_n447));
  INV_X1    g261(.A(G137), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT64), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT64), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G137), .ZN(new_n451));
  AND2_X1   g265(.A1(KEYINPUT11), .A2(G134), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(KEYINPUT11), .A2(G134), .ZN(new_n454));
  NOR2_X1   g268(.A1(KEYINPUT11), .A2(G134), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n454), .B1(new_n455), .B2(G137), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G131), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT65), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n453), .A2(new_n194), .A3(new_n456), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n457), .A2(KEYINPUT65), .A3(G131), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n411), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n420), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT10), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(KEYINPUT10), .B(new_n464), .C1(new_n359), .C2(new_n360), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n447), .A2(new_n463), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n463), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n403), .A2(KEYINPUT66), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n386), .A2(new_n442), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n473), .B1(new_n381), .B2(new_n382), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n467), .A2(new_n468), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(G110), .B(G140), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n188), .A2(G227), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n477), .B(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n470), .A2(new_n476), .A3(new_n480), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n474), .A2(new_n475), .A3(new_n471), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n465), .B1(new_n345), .B2(new_n464), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(KEYINPUT12), .A3(new_n471), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT12), .B1(new_n483), .B2(new_n471), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n482), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g301(.A(G469), .B(new_n481), .C1(new_n487), .C2(new_n480), .ZN(new_n488));
  INV_X1    g302(.A(G469), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n489), .A2(new_n254), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n463), .B1(new_n447), .B2(new_n469), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n479), .B1(new_n493), .B2(new_n482), .ZN(new_n494));
  INV_X1    g308(.A(new_n484), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n470), .B(new_n480), .C1(new_n495), .C2(new_n485), .ZN(new_n496));
  AOI211_X1 g310(.A(G469), .B(G902), .C1(new_n494), .C2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n440), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n324), .A2(new_n436), .A3(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT26), .B(G101), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n187), .A2(new_n188), .A3(G210), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n501), .B(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n503), .B(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n449), .A2(new_n451), .A3(new_n279), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n194), .B1(G134), .B2(G137), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n460), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n411), .B1(new_n509), .B2(KEYINPUT68), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT68), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n460), .A2(new_n511), .A3(new_n508), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n461), .A2(new_n462), .A3(new_n442), .A4(new_n472), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n514), .A3(new_n367), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT28), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n514), .A2(KEYINPUT67), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT67), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n446), .A2(new_n519), .A3(new_n462), .A4(new_n461), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n518), .A2(new_n367), .A3(new_n520), .A4(new_n513), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n461), .A2(new_n462), .A3(new_n404), .ZN(new_n522));
  OR2_X1    g336(.A1(new_n509), .A2(new_n411), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n366), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT28), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n517), .B1(new_n527), .B2(KEYINPUT73), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT73), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n526), .A2(new_n529), .A3(KEYINPUT28), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n505), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT30), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(new_n510), .B2(new_n512), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n518), .A2(new_n520), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT69), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT69), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n518), .A2(new_n534), .A3(new_n520), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n524), .A2(new_n533), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n366), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT70), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n539), .A2(KEYINPUT70), .A3(new_n542), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n521), .A2(new_n505), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT72), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n548), .B(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT31), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT70), .B1(new_n539), .B2(new_n542), .ZN(new_n552));
  AOI211_X1 g366(.A(new_n544), .B(new_n541), .C1(new_n536), .C2(new_n538), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n550), .B(KEYINPUT31), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n532), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT32), .ZN(new_n557));
  NOR2_X1   g371(.A1(G472), .A2(G902), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT31), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n531), .B1(new_n562), .B2(new_n554), .ZN(new_n563));
  INV_X1    g377(.A(new_n558), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT32), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n521), .B1(new_n552), .B2(new_n553), .ZN(new_n566));
  INV_X1    g380(.A(new_n505), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n528), .A2(new_n505), .A3(new_n530), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT74), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT29), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n528), .A2(KEYINPUT74), .A3(new_n505), .A4(new_n530), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n568), .A2(new_n571), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n518), .A2(new_n520), .A3(new_n513), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n366), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(KEYINPUT75), .A3(new_n521), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT75), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n575), .A2(new_n578), .A3(new_n366), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(KEYINPUT28), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n517), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n582), .A2(new_n572), .A3(new_n567), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(G902), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n574), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n559), .A2(new_n565), .B1(G472), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT23), .ZN(new_n587));
  AOI22_X1  g401(.A1(KEYINPUT77), .A2(new_n587), .B1(new_n409), .B2(G119), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(KEYINPUT77), .B2(new_n587), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n346), .A2(G128), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n409), .A2(KEYINPUT23), .A3(G119), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT76), .ZN(new_n592));
  OR2_X1    g406(.A1(new_n591), .A2(KEYINPUT76), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n589), .A2(new_n590), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(G110), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n409), .A2(G119), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n590), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT24), .B(G110), .ZN(new_n598));
  OAI221_X1 g412(.A(new_n595), .B1(new_n597), .B2(new_n598), .C1(new_n239), .C2(new_n238), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n598), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n594), .B2(G110), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n213), .A2(new_n214), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n202), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT22), .B(G137), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n606));
  XOR2_X1   g420(.A(new_n605), .B(new_n606), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n604), .B(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n291), .B1(G234), .B2(new_n254), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(G902), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(new_n611), .B(KEYINPUT79), .Z(new_n612));
  NAND2_X1  g426(.A1(new_n608), .A2(new_n254), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT25), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT25), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n608), .A2(new_n615), .A3(new_n254), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n616), .A3(new_n609), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n500), .A2(new_n586), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(new_n336), .ZN(G3));
  NAND2_X1  g434(.A1(new_n436), .A2(new_n319), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n298), .A2(new_n303), .A3(new_n304), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n300), .B2(KEYINPUT100), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n302), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n301), .A2(new_n293), .A3(new_n624), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n626), .A2(new_n627), .A3(G478), .A4(new_n254), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n622), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n264), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n621), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n556), .A2(new_n558), .ZN(new_n632));
  INV_X1    g446(.A(new_n618), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n633), .A3(new_n499), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT99), .ZN(new_n636));
  INV_X1    g450(.A(G472), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n556), .A2(new_n254), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT98), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n556), .A2(KEYINPUT98), .A3(new_n254), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n636), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n639), .B1(new_n563), .B2(G902), .ZN(new_n643));
  AND4_X1   g457(.A1(new_n636), .A2(new_n641), .A3(new_n643), .A4(G472), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n631), .B(new_n635), .C1(new_n642), .C2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT34), .B(G104), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  NAND3_X1  g461(.A1(new_n640), .A2(new_n636), .A3(new_n641), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n641), .A2(new_n643), .A3(G472), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT99), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n621), .A2(new_n264), .A3(new_n313), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n651), .A2(new_n635), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  AND2_X1   g469(.A1(new_n321), .A2(new_n323), .ZN(new_n656));
  INV_X1    g470(.A(new_n607), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(KEYINPUT36), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n604), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n610), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n617), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n499), .A2(new_n436), .A3(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n632), .B(new_n663), .C1(new_n642), .C2(new_n644), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT37), .B(G110), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G12));
  OR2_X1    g480(.A1(new_n318), .A2(G900), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n315), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n313), .A2(new_n264), .A3(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n670), .A2(new_n499), .A3(new_n436), .A4(new_n661), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n586), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(new_n409), .ZN(G30));
  NAND2_X1  g487(.A1(new_n434), .A2(new_n435), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT38), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR4_X1   g490(.A1(new_n265), .A2(new_n661), .A3(new_n313), .A4(new_n326), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n668), .B(KEYINPUT39), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n498), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT40), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n677), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AOI211_X1 g496(.A(new_n676), .B(new_n682), .C1(new_n681), .C2(new_n680), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n559), .A2(new_n565), .ZN(new_n684));
  INV_X1    g498(.A(new_n560), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n577), .A2(new_n567), .A3(new_n579), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n254), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(G472), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G143), .ZN(G45));
  NAND3_X1  g505(.A1(new_n264), .A2(new_n629), .A3(new_n668), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n499), .A2(new_n436), .A3(new_n693), .A4(new_n661), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n586), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(new_n395), .ZN(G48));
  NAND2_X1  g510(.A1(new_n585), .A2(G472), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n557), .B1(new_n556), .B2(new_n558), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n563), .A2(KEYINPUT32), .A3(new_n564), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n494), .A2(new_n496), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n254), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(G469), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n701), .A2(new_n489), .A3(new_n254), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n440), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(KEYINPUT101), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT101), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n703), .A2(new_n707), .A3(new_n440), .A4(new_n704), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n700), .A2(new_n633), .A3(new_n631), .A4(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT41), .B(G113), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT102), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n710), .B(new_n712), .ZN(G15));
  NAND4_X1  g527(.A1(new_n700), .A2(new_n633), .A3(new_n652), .A4(new_n709), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  INV_X1    g529(.A(new_n435), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n432), .B1(new_n419), .B2(new_n430), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n661), .B(new_n325), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n705), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n700), .A2(new_n324), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G119), .ZN(G21));
  OAI21_X1  g535(.A(G472), .B1(new_n563), .B2(G902), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n582), .A2(new_n567), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n723), .B1(new_n551), .B2(new_n555), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n558), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT103), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n618), .B(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n706), .A2(new_n319), .A3(new_n708), .ZN(new_n730));
  INV_X1    g544(.A(new_n313), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n436), .A2(new_n264), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G122), .ZN(G24));
  INV_X1    g549(.A(KEYINPUT104), .ZN(new_n736));
  INV_X1    g550(.A(new_n705), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n737), .A2(new_n436), .A3(new_n693), .A4(new_n661), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n736), .B1(new_n726), .B2(new_n738), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n718), .A2(new_n692), .A3(new_n705), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n740), .A2(KEYINPUT104), .A3(new_n725), .A4(new_n722), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G125), .ZN(G27));
  NAND3_X1  g557(.A1(new_n434), .A2(new_n325), .A3(new_n435), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n498), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n700), .A2(new_n633), .A3(new_n693), .A4(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT42), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n586), .A2(new_n728), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n744), .A2(new_n498), .A3(new_n692), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n749), .A2(KEYINPUT42), .ZN(new_n750));
  AOI22_X1  g564(.A1(new_n746), .A2(new_n747), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n194), .ZN(G33));
  NAND4_X1  g566(.A1(new_n700), .A2(new_n633), .A3(new_n670), .A4(new_n745), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G134), .ZN(G36));
  OAI21_X1  g568(.A(new_n481), .B1(new_n487), .B2(new_n480), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT105), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n489), .B1(new_n755), .B2(new_n756), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n490), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n761), .A2(KEYINPUT46), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n704), .B1(new_n761), .B2(KEYINPUT46), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n440), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n764), .A2(new_n679), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n651), .A2(new_n632), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT106), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT43), .ZN(new_n768));
  XOR2_X1   g582(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n769));
  INV_X1    g583(.A(new_n629), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n770), .A2(new_n264), .ZN(new_n771));
  MUX2_X1   g585(.A(new_n768), .B(new_n769), .S(new_n771), .Z(new_n772));
  NAND3_X1  g586(.A1(new_n766), .A2(new_n661), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n744), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT107), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n765), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n773), .A2(new_n774), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT108), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n778), .B(new_n780), .C1(new_n777), .C2(new_n776), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G137), .ZN(G39));
  NOR2_X1   g596(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n783));
  NAND2_X1  g597(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n764), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n786), .B1(new_n764), .B2(new_n785), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n700), .A2(new_n633), .A3(new_n692), .A4(new_n744), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(new_n199), .ZN(G42));
  INV_X1    g605(.A(new_n728), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n792), .A2(new_n325), .A3(new_n440), .A4(new_n771), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n703), .A2(new_n704), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT49), .ZN(new_n795));
  OR4_X1    g609(.A1(new_n689), .A2(new_n793), .A3(new_n675), .A4(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n315), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n772), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n744), .A2(new_n705), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n748), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT48), .ZN(new_n802));
  INV_X1    g616(.A(G952), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n799), .A2(new_n633), .A3(new_n797), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n689), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n630), .ZN(new_n806));
  AOI211_X1 g620(.A(new_n803), .B(G953), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n798), .A2(new_n729), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n737), .A2(new_n436), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n802), .B(new_n807), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n705), .A2(new_n325), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n676), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI211_X1 g627(.A(new_n813), .B(new_n808), .C1(new_n811), .C2(new_n812), .ZN(new_n814));
  XOR2_X1   g628(.A(new_n814), .B(KEYINPUT50), .Z(new_n815));
  NAND2_X1  g629(.A1(new_n562), .A2(new_n554), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n564), .B1(new_n816), .B2(new_n723), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n817), .B1(new_n638), .B2(G472), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n800), .A2(new_n661), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n805), .A2(new_n265), .A3(new_n770), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT51), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n815), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n787), .B1(new_n440), .B2(new_n794), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n808), .A2(new_n744), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n826), .A2(KEYINPUT114), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(KEYINPUT114), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n824), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n810), .B1(new_n823), .B2(new_n829), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n829), .B(KEYINPUT115), .Z(new_n831));
  XNOR2_X1  g645(.A(new_n815), .B(KEYINPUT117), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n831), .A2(new_n821), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n830), .B1(new_n833), .B2(KEYINPUT51), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT110), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n653), .A2(new_n664), .ZN(new_n836));
  OR3_X1    g650(.A1(new_n500), .A2(new_n586), .A3(new_n618), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n645), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n835), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n634), .B1(new_n648), .B2(new_n650), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n619), .B1(new_n840), .B2(new_n631), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(KEYINPUT110), .A3(new_n653), .A4(new_n664), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n671), .ZN(new_n844));
  INV_X1    g658(.A(new_n694), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n700), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n732), .A2(new_n498), .A3(new_n661), .A4(new_n669), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n689), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n742), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT52), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT111), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n818), .A2(new_n851), .A3(new_n661), .A4(new_n749), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n722), .A2(new_n749), .A3(new_n661), .A4(new_n725), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT111), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n265), .A2(new_n661), .A3(new_n313), .A4(new_n668), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n700), .A2(new_n745), .A3(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n855), .A2(new_n753), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n742), .A2(new_n846), .A3(new_n859), .A4(new_n848), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n850), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  AND4_X1   g675(.A1(new_n710), .A2(new_n714), .A3(new_n720), .A4(new_n734), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n746), .A2(new_n747), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n748), .A2(new_n750), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n843), .A2(new_n867), .A3(KEYINPUT53), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT53), .B1(new_n843), .B2(new_n867), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT54), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n871), .A2(KEYINPUT112), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n839), .A2(new_n842), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n684), .A2(new_n697), .B1(new_n671), .B2(new_n694), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n874), .B1(new_n739), .B2(new_n741), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n859), .B1(new_n875), .B2(new_n848), .ZN(new_n876));
  INV_X1    g690(.A(new_n860), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n862), .A2(KEYINPUT113), .A3(new_n865), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT113), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n710), .A2(new_n714), .A3(new_n720), .A4(new_n734), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n880), .B1(new_n881), .B2(new_n751), .ZN(new_n882));
  AND4_X1   g696(.A1(KEYINPUT53), .A2(new_n855), .A3(new_n753), .A4(new_n857), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n878), .A2(new_n879), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n873), .A2(new_n884), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n885), .A2(new_n869), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n871), .B(KEYINPUT112), .C1(KEYINPUT54), .C2(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n872), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n834), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n803), .A2(new_n188), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT118), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n796), .B1(new_n889), .B2(new_n891), .ZN(G75));
  AND2_X1   g706(.A1(new_n886), .A2(G902), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(G210), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n392), .A2(new_n394), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(new_n418), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT55), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n894), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT119), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n188), .A2(G952), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n898), .B1(new_n894), .B2(new_n895), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(G51));
  XNOR2_X1  g717(.A(new_n886), .B(KEYINPUT54), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n490), .B(KEYINPUT57), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n701), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n893), .A2(new_n760), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n901), .B1(new_n907), .B2(new_n908), .ZN(G54));
  NAND2_X1  g723(.A1(KEYINPUT58), .A2(G475), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT120), .Z(new_n911));
  AND3_X1   g725(.A1(new_n893), .A2(new_n248), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n248), .B1(new_n893), .B2(new_n911), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n912), .A2(new_n913), .A3(new_n901), .ZN(G60));
  AND2_X1   g728(.A1(new_n626), .A2(new_n627), .ZN(new_n915));
  NAND2_X1  g729(.A1(G478), .A2(G902), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT59), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n915), .B1(new_n888), .B2(new_n917), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n904), .A2(new_n915), .A3(new_n917), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n901), .A3(new_n919), .ZN(G63));
  XNOR2_X1  g734(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n291), .A2(new_n254), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n923), .B1(new_n885), .B2(new_n869), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT122), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI211_X1 g740(.A(KEYINPUT122), .B(new_n923), .C1(new_n885), .C2(new_n869), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n659), .ZN(new_n929));
  INV_X1    g743(.A(new_n901), .ZN(new_n930));
  INV_X1    g744(.A(new_n608), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n926), .A2(new_n931), .A3(new_n927), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n929), .A2(KEYINPUT61), .A3(new_n930), .A4(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT124), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n930), .ZN(new_n935));
  AOI22_X1  g749(.A1(new_n935), .A2(KEYINPUT123), .B1(new_n659), .B2(new_n928), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT123), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n932), .A2(new_n937), .A3(new_n930), .ZN(new_n938));
  AOI211_X1 g752(.A(new_n934), .B(KEYINPUT61), .C1(new_n936), .C2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n935), .A2(KEYINPUT123), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n938), .A3(new_n929), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT124), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n933), .B1(new_n939), .B2(new_n943), .ZN(G66));
  OAI21_X1  g758(.A(G953), .B1(new_n316), .B2(new_n416), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n873), .A2(new_n881), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n945), .B1(new_n946), .B2(G953), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n896), .B1(G898), .B2(new_n188), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(G69));
  NOR4_X1   g763(.A1(new_n765), .A2(new_n586), .A3(new_n728), .A4(new_n732), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT125), .Z(new_n951));
  OAI211_X1 g765(.A(new_n753), .B(new_n875), .C1(new_n787), .C2(new_n789), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n951), .A2(new_n751), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n953), .A2(new_n781), .A3(new_n188), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n539), .A2(new_n540), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(new_n208), .Z(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(G900), .B2(G953), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n690), .A2(new_n875), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n313), .A2(new_n264), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n680), .B1(new_n806), .B2(new_n962), .ZN(new_n963));
  NOR4_X1   g777(.A1(new_n586), .A2(new_n618), .A3(new_n744), .A4(new_n963), .ZN(new_n964));
  NOR4_X1   g778(.A1(new_n790), .A2(new_n960), .A3(new_n961), .A4(new_n964), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n781), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n956), .B1(new_n966), .B2(G953), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n958), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(G72));
  NAND3_X1  g784(.A1(new_n547), .A2(new_n567), .A3(new_n521), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n953), .A2(new_n781), .A3(new_n946), .ZN(new_n972));
  NAND2_X1  g786(.A1(G472), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT63), .Z(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(KEYINPUT126), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n972), .A2(new_n977), .A3(new_n974), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n971), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n974), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n980), .B1(new_n568), .B2(new_n560), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT127), .Z(new_n982));
  AOI21_X1  g796(.A(new_n901), .B1(new_n870), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n980), .B1(new_n966), .B2(new_n946), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n566), .A2(new_n505), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n979), .A2(new_n986), .ZN(G57));
endmodule


