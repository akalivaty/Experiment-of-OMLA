

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U554 ( .A1(n547), .A2(G2104), .ZN(n888) );
  AND2_X1 U555 ( .A1(G2104), .A2(G2105), .ZN(n886) );
  BUF_X1 U556 ( .A(n552), .Z(n543) );
  NOR2_X1 U557 ( .A1(n719), .A2(n718), .ZN(n720) );
  INV_X1 U558 ( .A(KEYINPUT28), .ZN(n700) );
  NOR2_X1 U559 ( .A1(G168), .A2(n735), .ZN(n737) );
  BUF_X1 U560 ( .A(n543), .Z(n889) );
  XOR2_X1 U561 ( .A(KEYINPUT17), .B(n542), .Z(n523) );
  XOR2_X1 U562 ( .A(KEYINPUT73), .B(n592), .Z(n524) );
  XOR2_X1 U563 ( .A(KEYINPUT65), .B(n553), .Z(n525) );
  AND2_X1 U564 ( .A1(n817), .A2(n833), .ZN(n526) );
  AND2_X1 U565 ( .A1(n787), .A2(n786), .ZN(n527) );
  NOR2_X1 U566 ( .A1(n756), .A2(n757), .ZN(n733) );
  NOR2_X1 U567 ( .A1(n699), .A2(n698), .ZN(n702) );
  INV_X1 U568 ( .A(n746), .ZN(n726) );
  INV_X1 U569 ( .A(KEYINPUT98), .ZN(n736) );
  INV_X1 U570 ( .A(KEYINPUT29), .ZN(n724) );
  INV_X1 U571 ( .A(KEYINPUT99), .ZN(n744) );
  XNOR2_X1 U572 ( .A(n745), .B(n744), .ZN(n751) );
  INV_X1 U573 ( .A(KEYINPUT100), .ZN(n774) );
  NAND2_X1 U574 ( .A1(n694), .A2(n789), .ZN(n746) );
  NOR2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n542) );
  OR2_X1 U576 ( .A1(n818), .A2(n526), .ZN(n819) );
  NOR2_X2 U577 ( .A1(n667), .A2(n533), .ZN(n651) );
  NOR2_X2 U578 ( .A1(G2104), .A2(n547), .ZN(n885) );
  XNOR2_X1 U579 ( .A(n597), .B(KEYINPUT15), .ZN(n962) );
  XNOR2_X1 U580 ( .A(KEYINPUT7), .B(KEYINPUT76), .ZN(n541) );
  NOR2_X1 U581 ( .A1(G651), .A2(G543), .ZN(n656) );
  NAND2_X1 U582 ( .A1(n656), .A2(G89), .ZN(n528) );
  XNOR2_X1 U583 ( .A(n528), .B(KEYINPUT4), .ZN(n530) );
  XOR2_X1 U584 ( .A(KEYINPUT0), .B(G543), .Z(n667) );
  INV_X1 U585 ( .A(G651), .ZN(n533) );
  NAND2_X1 U586 ( .A1(G76), .A2(n651), .ZN(n529) );
  NAND2_X1 U587 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U588 ( .A(KEYINPUT5), .B(n531), .ZN(n539) );
  NOR2_X1 U589 ( .A1(G651), .A2(n667), .ZN(n662) );
  NAND2_X1 U590 ( .A1(n662), .A2(G51), .ZN(n532) );
  XOR2_X1 U591 ( .A(KEYINPUT75), .B(n532), .Z(n536) );
  NOR2_X1 U592 ( .A1(G543), .A2(n533), .ZN(n534) );
  XOR2_X1 U593 ( .A(KEYINPUT1), .B(n534), .Z(n666) );
  NAND2_X1 U594 ( .A1(n666), .A2(G63), .ZN(n535) );
  NAND2_X1 U595 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U596 ( .A(KEYINPUT6), .B(n537), .Z(n538) );
  NAND2_X1 U597 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U598 ( .A(n541), .B(n540), .ZN(G168) );
  INV_X1 U599 ( .A(G2105), .ZN(n547) );
  NAND2_X1 U600 ( .A1(n888), .A2(G102), .ZN(n545) );
  XNOR2_X1 U601 ( .A(KEYINPUT66), .B(n523), .ZN(n552) );
  NAND2_X1 U602 ( .A1(G138), .A2(n543), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U604 ( .A(KEYINPUT90), .B(n546), .ZN(n551) );
  NAND2_X1 U605 ( .A1(G126), .A2(n885), .ZN(n549) );
  NAND2_X1 U606 ( .A1(G114), .A2(n886), .ZN(n548) );
  NAND2_X1 U607 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U608 ( .A1(n551), .A2(n550), .ZN(G164) );
  AND2_X1 U609 ( .A1(n552), .A2(G137), .ZN(n556) );
  NAND2_X1 U610 ( .A1(n885), .A2(G125), .ZN(n554) );
  NAND2_X1 U611 ( .A1(G113), .A2(n886), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n525), .ZN(n555) );
  NOR2_X1 U613 ( .A1(n556), .A2(n555), .ZN(n559) );
  NAND2_X1 U614 ( .A1(G101), .A2(n888), .ZN(n557) );
  XOR2_X1 U615 ( .A(KEYINPUT23), .B(n557), .Z(n558) );
  AND2_X1 U616 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X2 U617 ( .A(KEYINPUT64), .B(n560), .ZN(G160) );
  NAND2_X1 U618 ( .A1(G64), .A2(n666), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G52), .A2(n662), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n562), .A2(n561), .ZN(n570) );
  NAND2_X1 U621 ( .A1(G77), .A2(n651), .ZN(n565) );
  NAND2_X1 U622 ( .A1(n656), .A2(G90), .ZN(n563) );
  XOR2_X1 U623 ( .A(KEYINPUT67), .B(n563), .Z(n564) );
  NAND2_X1 U624 ( .A1(n565), .A2(n564), .ZN(n568) );
  XNOR2_X1 U625 ( .A(KEYINPUT68), .B(KEYINPUT69), .ZN(n566) );
  XNOR2_X1 U626 ( .A(n566), .B(KEYINPUT9), .ZN(n567) );
  XNOR2_X1 U627 ( .A(n568), .B(n567), .ZN(n569) );
  NOR2_X1 U628 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U629 ( .A(n571), .B(KEYINPUT70), .ZN(G171) );
  INV_X1 U630 ( .A(G171), .ZN(G301) );
  NAND2_X1 U631 ( .A1(G72), .A2(n651), .ZN(n573) );
  NAND2_X1 U632 ( .A1(G85), .A2(n656), .ZN(n572) );
  NAND2_X1 U633 ( .A1(n573), .A2(n572), .ZN(n577) );
  NAND2_X1 U634 ( .A1(G60), .A2(n666), .ZN(n575) );
  NAND2_X1 U635 ( .A1(G47), .A2(n662), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n575), .A2(n574), .ZN(n576) );
  OR2_X1 U637 ( .A1(n577), .A2(n576), .ZN(G290) );
  AND2_X1 U638 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U639 ( .A(G57), .ZN(G237) );
  INV_X1 U640 ( .A(G132), .ZN(G219) );
  INV_X1 U641 ( .A(G82), .ZN(G220) );
  NAND2_X1 U642 ( .A1(G7), .A2(G661), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U644 ( .A(G223), .ZN(n839) );
  NAND2_X1 U645 ( .A1(n839), .A2(G567), .ZN(n579) );
  XOR2_X1 U646 ( .A(KEYINPUT11), .B(n579), .Z(G234) );
  NAND2_X1 U647 ( .A1(n651), .A2(G68), .ZN(n580) );
  XNOR2_X1 U648 ( .A(KEYINPUT72), .B(n580), .ZN(n583) );
  NAND2_X1 U649 ( .A1(n656), .A2(G81), .ZN(n581) );
  XNOR2_X1 U650 ( .A(KEYINPUT12), .B(n581), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U652 ( .A(n584), .B(KEYINPUT13), .ZN(n586) );
  NAND2_X1 U653 ( .A1(G43), .A2(n662), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U655 ( .A1(n666), .A2(G56), .ZN(n587) );
  XOR2_X1 U656 ( .A(KEYINPUT14), .B(n587), .Z(n588) );
  NOR2_X1 U657 ( .A1(n589), .A2(n588), .ZN(n970) );
  NAND2_X1 U658 ( .A1(n970), .A2(G860), .ZN(G153) );
  NAND2_X1 U659 ( .A1(G301), .A2(G868), .ZN(n599) );
  NAND2_X1 U660 ( .A1(G66), .A2(n666), .ZN(n591) );
  NAND2_X1 U661 ( .A1(G92), .A2(n656), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n596) );
  NAND2_X1 U663 ( .A1(n651), .A2(G79), .ZN(n592) );
  NAND2_X1 U664 ( .A1(n662), .A2(G54), .ZN(n593) );
  NAND2_X1 U665 ( .A1(n524), .A2(n593), .ZN(n594) );
  XNOR2_X1 U666 ( .A(KEYINPUT74), .B(n594), .ZN(n595) );
  NOR2_X1 U667 ( .A1(n596), .A2(n595), .ZN(n597) );
  INV_X1 U668 ( .A(G868), .ZN(n678) );
  NAND2_X1 U669 ( .A1(n962), .A2(n678), .ZN(n598) );
  NAND2_X1 U670 ( .A1(n599), .A2(n598), .ZN(G284) );
  XOR2_X1 U671 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U672 ( .A1(G65), .A2(n666), .ZN(n601) );
  NAND2_X1 U673 ( .A1(G53), .A2(n662), .ZN(n600) );
  NAND2_X1 U674 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U675 ( .A(KEYINPUT71), .B(n602), .ZN(n606) );
  NAND2_X1 U676 ( .A1(G78), .A2(n651), .ZN(n604) );
  NAND2_X1 U677 ( .A1(G91), .A2(n656), .ZN(n603) );
  AND2_X1 U678 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n606), .A2(n605), .ZN(G299) );
  XNOR2_X1 U680 ( .A(KEYINPUT77), .B(G868), .ZN(n607) );
  NOR2_X1 U681 ( .A1(G286), .A2(n607), .ZN(n610) );
  NOR2_X1 U682 ( .A1(G868), .A2(G299), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n608), .B(KEYINPUT78), .ZN(n609) );
  NOR2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U685 ( .A(KEYINPUT79), .B(n611), .Z(G297) );
  INV_X1 U686 ( .A(G860), .ZN(n612) );
  NAND2_X1 U687 ( .A1(n612), .A2(G559), .ZN(n613) );
  INV_X1 U688 ( .A(n962), .ZN(n635) );
  NAND2_X1 U689 ( .A1(n613), .A2(n635), .ZN(n614) );
  XNOR2_X1 U690 ( .A(n614), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U691 ( .A1(n635), .A2(G868), .ZN(n615) );
  NOR2_X1 U692 ( .A1(G559), .A2(n615), .ZN(n617) );
  INV_X1 U693 ( .A(n970), .ZN(n638) );
  NOR2_X1 U694 ( .A1(G868), .A2(n638), .ZN(n616) );
  NOR2_X1 U695 ( .A1(n617), .A2(n616), .ZN(G282) );
  NAND2_X1 U696 ( .A1(G123), .A2(n885), .ZN(n618) );
  XNOR2_X1 U697 ( .A(n618), .B(KEYINPUT18), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n888), .A2(G99), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n886), .A2(G111), .ZN(n622) );
  NAND2_X1 U701 ( .A1(G135), .A2(n889), .ZN(n621) );
  NAND2_X1 U702 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U703 ( .A1(n624), .A2(n623), .ZN(n1017) );
  XNOR2_X1 U704 ( .A(G2096), .B(n1017), .ZN(n626) );
  INV_X1 U705 ( .A(G2100), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(G156) );
  NAND2_X1 U707 ( .A1(G93), .A2(n656), .ZN(n627) );
  XNOR2_X1 U708 ( .A(n627), .B(KEYINPUT82), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G67), .A2(n666), .ZN(n629) );
  NAND2_X1 U710 ( .A1(G80), .A2(n651), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U712 ( .A1(G55), .A2(n662), .ZN(n630) );
  XNOR2_X1 U713 ( .A(KEYINPUT83), .B(n630), .ZN(n631) );
  NOR2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U715 ( .A1(n634), .A2(n633), .ZN(n677) );
  NAND2_X1 U716 ( .A1(G559), .A2(n635), .ZN(n636) );
  XNOR2_X1 U717 ( .A(n636), .B(KEYINPUT80), .ZN(n637) );
  XNOR2_X1 U718 ( .A(n638), .B(n637), .ZN(n675) );
  NOR2_X1 U719 ( .A1(G860), .A2(n675), .ZN(n639) );
  XNOR2_X1 U720 ( .A(n639), .B(KEYINPUT81), .ZN(n640) );
  XNOR2_X1 U721 ( .A(n677), .B(n640), .ZN(G145) );
  NAND2_X1 U722 ( .A1(G88), .A2(n656), .ZN(n641) );
  XNOR2_X1 U723 ( .A(n641), .B(KEYINPUT88), .ZN(n648) );
  NAND2_X1 U724 ( .A1(G62), .A2(n666), .ZN(n643) );
  NAND2_X1 U725 ( .A1(G75), .A2(n651), .ZN(n642) );
  NAND2_X1 U726 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U727 ( .A1(G50), .A2(n662), .ZN(n644) );
  XNOR2_X1 U728 ( .A(KEYINPUT87), .B(n644), .ZN(n645) );
  NOR2_X1 U729 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U731 ( .A(KEYINPUT89), .B(n649), .Z(G303) );
  INV_X1 U732 ( .A(G303), .ZN(G166) );
  NAND2_X1 U733 ( .A1(G61), .A2(n666), .ZN(n650) );
  XNOR2_X1 U734 ( .A(n650), .B(KEYINPUT84), .ZN(n661) );
  NAND2_X1 U735 ( .A1(G73), .A2(n651), .ZN(n652) );
  XNOR2_X1 U736 ( .A(n652), .B(KEYINPUT86), .ZN(n653) );
  XNOR2_X1 U737 ( .A(n653), .B(KEYINPUT2), .ZN(n655) );
  NAND2_X1 U738 ( .A1(G48), .A2(n662), .ZN(n654) );
  NAND2_X1 U739 ( .A1(n655), .A2(n654), .ZN(n659) );
  NAND2_X1 U740 ( .A1(G86), .A2(n656), .ZN(n657) );
  XNOR2_X1 U741 ( .A(KEYINPUT85), .B(n657), .ZN(n658) );
  NOR2_X1 U742 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U743 ( .A1(n661), .A2(n660), .ZN(G305) );
  NAND2_X1 U744 ( .A1(G49), .A2(n662), .ZN(n664) );
  NAND2_X1 U745 ( .A1(G74), .A2(G651), .ZN(n663) );
  NAND2_X1 U746 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U747 ( .A1(n666), .A2(n665), .ZN(n669) );
  NAND2_X1 U748 ( .A1(n667), .A2(G87), .ZN(n668) );
  NAND2_X1 U749 ( .A1(n669), .A2(n668), .ZN(G288) );
  INV_X1 U750 ( .A(G299), .ZN(n967) );
  XNOR2_X1 U751 ( .A(n967), .B(G166), .ZN(n674) );
  XNOR2_X1 U752 ( .A(KEYINPUT19), .B(G305), .ZN(n670) );
  XNOR2_X1 U753 ( .A(n670), .B(G288), .ZN(n671) );
  XNOR2_X1 U754 ( .A(n671), .B(G290), .ZN(n672) );
  XNOR2_X1 U755 ( .A(n672), .B(n677), .ZN(n673) );
  XNOR2_X1 U756 ( .A(n674), .B(n673), .ZN(n913) );
  XOR2_X1 U757 ( .A(n675), .B(n913), .Z(n676) );
  NAND2_X1 U758 ( .A1(n676), .A2(G868), .ZN(n680) );
  NAND2_X1 U759 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U760 ( .A1(n680), .A2(n679), .ZN(G295) );
  NAND2_X1 U761 ( .A1(G2078), .A2(G2084), .ZN(n681) );
  XOR2_X1 U762 ( .A(KEYINPUT20), .B(n681), .Z(n682) );
  NAND2_X1 U763 ( .A1(G2090), .A2(n682), .ZN(n683) );
  XNOR2_X1 U764 ( .A(KEYINPUT21), .B(n683), .ZN(n684) );
  NAND2_X1 U765 ( .A1(n684), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U766 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U767 ( .A1(G220), .A2(G219), .ZN(n685) );
  XOR2_X1 U768 ( .A(KEYINPUT22), .B(n685), .Z(n686) );
  NOR2_X1 U769 ( .A1(G218), .A2(n686), .ZN(n687) );
  NAND2_X1 U770 ( .A1(G96), .A2(n687), .ZN(n845) );
  NAND2_X1 U771 ( .A1(n845), .A2(G2106), .ZN(n691) );
  NAND2_X1 U772 ( .A1(G69), .A2(G120), .ZN(n688) );
  NOR2_X1 U773 ( .A1(G237), .A2(n688), .ZN(n689) );
  NAND2_X1 U774 ( .A1(G108), .A2(n689), .ZN(n846) );
  NAND2_X1 U775 ( .A1(n846), .A2(G567), .ZN(n690) );
  NAND2_X1 U776 ( .A1(n691), .A2(n690), .ZN(n869) );
  NAND2_X1 U777 ( .A1(G661), .A2(G483), .ZN(n692) );
  NOR2_X1 U778 ( .A1(n869), .A2(n692), .ZN(n842) );
  NAND2_X1 U779 ( .A1(n842), .A2(G36), .ZN(G176) );
  INV_X1 U780 ( .A(KEYINPUT96), .ZN(n693) );
  NAND2_X1 U781 ( .A1(G40), .A2(G160), .ZN(n788) );
  XNOR2_X1 U782 ( .A(n693), .B(n788), .ZN(n694) );
  NOR2_X1 U783 ( .A1(G164), .A2(G1384), .ZN(n789) );
  NAND2_X1 U784 ( .A1(G8), .A2(n746), .ZN(n784) );
  NOR2_X1 U785 ( .A1(G1981), .A2(G305), .ZN(n695) );
  XOR2_X1 U786 ( .A(n695), .B(KEYINPUT24), .Z(n696) );
  NOR2_X1 U787 ( .A1(n784), .A2(n696), .ZN(n778) );
  XNOR2_X1 U788 ( .A(G1981), .B(G305), .ZN(n979) );
  NAND2_X1 U789 ( .A1(n726), .A2(G2072), .ZN(n697) );
  XNOR2_X1 U790 ( .A(n697), .B(KEYINPUT27), .ZN(n699) );
  INV_X1 U791 ( .A(G1956), .ZN(n996) );
  NOR2_X1 U792 ( .A1(n996), .A2(n726), .ZN(n698) );
  NOR2_X1 U793 ( .A1(n702), .A2(n967), .ZN(n701) );
  XNOR2_X1 U794 ( .A(n701), .B(n700), .ZN(n723) );
  NAND2_X1 U795 ( .A1(n702), .A2(n967), .ZN(n721) );
  INV_X1 U796 ( .A(G1341), .ZN(n995) );
  NAND2_X1 U797 ( .A1(G1348), .A2(n962), .ZN(n973) );
  NAND2_X1 U798 ( .A1(n995), .A2(n973), .ZN(n703) );
  NAND2_X1 U799 ( .A1(n746), .A2(n703), .ZN(n706) );
  NAND2_X1 U800 ( .A1(n726), .A2(G1996), .ZN(n704) );
  XNOR2_X1 U801 ( .A(KEYINPUT26), .B(KEYINPUT97), .ZN(n707) );
  NAND2_X1 U802 ( .A1(n704), .A2(n707), .ZN(n705) );
  NAND2_X1 U803 ( .A1(n706), .A2(n705), .ZN(n714) );
  NAND2_X1 U804 ( .A1(n962), .A2(G2067), .ZN(n710) );
  INV_X1 U805 ( .A(n707), .ZN(n708) );
  NAND2_X1 U806 ( .A1(G1996), .A2(n708), .ZN(n709) );
  NAND2_X1 U807 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U808 ( .A1(n711), .A2(n726), .ZN(n712) );
  NAND2_X1 U809 ( .A1(n970), .A2(n712), .ZN(n713) );
  NOR2_X1 U810 ( .A1(n714), .A2(n713), .ZN(n719) );
  NAND2_X1 U811 ( .A1(G1348), .A2(n746), .ZN(n716) );
  NAND2_X1 U812 ( .A1(G2067), .A2(n726), .ZN(n715) );
  NAND2_X1 U813 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U814 ( .A1(n717), .A2(n962), .ZN(n718) );
  NAND2_X1 U815 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U816 ( .A1(n723), .A2(n722), .ZN(n725) );
  XNOR2_X1 U817 ( .A(n725), .B(n724), .ZN(n730) );
  XOR2_X1 U818 ( .A(G2078), .B(KEYINPUT25), .Z(n945) );
  NOR2_X1 U819 ( .A1(n945), .A2(n746), .ZN(n728) );
  NOR2_X1 U820 ( .A1(n726), .A2(G1961), .ZN(n727) );
  NOR2_X1 U821 ( .A1(n728), .A2(n727), .ZN(n738) );
  OR2_X1 U822 ( .A1(n738), .A2(G301), .ZN(n729) );
  NAND2_X1 U823 ( .A1(n730), .A2(n729), .ZN(n743) );
  INV_X1 U824 ( .A(G8), .ZN(n731) );
  NOR2_X1 U825 ( .A1(n731), .A2(G1966), .ZN(n732) );
  AND2_X1 U826 ( .A1(n746), .A2(n732), .ZN(n756) );
  NOR2_X1 U827 ( .A1(G2084), .A2(n746), .ZN(n757) );
  NAND2_X1 U828 ( .A1(G8), .A2(n733), .ZN(n734) );
  XNOR2_X1 U829 ( .A(KEYINPUT30), .B(n734), .ZN(n735) );
  XNOR2_X1 U830 ( .A(n737), .B(n736), .ZN(n740) );
  NAND2_X1 U831 ( .A1(G301), .A2(n738), .ZN(n739) );
  NAND2_X1 U832 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U833 ( .A(KEYINPUT31), .B(n741), .ZN(n742) );
  NAND2_X1 U834 ( .A1(n743), .A2(n742), .ZN(n754) );
  NAND2_X1 U835 ( .A1(n754), .A2(G286), .ZN(n745) );
  NOR2_X1 U836 ( .A1(G1971), .A2(n784), .ZN(n748) );
  NOR2_X1 U837 ( .A1(G2090), .A2(n746), .ZN(n747) );
  NOR2_X1 U838 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U839 ( .A1(G303), .A2(n749), .ZN(n750) );
  NAND2_X1 U840 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U841 ( .A1(n752), .A2(G8), .ZN(n753) );
  XNOR2_X1 U842 ( .A(KEYINPUT32), .B(n753), .ZN(n780) );
  INV_X1 U843 ( .A(n754), .ZN(n755) );
  NOR2_X1 U844 ( .A1(n756), .A2(n755), .ZN(n759) );
  NAND2_X1 U845 ( .A1(G8), .A2(n757), .ZN(n758) );
  NAND2_X1 U846 ( .A1(n759), .A2(n758), .ZN(n779) );
  NAND2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n763) );
  AND2_X1 U848 ( .A1(n779), .A2(n763), .ZN(n761) );
  INV_X1 U849 ( .A(KEYINPUT33), .ZN(n760) );
  AND2_X1 U850 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U851 ( .A1(n780), .A2(n762), .ZN(n773) );
  INV_X1 U852 ( .A(n763), .ZN(n959) );
  NOR2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n768) );
  NOR2_X1 U854 ( .A1(G1971), .A2(G303), .ZN(n764) );
  NOR2_X1 U855 ( .A1(n768), .A2(n764), .ZN(n968) );
  OR2_X1 U856 ( .A1(n959), .A2(n968), .ZN(n765) );
  OR2_X1 U857 ( .A1(KEYINPUT33), .A2(n765), .ZN(n766) );
  OR2_X1 U858 ( .A1(n784), .A2(n766), .ZN(n771) );
  INV_X1 U859 ( .A(n784), .ZN(n767) );
  NAND2_X1 U860 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U861 ( .A1(n769), .A2(KEYINPUT33), .ZN(n770) );
  AND2_X1 U862 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n775) );
  XNOR2_X1 U864 ( .A(n775), .B(n774), .ZN(n776) );
  NOR2_X1 U865 ( .A1(n979), .A2(n776), .ZN(n777) );
  NOR2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n787) );
  NAND2_X1 U867 ( .A1(n779), .A2(n780), .ZN(n783) );
  NOR2_X1 U868 ( .A1(G2090), .A2(G303), .ZN(n781) );
  NAND2_X1 U869 ( .A1(G8), .A2(n781), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n785) );
  NAND2_X1 U871 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U872 ( .A1(n789), .A2(n788), .ZN(n833) );
  XNOR2_X1 U873 ( .A(G2067), .B(KEYINPUT37), .ZN(n831) );
  NAND2_X1 U874 ( .A1(G140), .A2(n889), .ZN(n790) );
  XOR2_X1 U875 ( .A(KEYINPUT91), .B(n790), .Z(n792) );
  NAND2_X1 U876 ( .A1(n888), .A2(G104), .ZN(n791) );
  NAND2_X1 U877 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U878 ( .A(KEYINPUT34), .B(n793), .ZN(n799) );
  NAND2_X1 U879 ( .A1(G128), .A2(n885), .ZN(n795) );
  NAND2_X1 U880 ( .A1(G116), .A2(n886), .ZN(n794) );
  NAND2_X1 U881 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U882 ( .A(KEYINPUT92), .B(n796), .Z(n797) );
  XNOR2_X1 U883 ( .A(KEYINPUT35), .B(n797), .ZN(n798) );
  NOR2_X1 U884 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U885 ( .A(KEYINPUT36), .B(n800), .ZN(n910) );
  NOR2_X1 U886 ( .A1(n831), .A2(n910), .ZN(n1040) );
  NAND2_X1 U887 ( .A1(n833), .A2(n1040), .ZN(n801) );
  XOR2_X1 U888 ( .A(KEYINPUT93), .B(n801), .Z(n828) );
  INV_X1 U889 ( .A(n828), .ZN(n818) );
  NAND2_X1 U890 ( .A1(G105), .A2(n888), .ZN(n802) );
  XNOR2_X1 U891 ( .A(n802), .B(KEYINPUT38), .ZN(n809) );
  NAND2_X1 U892 ( .A1(G129), .A2(n885), .ZN(n804) );
  NAND2_X1 U893 ( .A1(G117), .A2(n886), .ZN(n803) );
  NAND2_X1 U894 ( .A1(n804), .A2(n803), .ZN(n807) );
  NAND2_X1 U895 ( .A1(G141), .A2(n889), .ZN(n805) );
  XNOR2_X1 U896 ( .A(KEYINPUT95), .B(n805), .ZN(n806) );
  NOR2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U898 ( .A1(n809), .A2(n808), .ZN(n907) );
  AND2_X1 U899 ( .A1(n907), .A2(G1996), .ZN(n1020) );
  NAND2_X1 U900 ( .A1(G119), .A2(n885), .ZN(n811) );
  NAND2_X1 U901 ( .A1(G107), .A2(n886), .ZN(n810) );
  NAND2_X1 U902 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U903 ( .A(KEYINPUT94), .B(n812), .ZN(n816) );
  NAND2_X1 U904 ( .A1(n888), .A2(G95), .ZN(n814) );
  NAND2_X1 U905 ( .A1(G131), .A2(n889), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n900) );
  INV_X1 U908 ( .A(G1991), .ZN(n823) );
  NOR2_X1 U909 ( .A1(n900), .A2(n823), .ZN(n1018) );
  OR2_X1 U910 ( .A1(n1020), .A2(n1018), .ZN(n817) );
  NOR2_X1 U911 ( .A1(n527), .A2(n819), .ZN(n821) );
  XNOR2_X1 U912 ( .A(G1986), .B(G290), .ZN(n958) );
  NAND2_X1 U913 ( .A1(n958), .A2(n833), .ZN(n820) );
  NAND2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n836) );
  NOR2_X1 U915 ( .A1(G1996), .A2(n907), .ZN(n822) );
  XOR2_X1 U916 ( .A(KEYINPUT101), .B(n822), .Z(n1024) );
  AND2_X1 U917 ( .A1(n823), .A2(n900), .ZN(n1019) );
  NOR2_X1 U918 ( .A1(G1986), .A2(G290), .ZN(n824) );
  NOR2_X1 U919 ( .A1(n1019), .A2(n824), .ZN(n825) );
  NOR2_X1 U920 ( .A1(n526), .A2(n825), .ZN(n826) );
  NOR2_X1 U921 ( .A1(n1024), .A2(n826), .ZN(n827) );
  XNOR2_X1 U922 ( .A(n827), .B(KEYINPUT39), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U924 ( .A(n830), .B(KEYINPUT102), .ZN(n832) );
  NAND2_X1 U925 ( .A1(n831), .A2(n910), .ZN(n1037) );
  NAND2_X1 U926 ( .A1(n832), .A2(n1037), .ZN(n834) );
  NAND2_X1 U927 ( .A1(n834), .A2(n833), .ZN(n835) );
  NAND2_X1 U928 ( .A1(n836), .A2(n835), .ZN(n838) );
  XOR2_X1 U929 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n837) );
  XNOR2_X1 U930 ( .A(n838), .B(n837), .ZN(G329) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n839), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n840) );
  NAND2_X1 U933 ( .A1(G661), .A2(n840), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n841) );
  XNOR2_X1 U935 ( .A(KEYINPUT106), .B(n841), .ZN(n843) );
  NAND2_X1 U936 ( .A1(n843), .A2(n842), .ZN(n844) );
  XOR2_X1 U937 ( .A(KEYINPUT107), .B(n844), .Z(G188) );
  INV_X1 U939 ( .A(G120), .ZN(G236) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  INV_X1 U941 ( .A(G69), .ZN(G235) );
  NOR2_X1 U942 ( .A1(n846), .A2(n845), .ZN(G325) );
  INV_X1 U943 ( .A(G325), .ZN(G261) );
  XOR2_X1 U944 ( .A(G2096), .B(G2678), .Z(n848) );
  XNOR2_X1 U945 ( .A(G2090), .B(KEYINPUT43), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U947 ( .A(n849), .B(KEYINPUT42), .Z(n851) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2072), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U950 ( .A(KEYINPUT108), .B(G2100), .Z(n853) );
  XNOR2_X1 U951 ( .A(G2078), .B(G2084), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(G227) );
  XOR2_X1 U954 ( .A(KEYINPUT109), .B(KEYINPUT112), .Z(n857) );
  XNOR2_X1 U955 ( .A(KEYINPUT41), .B(KEYINPUT111), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U957 ( .A(n858), .B(KEYINPUT110), .Z(n860) );
  XNOR2_X1 U958 ( .A(G1996), .B(G1991), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n868) );
  XOR2_X1 U960 ( .A(G1976), .B(G1971), .Z(n862) );
  XNOR2_X1 U961 ( .A(G1986), .B(G1961), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U963 ( .A(G2474), .B(G1981), .Z(n864) );
  XNOR2_X1 U964 ( .A(G1966), .B(G1956), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U966 ( .A(n866), .B(n865), .Z(n867) );
  XNOR2_X1 U967 ( .A(n868), .B(n867), .ZN(G229) );
  INV_X1 U968 ( .A(n869), .ZN(G319) );
  NAND2_X1 U969 ( .A1(G124), .A2(n885), .ZN(n870) );
  XNOR2_X1 U970 ( .A(n870), .B(KEYINPUT44), .ZN(n872) );
  NAND2_X1 U971 ( .A1(n888), .A2(G100), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n876) );
  NAND2_X1 U973 ( .A1(n886), .A2(G112), .ZN(n874) );
  NAND2_X1 U974 ( .A1(G136), .A2(n889), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U976 ( .A1(n876), .A2(n875), .ZN(G162) );
  NAND2_X1 U977 ( .A1(n888), .A2(G103), .ZN(n878) );
  NAND2_X1 U978 ( .A1(G139), .A2(n889), .ZN(n877) );
  NAND2_X1 U979 ( .A1(n878), .A2(n877), .ZN(n883) );
  NAND2_X1 U980 ( .A1(G127), .A2(n885), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G115), .A2(n886), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U983 ( .A(KEYINPUT47), .B(n881), .Z(n882) );
  NOR2_X1 U984 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U985 ( .A(KEYINPUT115), .B(n884), .Z(n1031) );
  NAND2_X1 U986 ( .A1(G130), .A2(n885), .ZN(n897) );
  NAND2_X1 U987 ( .A1(n886), .A2(G118), .ZN(n887) );
  XNOR2_X1 U988 ( .A(KEYINPUT113), .B(n887), .ZN(n895) );
  NAND2_X1 U989 ( .A1(n888), .A2(G106), .ZN(n891) );
  NAND2_X1 U990 ( .A1(G142), .A2(n889), .ZN(n890) );
  NAND2_X1 U991 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U992 ( .A(KEYINPUT45), .B(n892), .Z(n893) );
  XNOR2_X1 U993 ( .A(KEYINPUT114), .B(n893), .ZN(n894) );
  NOR2_X1 U994 ( .A1(n895), .A2(n894), .ZN(n896) );
  NAND2_X1 U995 ( .A1(n897), .A2(n896), .ZN(n898) );
  XNOR2_X1 U996 ( .A(n898), .B(G162), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n1031), .B(n899), .ZN(n902) );
  XNOR2_X1 U998 ( .A(G160), .B(n900), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n906) );
  XOR2_X1 U1000 ( .A(KEYINPUT48), .B(KEYINPUT116), .Z(n904) );
  XNOR2_X1 U1001 ( .A(n1017), .B(KEYINPUT46), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1003 ( .A(n906), .B(n905), .Z(n909) );
  XOR2_X1 U1004 ( .A(G164), .B(n907), .Z(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n911) );
  XOR2_X1 U1006 ( .A(n911), .B(n910), .Z(n912) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n912), .ZN(G395) );
  XNOR2_X1 U1008 ( .A(n913), .B(n962), .ZN(n914) );
  XNOR2_X1 U1009 ( .A(n914), .B(G286), .ZN(n916) );
  XOR2_X1 U1010 ( .A(n970), .B(G301), .Z(n915) );
  XNOR2_X1 U1011 ( .A(n916), .B(n915), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n917), .ZN(G397) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n919) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(KEYINPUT118), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(n919), .B(n918), .ZN(n920) );
  XOR2_X1 U1016 ( .A(KEYINPUT117), .B(n920), .Z(n933) );
  XNOR2_X1 U1017 ( .A(G2451), .B(G2427), .ZN(n930) );
  XOR2_X1 U1018 ( .A(KEYINPUT105), .B(G2443), .Z(n922) );
  XNOR2_X1 U1019 ( .A(G2435), .B(G2438), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(n922), .B(n921), .ZN(n926) );
  XOR2_X1 U1021 ( .A(G2454), .B(G2430), .Z(n924) );
  XNOR2_X1 U1022 ( .A(G1348), .B(G1341), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(n924), .B(n923), .ZN(n925) );
  XOR2_X1 U1024 ( .A(n926), .B(n925), .Z(n928) );
  XNOR2_X1 U1025 ( .A(G2446), .B(KEYINPUT104), .ZN(n927) );
  XNOR2_X1 U1026 ( .A(n928), .B(n927), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(n930), .B(n929), .ZN(n931) );
  NAND2_X1 U1028 ( .A1(n931), .A2(G14), .ZN(n936) );
  NAND2_X1 U1029 ( .A1(G319), .A2(n936), .ZN(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(G395), .A2(G397), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(G225) );
  INV_X1 U1033 ( .A(G225), .ZN(G308) );
  INV_X1 U1034 ( .A(G108), .ZN(G238) );
  INV_X1 U1035 ( .A(n936), .ZN(G401) );
  XOR2_X1 U1036 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n1048) );
  INV_X1 U1037 ( .A(KEYINPUT55), .ZN(n1042) );
  XNOR2_X1 U1038 ( .A(G2090), .B(G35), .ZN(n950) );
  XNOR2_X1 U1039 ( .A(G1991), .B(G25), .ZN(n938) );
  XNOR2_X1 U1040 ( .A(G33), .B(G2072), .ZN(n937) );
  NOR2_X1 U1041 ( .A1(n938), .A2(n937), .ZN(n944) );
  XOR2_X1 U1042 ( .A(G32), .B(G1996), .Z(n939) );
  NAND2_X1 U1043 ( .A1(n939), .A2(G28), .ZN(n942) );
  XNOR2_X1 U1044 ( .A(KEYINPUT120), .B(G2067), .ZN(n940) );
  XNOR2_X1 U1045 ( .A(G26), .B(n940), .ZN(n941) );
  NOR2_X1 U1046 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1047 ( .A1(n944), .A2(n943), .ZN(n947) );
  XNOR2_X1 U1048 ( .A(G27), .B(n945), .ZN(n946) );
  NOR2_X1 U1049 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1050 ( .A(KEYINPUT53), .B(n948), .ZN(n949) );
  NOR2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n953) );
  XOR2_X1 U1052 ( .A(G2084), .B(KEYINPUT54), .Z(n951) );
  XNOR2_X1 U1053 ( .A(G34), .B(n951), .ZN(n952) );
  NAND2_X1 U1054 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1055 ( .A(n1042), .B(n954), .ZN(n956) );
  INV_X1 U1056 ( .A(G29), .ZN(n955) );
  NAND2_X1 U1057 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1058 ( .A1(G11), .A2(n957), .ZN(n1016) );
  XNOR2_X1 U1059 ( .A(G16), .B(KEYINPUT56), .ZN(n984) );
  NOR2_X1 U1060 ( .A1(n959), .A2(n958), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(G171), .B(G1961), .ZN(n961) );
  NAND2_X1 U1062 ( .A1(G1971), .A2(G303), .ZN(n960) );
  NAND2_X1 U1063 ( .A1(n961), .A2(n960), .ZN(n964) );
  NOR2_X1 U1064 ( .A1(G1348), .A2(n962), .ZN(n963) );
  NOR2_X1 U1065 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1066 ( .A1(n966), .A2(n965), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(n967), .B(G1956), .ZN(n969) );
  NAND2_X1 U1068 ( .A1(n969), .A2(n968), .ZN(n972) );
  XOR2_X1 U1069 ( .A(n970), .B(G1341), .Z(n971) );
  NOR2_X1 U1070 ( .A1(n972), .A2(n971), .ZN(n974) );
  NAND2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(G1966), .B(KEYINPUT121), .ZN(n977) );
  XNOR2_X1 U1074 ( .A(n977), .B(G168), .ZN(n978) );
  NOR2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1076 ( .A(KEYINPUT57), .B(n980), .Z(n981) );
  NAND2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n1014) );
  INV_X1 U1079 ( .A(G16), .ZN(n1012) );
  XNOR2_X1 U1080 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n1010) );
  XNOR2_X1 U1081 ( .A(G1971), .B(G22), .ZN(n986) );
  XNOR2_X1 U1082 ( .A(G23), .B(G1976), .ZN(n985) );
  NOR2_X1 U1083 ( .A1(n986), .A2(n985), .ZN(n988) );
  XOR2_X1 U1084 ( .A(G1986), .B(G24), .Z(n987) );
  NAND2_X1 U1085 ( .A1(n988), .A2(n987), .ZN(n990) );
  XOR2_X1 U1086 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n989) );
  XNOR2_X1 U1087 ( .A(n990), .B(n989), .ZN(n1008) );
  XOR2_X1 U1088 ( .A(G1981), .B(G6), .Z(n994) );
  XNOR2_X1 U1089 ( .A(KEYINPUT59), .B(KEYINPUT122), .ZN(n991) );
  XNOR2_X1 U1090 ( .A(n991), .B(G4), .ZN(n992) );
  XNOR2_X1 U1091 ( .A(G1348), .B(n992), .ZN(n993) );
  NAND2_X1 U1092 ( .A1(n994), .A2(n993), .ZN(n1000) );
  XNOR2_X1 U1093 ( .A(n995), .B(G19), .ZN(n998) );
  XNOR2_X1 U1094 ( .A(n996), .B(G20), .ZN(n997) );
  NAND2_X1 U1095 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1096 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1097 ( .A(KEYINPUT60), .B(n1001), .ZN(n1005) );
  XNOR2_X1 U1098 ( .A(G1966), .B(G21), .ZN(n1003) );
  XNOR2_X1 U1099 ( .A(G1961), .B(G5), .ZN(n1002) );
  NOR2_X1 U1100 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1101 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1102 ( .A(KEYINPUT123), .B(n1006), .ZN(n1007) );
  NAND2_X1 U1103 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1104 ( .A(n1010), .B(n1009), .ZN(n1011) );
  NAND2_X1 U1105 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1106 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1107 ( .A1(n1016), .A2(n1015), .ZN(n1046) );
  NOR2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1030) );
  XNOR2_X1 U1109 ( .A(G2084), .B(G160), .ZN(n1022) );
  NOR2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1028) );
  XOR2_X1 U1112 ( .A(G2090), .B(G162), .Z(n1023) );
  NOR2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1114 ( .A(KEYINPUT119), .B(n1025), .Z(n1026) );
  XNOR2_X1 U1115 ( .A(n1026), .B(KEYINPUT51), .ZN(n1027) );
  NOR2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1036) );
  XOR2_X1 U1118 ( .A(G2072), .B(n1031), .Z(n1033) );
  XOR2_X1 U1119 ( .A(G164), .B(G2078), .Z(n1032) );
  NOR2_X1 U1120 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XOR2_X1 U1121 ( .A(KEYINPUT50), .B(n1034), .Z(n1035) );
  NOR2_X1 U1122 ( .A1(n1036), .A2(n1035), .ZN(n1038) );
  NAND2_X1 U1123 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NOR2_X1 U1124 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XNOR2_X1 U1125 ( .A(KEYINPUT52), .B(n1041), .ZN(n1043) );
  NAND2_X1 U1126 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  NAND2_X1 U1127 ( .A1(n1044), .A2(G29), .ZN(n1045) );
  NAND2_X1 U1128 ( .A1(n1046), .A2(n1045), .ZN(n1047) );
  XOR2_X1 U1129 ( .A(n1048), .B(n1047), .Z(G150) );
  INV_X1 U1130 ( .A(G150), .ZN(G311) );
endmodule

