//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT66), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT67), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT68), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  AND2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(G125), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n464), .A2(new_n469), .ZN(G160));
  OAI21_X1  g045(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G112), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n471), .B1(new_n472), .B2(G2105), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n460), .A2(new_n461), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(new_n459), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT69), .ZN(new_n477));
  OR2_X1    g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(G2105), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI211_X1 g055(.A(new_n473), .B(new_n477), .C1(G136), .C2(new_n480), .ZN(G162));
  INV_X1    g056(.A(G138), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n483), .B1(new_n460), .B2(new_n461), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT72), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n483), .B(KEYINPUT72), .C1(new_n461), .C2(new_n460), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n486), .A2(KEYINPUT4), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n484), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n474), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n492), .A2(G126), .A3(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT70), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n459), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT70), .B(G114), .ZN(new_n503));
  NOR3_X1   g078(.A1(new_n503), .A2(KEYINPUT71), .A3(new_n459), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n493), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n491), .A2(new_n505), .ZN(G164));
  NAND2_X1  g081(.A1(G75), .A2(G543), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n507), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n510), .A2(new_n520), .A3(G88), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n519), .A2(new_n521), .A3(KEYINPUT73), .ZN(new_n522));
  AOI21_X1  g097(.A(KEYINPUT73), .B1(new_n519), .B2(new_n521), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n514), .B1(new_n522), .B2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND2_X1  g100(.A1(new_n520), .A2(G89), .ZN(new_n526));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n511), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n520), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G51), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n528), .A2(new_n533), .ZN(G168));
  AOI22_X1  g109(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G651), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n510), .A2(new_n520), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n538), .A2(new_n539), .B1(new_n531), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n537), .A2(new_n541), .ZN(G171));
  AOI22_X1  g117(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n536), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT74), .B(G43), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n538), .A2(new_n545), .B1(new_n531), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  XNOR2_X1  g129(.A(KEYINPUT76), .B(G65), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n511), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n538), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n556), .A2(G651), .B1(new_n557), .B2(G91), .ZN(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT9), .B1(new_n531), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n518), .A2(new_n561), .A3(G53), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(KEYINPUT75), .B1(new_n560), .B2(new_n562), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n558), .B1(new_n565), .B2(new_n566), .ZN(G299));
  OR2_X1    g142(.A1(new_n537), .A2(new_n541), .ZN(G301));
  INV_X1    g143(.A(G168), .ZN(G286));
  NAND2_X1  g144(.A1(new_n557), .A2(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n518), .A2(G49), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n508), .B2(new_n509), .ZN(new_n575));
  AND2_X1   g150(.A1(G73), .A2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n510), .A2(new_n520), .A3(G86), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n518), .A2(G48), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G305));
  NAND2_X1  g155(.A1(new_n557), .A2(G85), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  XNOR2_X1  g157(.A(KEYINPUT77), .B(G47), .ZN(new_n583));
  OAI221_X1 g158(.A(new_n581), .B1(new_n536), .B2(new_n582), .C1(new_n531), .C2(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  AND3_X1   g160(.A1(new_n510), .A2(new_n520), .A3(G92), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT10), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n511), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(G54), .B2(new_n518), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n585), .B1(new_n593), .B2(G868), .ZN(G284));
  OAI21_X1  g169(.A(new_n585), .B1(new_n593), .B2(G868), .ZN(G321));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  INV_X1    g171(.A(G299), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G297));
  OAI21_X1  g173(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n593), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n593), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n492), .A2(new_n467), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT13), .ZN(new_n608));
  INV_X1    g183(.A(G2100), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n475), .A2(G123), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n480), .A2(G135), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n459), .A2(G111), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n612), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G2096), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n610), .A2(new_n611), .A3(new_n618), .ZN(G156));
  INV_X1    g194(.A(KEYINPUT14), .ZN(new_n620));
  XNOR2_X1  g195(.A(G2427), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2430), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n623), .B2(new_n622), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2451), .B(G2454), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT16), .ZN(new_n627));
  XNOR2_X1  g202(.A(G1341), .B(G1348), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n625), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  AND3_X1   g208(.A1(new_n632), .A2(G14), .A3(new_n633), .ZN(G401));
  INV_X1    g209(.A(KEYINPUT18), .ZN(new_n635));
  XOR2_X1   g210(.A(G2084), .B(G2090), .Z(new_n636));
  XNOR2_X1  g211(.A(G2067), .B(G2678), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(KEYINPUT17), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n636), .A2(new_n637), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n635), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(new_n609), .ZN(new_n642));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n638), .B2(KEYINPUT18), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(new_n617), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(new_n645), .ZN(G227));
  XNOR2_X1  g221(.A(G1961), .B(G1966), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT78), .ZN(new_n648));
  XOR2_X1   g223(.A(G1956), .B(G2474), .Z(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1971), .B(G1976), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT19), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n648), .A2(new_n649), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n650), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n652), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT20), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n653), .A2(KEYINPUT20), .A3(new_n652), .ZN(new_n658));
  OAI221_X1 g233(.A(new_n654), .B1(new_n652), .B2(new_n650), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G1991), .B(G1996), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1981), .B(G1986), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n661), .A2(new_n663), .ZN(new_n666));
  AND3_X1   g241(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n665), .B1(new_n664), .B2(new_n666), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(G229));
  INV_X1    g244(.A(G29), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(G32), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n475), .A2(G129), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n467), .A2(G105), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(G141), .B2(new_n480), .ZN(new_n675));
  NAND3_X1  g250(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT91), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT26), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n671), .B1(new_n680), .B2(new_n670), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT92), .Z(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT27), .B(G1996), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(G160), .A2(G29), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT90), .B(KEYINPUT24), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G34), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n686), .B1(G29), .B2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G2084), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  NOR2_X1   g267(.A1(G168), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(new_n692), .B2(G21), .ZN(new_n694));
  INV_X1    g269(.A(G1966), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n691), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n695), .B2(new_n694), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n692), .A2(G5), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G171), .B2(new_n692), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G1961), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT30), .B(G28), .ZN(new_n701));
  OR2_X1    g276(.A1(KEYINPUT31), .A2(G11), .ZN(new_n702));
  NAND2_X1  g277(.A1(KEYINPUT31), .A2(G11), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n701), .A2(new_n670), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI221_X1 g279(.A(new_n704), .B1(new_n670), .B2(new_n616), .C1(new_n689), .C2(new_n690), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n684), .A2(new_n685), .A3(new_n697), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n670), .A2(G35), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT95), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G162), .B2(new_n670), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT29), .B(G2090), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT82), .B(G16), .Z(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n714), .A2(G19), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n548), .B2(new_n714), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT86), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1341), .ZN(new_n718));
  INV_X1    g293(.A(G2072), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n670), .A2(G33), .ZN(new_n720));
  NAND2_X1  g295(.A1(G115), .A2(G2104), .ZN(new_n721));
  INV_X1    g296(.A(G127), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n474), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT88), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n459), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(new_n724), .B2(new_n723), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT25), .ZN(new_n727));
  NAND2_X1  g302(.A1(G103), .A2(G2104), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(G2105), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n459), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n480), .A2(G139), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n720), .B1(new_n732), .B2(G29), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n712), .B(new_n718), .C1(new_n719), .C2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n713), .A2(G20), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT96), .B(KEYINPUT23), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n597), .B2(new_n692), .ZN(new_n738));
  INV_X1    g313(.A(G1956), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n733), .A2(new_n719), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT89), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n692), .A2(G4), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n593), .B2(new_n692), .ZN(new_n745));
  INV_X1    g320(.A(G1348), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n670), .A2(G26), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT28), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n480), .A2(G140), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n753));
  INV_X1    g328(.A(G116), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(G2105), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n475), .B2(G128), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n749), .B1(new_n757), .B2(G29), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2067), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n670), .A2(G27), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT93), .Z(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G164), .B2(new_n670), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT94), .B(G2078), .Z(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n747), .A2(new_n759), .A3(new_n764), .ZN(new_n765));
  NOR4_X1   g340(.A1(new_n707), .A2(new_n734), .A3(new_n743), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT97), .ZN(new_n767));
  NAND2_X1  g342(.A1(G166), .A2(new_n714), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G22), .B2(new_n714), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(KEYINPUT84), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(KEYINPUT84), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G1971), .ZN(new_n773));
  INV_X1    g348(.A(G1971), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n770), .A2(new_n774), .A3(new_n771), .ZN(new_n775));
  MUX2_X1   g350(.A(G6), .B(G305), .S(G16), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT83), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT32), .B(G1981), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n692), .A2(G23), .ZN(new_n780));
  INV_X1    g355(.A(G288), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(new_n692), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT33), .B(G1976), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n773), .A2(new_n775), .A3(new_n779), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(KEYINPUT34), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT85), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n785), .A2(KEYINPUT34), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n475), .A2(G119), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n480), .A2(G131), .ZN(new_n791));
  OR2_X1    g366(.A1(G95), .A2(G2105), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n792), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n790), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT79), .ZN(new_n795));
  MUX2_X1   g370(.A(G25), .B(new_n795), .S(G29), .Z(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT35), .B(G1991), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT80), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n796), .B(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT81), .ZN(new_n800));
  MUX2_X1   g375(.A(G24), .B(G290), .S(new_n714), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1986), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n789), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n788), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(KEYINPUT36), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT36), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n788), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n767), .B1(new_n805), .B2(new_n807), .ZN(G311));
  XOR2_X1   g383(.A(new_n766), .B(KEYINPUT97), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n805), .A2(new_n807), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(G150));
  NAND2_X1  g386(.A1(new_n593), .A2(G559), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT38), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(new_n536), .ZN(new_n815));
  INV_X1    g390(.A(G93), .ZN(new_n816));
  INV_X1    g391(.A(G55), .ZN(new_n817));
  OAI22_X1  g392(.A1(new_n538), .A2(new_n816), .B1(new_n531), .B2(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n544), .B2(new_n547), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n815), .A2(new_n818), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n548), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n813), .B(new_n823), .Z(new_n824));
  AND2_X1   g399(.A1(new_n824), .A2(KEYINPUT39), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(KEYINPUT39), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n825), .A2(new_n826), .A3(G860), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n819), .A2(G860), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT98), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT37), .Z(new_n830));
  OR2_X1    g405(.A1(new_n827), .A2(new_n830), .ZN(G145));
  NAND2_X1  g406(.A1(new_n475), .A2(G130), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n480), .A2(G142), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n459), .A2(G118), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n832), .B(new_n833), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n607), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n794), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n837), .A2(new_n838), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n840), .A2(KEYINPUT101), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n757), .B(G164), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n846), .A2(new_n679), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n732), .A2(KEYINPUT100), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n679), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n848), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n732), .A2(KEYINPUT100), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n847), .B2(new_n849), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n842), .B(new_n845), .C1(new_n850), .C2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n854), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n857));
  INV_X1    g432(.A(new_n843), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(G160), .B(KEYINPUT99), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n616), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(G162), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n855), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT102), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n855), .A2(new_n859), .A3(new_n865), .A4(new_n862), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n845), .A2(new_n842), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n868), .A2(new_n856), .A3(new_n857), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n862), .B1(new_n869), .B2(new_n855), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n870), .A2(G37), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n593), .B2(G299), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n593), .A2(G299), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n563), .B(new_n564), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n877), .A2(new_n592), .A3(KEYINPUT103), .A4(new_n558), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT41), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n597), .A2(new_n592), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n880), .B1(new_n593), .B2(G299), .ZN(new_n882));
  AOI22_X1  g457(.A1(new_n879), .A2(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n876), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n602), .B(new_n823), .ZN(new_n886));
  MUX2_X1   g461(.A(new_n883), .B(new_n885), .S(new_n886), .Z(new_n887));
  XNOR2_X1  g462(.A(G290), .B(G303), .ZN(new_n888));
  XNOR2_X1  g463(.A(G288), .B(G305), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT42), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n887), .B(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(G868), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(G868), .B2(new_n821), .ZN(G295));
  OAI21_X1  g469(.A(new_n893), .B1(G868), .B2(new_n821), .ZN(G331));
  NAND2_X1  g470(.A1(G301), .A2(KEYINPUT105), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n897));
  NAND2_X1  g472(.A1(G171), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n896), .A2(G168), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(G168), .B1(new_n896), .B2(new_n898), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n823), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OR3_X1    g478(.A1(new_n899), .A2(new_n900), .A3(new_n823), .ZN(new_n904));
  OAI211_X1 g479(.A(KEYINPUT106), .B(new_n823), .C1(new_n899), .C2(new_n900), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n884), .A4(new_n905), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n904), .A2(new_n901), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n906), .B(new_n890), .C1(new_n907), .C2(new_n883), .ZN(new_n908));
  AOI21_X1  g483(.A(G37), .B1(new_n908), .B2(KEYINPUT107), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n907), .A2(new_n883), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT107), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n910), .A2(new_n911), .A3(new_n890), .A4(new_n906), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n906), .B1(new_n907), .B2(new_n883), .ZN(new_n913));
  INV_X1    g488(.A(new_n890), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n909), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  XOR2_X1   g491(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n875), .A2(new_n882), .A3(new_n878), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(new_n885), .B2(KEYINPUT41), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n904), .A2(new_n884), .A3(new_n901), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n914), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n909), .A2(new_n912), .A3(new_n917), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n919), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n927), .A2(KEYINPUT44), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n909), .A2(new_n912), .A3(new_n925), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(new_n916), .B2(new_n918), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n928), .B1(KEYINPUT44), .B2(new_n931), .ZN(G397));
  INV_X1    g507(.A(KEYINPUT126), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n757), .B(G2067), .ZN(new_n934));
  INV_X1    g509(.A(G1384), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(new_n491), .B2(new_n505), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT45), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n465), .A2(new_n468), .ZN(new_n939));
  INV_X1    g514(.A(G125), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n478), .B2(new_n479), .ZN(new_n941));
  INV_X1    g516(.A(new_n463), .ZN(new_n942));
  OAI21_X1  g517(.A(G2105), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n939), .A2(new_n943), .A3(G40), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(G160), .A2(KEYINPUT108), .A3(G40), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n938), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n934), .A2(new_n949), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n950), .A2(KEYINPUT109), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(KEYINPUT109), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n679), .B(G1996), .ZN(new_n953));
  AOI22_X1  g528(.A1(new_n951), .A2(new_n952), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n794), .B(new_n798), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n949), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n949), .ZN(new_n957));
  XOR2_X1   g532(.A(G290), .B(G1986), .Z(new_n958));
  OAI211_X1 g533(.A(new_n954), .B(new_n956), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n959), .B(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n962));
  INV_X1    g537(.A(G8), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n500), .B1(new_n503), .B2(new_n459), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n496), .A2(G114), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n494), .A2(KEYINPUT70), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n499), .B(G2105), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(G2104), .A3(new_n967), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n488), .A2(new_n968), .A3(new_n493), .A4(new_n490), .ZN(new_n969));
  XOR2_X1   g544(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n970));
  AND3_X1   g545(.A1(new_n969), .A2(new_n935), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n972), .B1(new_n969), .B2(new_n935), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n971), .A2(new_n973), .A3(new_n948), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n946), .A2(new_n947), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n969), .A2(KEYINPUT45), .A3(new_n935), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n938), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  AOI22_X1  g552(.A1(new_n974), .A2(new_n690), .B1(new_n977), .B2(new_n695), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n963), .B1(new_n978), .B2(G168), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n695), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n936), .A2(KEYINPUT50), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n969), .A2(new_n935), .A3(new_n970), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n981), .A2(new_n975), .A3(new_n690), .A4(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(G286), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n962), .B1(new_n979), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n980), .A2(G168), .A3(new_n983), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(G8), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(KEYINPUT51), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT62), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n978), .A2(G168), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT51), .B1(new_n991), .B2(new_n988), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT62), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n979), .A2(new_n962), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n969), .A2(KEYINPUT45), .A3(new_n935), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT45), .B1(new_n969), .B2(new_n935), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n996), .A2(new_n997), .A3(new_n948), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n981), .A2(new_n975), .A3(new_n982), .ZN(new_n999));
  OAI22_X1  g574(.A1(new_n998), .A2(G1971), .B1(new_n999), .B2(G2090), .ZN(new_n1000));
  NOR2_X1   g575(.A1(G166), .A2(new_n963), .ZN(new_n1001));
  OR2_X1    g576(.A1(KEYINPUT112), .A2(KEYINPUT55), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(KEYINPUT112), .B(KEYINPUT55), .Z(new_n1004));
  OAI21_X1  g579(.A(new_n1003), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1000), .A2(new_n1005), .A3(G8), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n946), .A2(new_n969), .A3(new_n947), .A4(new_n935), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(G8), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n1009));
  INV_X1    g584(.A(G1981), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n577), .A2(new_n1010), .A3(new_n578), .A4(new_n579), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT115), .ZN(new_n1012));
  NAND2_X1  g587(.A1(G305), .A2(G1981), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1008), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1012), .A2(KEYINPUT49), .A3(new_n1013), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n781), .A2(G1976), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1007), .A2(G8), .A3(new_n1017), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n1015), .A2(new_n1016), .B1(KEYINPUT52), .B2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT113), .B(G1976), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(G288), .B2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1007), .A2(new_n1017), .A3(G8), .A4(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1022), .B(KEYINPUT114), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1006), .A2(new_n1019), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n1025));
  INV_X1    g600(.A(G2078), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n938), .A2(new_n975), .A3(new_n1026), .A4(new_n976), .ZN(new_n1027));
  INV_X1    g602(.A(G1961), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n1025), .A2(new_n1027), .B1(new_n999), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1025), .A2(G2078), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n998), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(G171), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n972), .B(new_n935), .C1(new_n491), .C2(new_n505), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n970), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n936), .A2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n969), .A2(KEYINPUT117), .A3(new_n972), .A4(new_n935), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1036), .A2(new_n1038), .A3(new_n975), .A4(new_n1039), .ZN(new_n1040));
  OAI22_X1  g615(.A1(new_n1040), .A2(G2090), .B1(new_n998), .B2(G1971), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1005), .B1(new_n1041), .B2(G8), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1024), .A2(new_n1033), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n990), .A2(new_n995), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n1045));
  INV_X1    g620(.A(G2090), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n974), .A2(new_n1046), .B1(new_n977), .B2(new_n774), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1045), .B1(new_n1047), .B2(new_n963), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1005), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1000), .A2(KEYINPUT118), .A3(G8), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n984), .A2(G8), .A3(G168), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT63), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1051), .A2(new_n1052), .A3(new_n1055), .A4(new_n1006), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1024), .A2(new_n1042), .A3(new_n1053), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1056), .B1(new_n1057), .B2(KEYINPUT63), .ZN(new_n1058));
  XOR2_X1   g633(.A(new_n1008), .B(KEYINPUT116), .Z(new_n1059));
  NAND2_X1  g634(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1060));
  INV_X1    g635(.A(G1976), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n781), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1059), .B1(new_n1062), .B2(new_n1012), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1006), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1063), .B1(new_n1052), .B2(new_n1064), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1044), .A2(new_n1058), .A3(new_n1065), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n488), .A2(new_n490), .ZN(new_n1067));
  OAI21_X1  g642(.A(G2105), .B1(new_n965), .B2(new_n966), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n466), .B1(new_n1068), .B2(new_n500), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1069), .A2(new_n967), .B1(G126), .B2(new_n475), .ZN(new_n1070));
  AOI21_X1  g645(.A(G1384), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n975), .A2(new_n1071), .A3(KEYINPUT120), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1007), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(G2067), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n999), .A2(new_n746), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n592), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1040), .A2(new_n739), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n996), .A2(new_n997), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n1082));
  XNOR2_X1  g657(.A(KEYINPUT56), .B(G2072), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1081), .A2(new_n1082), .A3(new_n975), .A4(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n938), .A2(new_n975), .A3(new_n976), .A4(new_n1083), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT119), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1080), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n558), .A2(new_n1088), .A3(new_n563), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1089), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  AOI211_X1 g667(.A(KEYINPUT121), .B(new_n1089), .C1(G299), .C2(KEYINPUT57), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1087), .A2(KEYINPUT122), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT122), .B1(new_n1087), .B2(new_n1094), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1079), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1085), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1098), .A2(new_n1082), .B1(new_n1040), .B2(new_n739), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(new_n1086), .A3(new_n1090), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT61), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1090), .B1(new_n1099), .B2(new_n1086), .ZN(new_n1103));
  AND4_X1   g678(.A1(new_n1086), .A2(new_n1080), .A3(new_n1084), .A4(new_n1090), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1077), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n592), .A2(KEYINPUT60), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1106), .A2(new_n1075), .A3(new_n1107), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT58), .B(G1341), .Z(new_n1109));
  NAND3_X1  g684(.A1(new_n1072), .A2(new_n1074), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1996), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n938), .A2(new_n975), .A3(new_n1111), .A4(new_n976), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n548), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT59), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(new_n1116), .A3(new_n548), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1108), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1106), .A2(new_n1075), .A3(new_n593), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT60), .B1(new_n1078), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1105), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1100), .A2(KEYINPUT61), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1096), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1087), .A2(new_n1094), .A3(KEYINPUT122), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1101), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1081), .A2(G40), .A3(G160), .A4(new_n1030), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1029), .A2(new_n1128), .A3(G301), .A4(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1029), .A2(G301), .A3(new_n1129), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT123), .ZN(new_n1132));
  AOI21_X1  g707(.A(G301), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1127), .B(new_n1130), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n992), .A2(new_n994), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1029), .A2(new_n1129), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(G171), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1137), .B(KEYINPUT54), .C1(G171), .C2(new_n1032), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1024), .A2(new_n1042), .ZN(new_n1139));
  AND4_X1   g714(.A1(new_n1134), .A2(new_n1135), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1126), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n961), .B1(new_n1066), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n757), .A2(G2067), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n795), .A2(new_n798), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1143), .B1(new_n954), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n957), .B1(new_n1145), .B2(KEYINPUT124), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(KEYINPUT124), .B2(new_n1145), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n949), .A2(new_n1111), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT46), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n949), .B1(new_n934), .B2(new_n679), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT47), .ZN(new_n1152));
  NOR2_X1   g727(.A1(G290), .A2(G1986), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n949), .A2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT125), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT48), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1156), .A2(new_n954), .A3(new_n956), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1147), .A2(new_n1152), .A3(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n933), .B1(new_n1142), .B2(new_n1158), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1147), .A2(new_n1152), .A3(new_n1157), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1134), .A2(new_n1135), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1161));
  OAI211_X1 g736(.A(KEYINPUT61), .B(new_n1100), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1162), .A2(new_n1105), .A3(new_n1120), .A4(new_n1118), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1161), .B1(new_n1163), .B2(new_n1101), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1044), .A2(new_n1058), .A3(new_n1065), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g741(.A(KEYINPUT126), .B(new_n1160), .C1(new_n1166), .C2(new_n961), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1159), .A2(new_n1167), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g743(.A(G319), .ZN(new_n1170));
  NOR3_X1   g744(.A1(G401), .A2(new_n1170), .A3(G227), .ZN(new_n1171));
  OAI21_X1  g745(.A(new_n1171), .B1(new_n667), .B2(new_n668), .ZN(new_n1172));
  AOI21_X1  g746(.A(new_n1172), .B1(new_n867), .B2(new_n871), .ZN(new_n1173));
  AND3_X1   g747(.A1(new_n927), .A2(new_n1173), .A3(KEYINPUT127), .ZN(new_n1174));
  AOI21_X1  g748(.A(KEYINPUT127), .B1(new_n927), .B2(new_n1173), .ZN(new_n1175));
  NOR2_X1   g749(.A1(new_n1174), .A2(new_n1175), .ZN(G308));
  NAND2_X1  g750(.A1(new_n927), .A2(new_n1173), .ZN(G225));
endmodule


