//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n451, new_n452, new_n454, new_n455,
    new_n456, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G234));
  INV_X1    g025(.A(G2106), .ZN(new_n451));
  NOR2_X1   g026(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR4_X1   g030(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  OAI22_X1  g033(.A1(new_n455), .A2(new_n451), .B1(new_n448), .B2(new_n456), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n466), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  OR2_X1    g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT69), .B1(new_n461), .B2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(new_n462), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n461), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G137), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n463), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n469), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NAND3_X1  g054(.A1(new_n471), .A2(G2105), .A3(new_n472), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n474), .A2(G136), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n468), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n482), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT70), .ZN(G162));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR4_X1   g063(.A1(new_n465), .A2(KEYINPUT4), .A3(new_n488), .A4(G2105), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n471), .A2(G138), .A3(new_n468), .A4(new_n472), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT72), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n490), .A2(KEYINPUT72), .A3(KEYINPUT4), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n489), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n471), .A2(G126), .A3(G2105), .A4(new_n472), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G114), .C2(new_n468), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n496), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n497), .A2(new_n496), .A3(new_n499), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n495), .A2(new_n503), .ZN(G164));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT5), .B1(new_n505), .B2(KEYINPUT73), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(new_n508), .A3(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n510), .A2(G62), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n516), .A2(new_n520), .ZN(G166));
  INV_X1    g096(.A(new_n514), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G51), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n528), .B2(new_n512), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  AND2_X1   g105(.A1(new_n510), .A2(new_n511), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n531), .A2(G90), .B1(new_n522), .B2(G52), .ZN(new_n532));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n506), .A2(new_n509), .ZN(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g113(.A(G651), .B1(new_n536), .B2(new_n537), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n532), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(KEYINPUT75), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(KEYINPUT75), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(G171));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n512), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n510), .A2(G56), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n517), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI211_X1 g123(.A(new_n545), .B(new_n548), .C1(G43), .C2(new_n522), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT76), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n552), .A2(new_n555), .ZN(G188));
  XNOR2_X1  g131(.A(KEYINPUT77), .B(KEYINPUT9), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n522), .A2(G53), .A3(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OAI211_X1 g135(.A(KEYINPUT77), .B(new_n559), .C1(new_n514), .C2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(G91), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n558), .B(new_n561), .C1(new_n562), .C2(new_n512), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n510), .A2(G65), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n517), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  INV_X1    g144(.A(G166), .ZN(G303));
  OAI21_X1  g145(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT78), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n531), .A2(G87), .B1(new_n522), .B2(G49), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n572), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  INV_X1    g151(.A(G86), .ZN(new_n577));
  INV_X1    g152(.A(G48), .ZN(new_n578));
  OAI22_X1  g153(.A1(new_n512), .A2(new_n577), .B1(new_n514), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n510), .A2(G61), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n517), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G305));
  INV_X1    g159(.A(G85), .ZN(new_n585));
  INV_X1    g160(.A(G47), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n512), .A2(new_n585), .B1(new_n514), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n510), .A2(G60), .ZN(new_n588));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n517), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(new_n531), .A2(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n534), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(new_n522), .B2(G54), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G171), .B2(new_n601), .ZN(G284));
  OAI21_X1  g178(.A(new_n602), .B1(G171), .B2(new_n601), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n567), .ZN(G297));
  OAI21_X1  g181(.A(new_n605), .B1(G868), .B2(new_n567), .ZN(G280));
  AND2_X1   g182(.A1(new_n595), .A2(new_n599), .ZN(new_n608));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n550), .ZN(new_n613));
  MUX2_X1   g188(.A(new_n612), .B(new_n613), .S(KEYINPUT79), .Z(G323));
  XOR2_X1   g189(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n615));
  XNOR2_X1  g190(.A(G323), .B(new_n615), .ZN(G282));
  NAND2_X1  g191(.A1(new_n474), .A2(G135), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n468), .A2(G111), .ZN(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(G123), .B2(new_n481), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT81), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2096), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n466), .A2(new_n476), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2100), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n623), .A2(new_n627), .ZN(G156));
  INV_X1    g203(.A(KEYINPUT14), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2435), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n632), .B2(new_n631), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT16), .B(G1341), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(G14), .B1(new_n634), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(new_n634), .B2(new_n640), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT82), .Z(G401));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT83), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT18), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n647), .B(KEYINPUT84), .Z(new_n651));
  NOR2_X1   g226(.A1(new_n651), .A2(new_n646), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(new_n644), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n646), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n644), .B(KEYINPUT17), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n653), .B(new_n654), .C1(new_n652), .C2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2096), .B(G2100), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  AND2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n667), .A2(KEYINPUT20), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(KEYINPUT20), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n664), .A2(new_n665), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  OR3_X1    g246(.A1(new_n663), .A2(new_n666), .A3(new_n670), .ZN(new_n672));
  NAND4_X1  g247(.A1(new_n668), .A2(new_n669), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1981), .B(G1986), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT86), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n673), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1991), .B(G1996), .Z(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n676), .B(new_n679), .ZN(G229));
  NOR2_X1   g255(.A1(G16), .A2(G23), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT87), .ZN(new_n682));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(G288), .B2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT33), .B(G1976), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(G22), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G166), .B2(new_n683), .ZN(new_n688));
  INV_X1    g263(.A(G1971), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n683), .A2(G6), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(new_n583), .B2(new_n683), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT32), .B(G1981), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n686), .A2(new_n690), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT34), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n481), .A2(G119), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n474), .A2(G131), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n468), .A2(G107), .ZN(new_n699));
  OAI21_X1  g274(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n697), .B(new_n698), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G25), .B(new_n701), .S(G29), .Z(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT35), .B(G1991), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n683), .A2(G24), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n591), .B2(new_n683), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1986), .ZN(new_n707));
  OR3_X1    g282(.A1(new_n696), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(KEYINPUT36), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(KEYINPUT88), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(KEYINPUT88), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n710), .A2(KEYINPUT36), .A3(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT89), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n709), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n713), .B2(new_n712), .ZN(new_n715));
  NOR2_X1   g290(.A1(G16), .A2(G19), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n550), .B2(G16), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(G1341), .Z(new_n718));
  NOR2_X1   g293(.A1(G286), .A2(new_n683), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT97), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G16), .B2(G21), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G1966), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT98), .B(KEYINPUT23), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n683), .A2(G20), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n567), .B2(new_n683), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1956), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT31), .B(G11), .ZN(new_n729));
  INV_X1    g304(.A(G28), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(KEYINPUT30), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT30), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(G28), .ZN(new_n734));
  AND2_X1   g309(.A1(KEYINPUT24), .A2(G34), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n732), .B1(KEYINPUT24), .B2(G34), .ZN(new_n736));
  OAI22_X1  g311(.A1(G160), .A2(new_n732), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI221_X1 g312(.A(new_n729), .B1(new_n731), .B2(new_n734), .C1(new_n737), .C2(G2084), .ZN(new_n738));
  AOI211_X1 g313(.A(new_n728), .B(new_n738), .C1(G2084), .C2(new_n737), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n683), .A2(G4), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n608), .B2(new_n683), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT90), .B(G1348), .Z(new_n742));
  AOI22_X1  g317(.A1(new_n622), .A2(G29), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n739), .B(new_n743), .C1(new_n741), .C2(new_n742), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n732), .A2(G33), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n476), .A2(G103), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT25), .Z(new_n747));
  INV_X1    g322(.A(G139), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(new_n473), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT92), .Z(new_n750));
  AOI22_X1  g325(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT93), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n468), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n752), .B2(new_n751), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n745), .B1(new_n755), .B2(G29), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2072), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n474), .A2(G141), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT94), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n481), .A2(G129), .ZN(new_n761));
  NAND3_X1  g336(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT26), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n764), .A2(new_n765), .B1(G105), .B2(new_n476), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n761), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n760), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT95), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n770), .A2(new_n732), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n732), .B2(G32), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT27), .B(G1996), .Z(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n757), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n723), .A2(new_n744), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G29), .A2(G35), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G162), .B2(G29), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT29), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n779), .A2(G2090), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n779), .A2(G2090), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n732), .A2(G27), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G164), .B2(new_n732), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G2078), .ZN(new_n784));
  NOR2_X1   g359(.A1(G5), .A2(G16), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G171), .B2(G16), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1961), .ZN(new_n787));
  NOR4_X1   g362(.A1(new_n780), .A2(new_n781), .A3(new_n784), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n772), .A2(new_n774), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT96), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n732), .A2(G26), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n481), .A2(G128), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n474), .A2(G140), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n468), .A2(G116), .ZN(new_n794));
  OAI21_X1  g369(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n792), .B(new_n793), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT91), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n791), .B1(new_n797), .B2(G29), .ZN(new_n798));
  MUX2_X1   g373(.A(new_n791), .B(new_n798), .S(KEYINPUT28), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G2067), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n776), .A2(new_n788), .A3(new_n790), .A4(new_n800), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT99), .Z(new_n802));
  AND2_X1   g377(.A1(new_n715), .A2(new_n802), .ZN(G311));
  NAND2_X1  g378(.A1(new_n715), .A2(new_n802), .ZN(G150));
  INV_X1    g379(.A(G93), .ZN(new_n805));
  INV_X1    g380(.A(G55), .ZN(new_n806));
  OAI22_X1  g381(.A1(new_n512), .A2(new_n805), .B1(new_n514), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n510), .A2(G67), .ZN(new_n808));
  NAND2_X1  g383(.A1(G80), .A2(G543), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n517), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G860), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT37), .ZN(new_n814));
  INV_X1    g389(.A(new_n811), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n549), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n550), .B2(new_n815), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT39), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n600), .A2(new_n609), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(new_n812), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n818), .A2(new_n820), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n814), .B1(new_n822), .B2(new_n823), .ZN(G145));
  XNOR2_X1  g399(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n768), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n755), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n770), .B(KEYINPUT102), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n829), .B2(new_n755), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n497), .A2(new_n499), .ZN(new_n831));
  INV_X1    g406(.A(new_n489), .ZN(new_n832));
  AND3_X1   g407(.A1(new_n490), .A2(KEYINPUT72), .A3(KEYINPUT4), .ZN(new_n833));
  AOI21_X1  g408(.A(KEYINPUT72), .B1(new_n490), .B2(KEYINPUT4), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT101), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n831), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n495), .A2(KEYINPUT101), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n797), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n830), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n474), .A2(G142), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n468), .A2(G118), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(G130), .B2(new_n481), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n625), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(new_n701), .Z(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n828), .B(new_n840), .C1(new_n829), .C2(new_n755), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n842), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT103), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n850), .B1(new_n842), .B2(new_n851), .ZN(new_n854));
  XNOR2_X1  g429(.A(G162), .B(KEYINPUT100), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n478), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n622), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n853), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G37), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n857), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n854), .B(KEYINPUT104), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n862), .B1(new_n863), .B2(new_n853), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n826), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n853), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(new_n857), .ZN(new_n867));
  AOI21_X1  g442(.A(G37), .B1(new_n853), .B2(new_n858), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n868), .A3(new_n825), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n865), .A2(new_n869), .ZN(G395));
  NAND2_X1  g445(.A1(new_n608), .A2(G299), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n600), .A2(new_n567), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT106), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT107), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n817), .B(new_n611), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n873), .A2(KEYINPUT41), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(new_n877), .B2(KEYINPUT41), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n883), .A2(new_n880), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(G166), .B(new_n583), .Z(new_n886));
  XNOR2_X1  g461(.A(G288), .B(new_n591), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT108), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(new_n889), .B2(KEYINPUT42), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(KEYINPUT42), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n890), .B(new_n891), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n885), .B(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n893), .A2(new_n601), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n811), .A2(G868), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n894), .A2(new_n895), .ZN(G295));
  OAI21_X1  g471(.A(KEYINPUT109), .B1(new_n894), .B2(new_n895), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT109), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n815), .A2(new_n601), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n898), .B(new_n899), .C1(new_n893), .C2(new_n601), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(G331));
  XNOR2_X1  g476(.A(G171), .B(G286), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n817), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n903), .A2(new_n874), .A3(new_n876), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(new_n883), .B2(new_n903), .ZN(new_n905));
  AOI21_X1  g480(.A(G37), .B1(new_n905), .B2(new_n888), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n888), .B1(new_n879), .B2(new_n903), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT41), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT110), .B1(new_n877), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n873), .A2(new_n908), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n873), .A2(KEYINPUT110), .A3(new_n908), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n903), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n907), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n906), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n905), .A2(new_n888), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT43), .B1(new_n918), .B2(new_n906), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT44), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n915), .A2(KEYINPUT43), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n916), .B1(new_n918), .B2(new_n906), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n920), .B1(new_n923), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g499(.A(KEYINPUT112), .ZN(new_n925));
  INV_X1    g500(.A(G1384), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n839), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n928));
  INV_X1    g503(.A(G40), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n478), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n931), .A2(KEYINPUT111), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT111), .ZN(new_n933));
  AOI21_X1  g508(.A(G1384), .B1(new_n837), .B2(new_n838), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n934), .A2(KEYINPUT45), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n933), .B1(new_n935), .B2(new_n930), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n925), .B1(new_n932), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n931), .A2(KEYINPUT111), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n935), .A2(new_n933), .A3(new_n930), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(KEYINPUT112), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n941), .A2(G1996), .A3(new_n768), .ZN(new_n942));
  INV_X1    g517(.A(G2067), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n797), .B(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n938), .A2(new_n939), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G1996), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n949), .A3(new_n770), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n942), .A2(new_n946), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n701), .A2(new_n703), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n701), .A2(new_n703), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n941), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n591), .B(G1986), .Z(new_n956));
  AOI21_X1  g531(.A(new_n955), .B1(new_n948), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G8), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n497), .A2(new_n496), .A3(new_n499), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(new_n500), .ZN(new_n960));
  AOI21_X1  g535(.A(G1384), .B1(new_n835), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT45), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n930), .B(new_n962), .C1(new_n934), .C2(KEYINPUT45), .ZN(new_n963));
  INV_X1    g538(.A(G1966), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n930), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n926), .B1(new_n495), .B2(new_n503), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT50), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n966), .B1(new_n968), .B2(KEYINPUT114), .ZN(new_n969));
  INV_X1    g544(.A(G2084), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n839), .A2(new_n971), .A3(new_n926), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT114), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n967), .A2(new_n973), .A3(KEYINPUT50), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n969), .A2(new_n970), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n958), .B1(new_n965), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT120), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT51), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT114), .B1(new_n961), .B2(new_n971), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n979), .A2(new_n974), .A3(new_n930), .ZN(new_n980));
  AOI211_X1 g555(.A(KEYINPUT50), .B(G1384), .C1(new_n837), .C2(new_n838), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n982), .A2(new_n970), .B1(new_n964), .B2(new_n963), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n958), .B1(new_n983), .B2(G168), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n978), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n965), .A2(new_n975), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(G8), .ZN(new_n987));
  NOR2_X1   g562(.A1(G168), .A2(new_n958), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n987), .A2(new_n977), .A3(KEYINPUT51), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n986), .A2(new_n988), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n985), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT62), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT124), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT62), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n985), .A2(new_n995), .A3(new_n990), .A4(new_n991), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n839), .A2(KEYINPUT45), .A3(new_n926), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT113), .B1(new_n961), .B2(KEYINPUT45), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n967), .A2(new_n1000), .A3(new_n928), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n998), .A2(new_n930), .A3(new_n999), .A4(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n997), .B1(new_n1002), .B2(G2078), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n966), .B1(new_n927), .B2(new_n928), .ZN(new_n1004));
  INV_X1    g579(.A(G2078), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1004), .A2(KEYINPUT53), .A3(new_n1005), .A4(new_n962), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n969), .A2(new_n972), .A3(new_n974), .ZN(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT121), .B(G1961), .Z(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1003), .A2(new_n1006), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(G171), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n996), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(G303), .A2(G8), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT55), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n930), .B1(new_n967), .B2(KEYINPUT50), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n927), .B2(KEYINPUT50), .ZN(new_n1018));
  INV_X1    g593(.A(G2090), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n1002), .A2(new_n689), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n958), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1002), .A2(new_n689), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT116), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1016), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n982), .A2(new_n1019), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n1023), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(G8), .A3(new_n1016), .ZN(new_n1030));
  XOR2_X1   g605(.A(new_n583), .B(G1981), .Z(new_n1031));
  XNOR2_X1  g606(.A(new_n1031), .B(KEYINPUT49), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n934), .A2(new_n930), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(G8), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1976), .ZN(new_n1035));
  NOR2_X1   g610(.A1(G288), .A2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1036), .B(KEYINPUT115), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(new_n1033), .A3(G8), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT52), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT52), .B1(G288), .B2(new_n1035), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1037), .A2(new_n1033), .A3(G8), .A4(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1034), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1030), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT122), .B1(new_n1027), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(G8), .B1(new_n1025), .B2(KEYINPUT116), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1015), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT122), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n958), .B1(new_n1028), .B2(new_n1023), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1042), .B1(new_n1050), .B2(new_n1016), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1048), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1045), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT124), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n992), .A2(new_n1054), .A3(KEYINPUT62), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n994), .A2(new_n1013), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1033), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1057), .A2(new_n958), .ZN(new_n1058));
  AOI211_X1 g633(.A(G1976), .B(G288), .C1(new_n1058), .C2(new_n1032), .ZN(new_n1059));
  NOR2_X1   g634(.A1(G305), .A2(G1981), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n1030), .B2(new_n1042), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1048), .A2(G168), .A3(new_n1051), .A4(new_n976), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT63), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n987), .A2(new_n1064), .A3(G286), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1051), .B(new_n1066), .C1(new_n1016), .C2(new_n1050), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1062), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1056), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G1956), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n934), .A2(new_n971), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1070), .B1(new_n1071), .B2(new_n1017), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n961), .A2(KEYINPUT45), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n966), .B1(new_n1073), .B2(new_n1000), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT56), .B(G2072), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(new_n998), .A3(new_n999), .A4(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n567), .B(KEYINPUT57), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1072), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1348), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1007), .A2(new_n1079), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n934), .A2(new_n943), .A3(new_n930), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n608), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1072), .A2(new_n1076), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1077), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1078), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT61), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1077), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1089), .B1(new_n1078), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1072), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1087), .A2(KEYINPUT61), .A3(new_n1092), .ZN(new_n1093));
  XOR2_X1   g668(.A(KEYINPUT117), .B(G1996), .Z(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT58), .B(G1341), .ZN(new_n1095));
  OAI22_X1  g670(.A1(new_n1002), .A2(new_n1094), .B1(new_n1057), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n550), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1096), .A2(KEYINPUT59), .A3(new_n550), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1091), .A2(new_n1093), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT60), .ZN(new_n1103));
  AOI211_X1 g678(.A(new_n1103), .B(new_n1081), .C1(new_n1007), .C2(new_n1079), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1102), .B1(new_n1104), .B2(new_n600), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n600), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1080), .A2(KEYINPUT60), .A3(new_n1082), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1107), .A2(KEYINPUT119), .A3(new_n608), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1083), .A2(new_n1103), .ZN(new_n1110));
  AOI22_X1  g685(.A1(KEYINPUT118), .A2(new_n1101), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1112), .A2(new_n1113), .A3(new_n1093), .A4(new_n1091), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1088), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1004), .A2(KEYINPUT53), .A3(new_n1005), .A4(new_n998), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1003), .A2(new_n1009), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(G171), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1003), .A2(new_n1006), .A3(new_n1009), .A4(G301), .ZN(new_n1120));
  AND4_X1   g695(.A1(new_n1116), .A2(new_n1119), .A3(KEYINPUT54), .A4(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1122), .B1(new_n1118), .B2(G171), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1116), .B1(new_n1123), .B2(new_n1120), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n978), .A2(new_n984), .B1(new_n986), .B2(new_n988), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1011), .B1(G171), .B2(new_n1118), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n990), .A2(new_n1126), .B1(new_n1127), .B2(new_n1122), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1053), .A2(new_n1125), .A3(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1115), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n957), .B1(new_n1069), .B2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n942), .A2(new_n946), .A3(new_n952), .A4(new_n950), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n797), .A2(G2067), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n941), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n947), .A2(G1986), .A3(G290), .ZN(new_n1136));
  XOR2_X1   g711(.A(new_n1136), .B(KEYINPUT48), .Z(new_n1137));
  NAND3_X1  g712(.A1(new_n1137), .A2(new_n951), .A3(new_n954), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT47), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n938), .A2(KEYINPUT112), .A3(new_n939), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT112), .B1(new_n938), .B2(new_n939), .ZN(new_n1141));
  OAI22_X1  g716(.A1(new_n1140), .A2(new_n1141), .B1(new_n768), .B2(new_n945), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n941), .B(KEYINPUT125), .C1(new_n768), .C2(new_n945), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n938), .A2(new_n949), .A3(new_n939), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT46), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1147), .B(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1139), .B1(new_n1146), .B2(new_n1150), .ZN(new_n1151));
  AOI211_X1 g726(.A(KEYINPUT47), .B(new_n1149), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1135), .B(new_n1138), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT126), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1146), .A2(new_n1150), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(KEYINPUT47), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1146), .A2(new_n1139), .A3(new_n1150), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1158), .A2(new_n1159), .A3(new_n1135), .A4(new_n1138), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1154), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1131), .A2(new_n1161), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g737(.A1(new_n659), .A2(G319), .ZN(new_n1164));
  NOR2_X1   g738(.A1(new_n1164), .A2(G401), .ZN(new_n1165));
  XNOR2_X1  g739(.A(new_n1165), .B(KEYINPUT127), .ZN(new_n1166));
  NOR2_X1   g740(.A1(new_n1166), .A2(G229), .ZN(new_n1167));
  OAI21_X1  g741(.A(new_n1167), .B1(new_n921), .B2(new_n922), .ZN(new_n1168));
  AOI21_X1  g742(.A(new_n1168), .B1(new_n867), .B2(new_n868), .ZN(G308));
  OAI221_X1 g743(.A(new_n1167), .B1(new_n921), .B2(new_n922), .C1(new_n861), .C2(new_n864), .ZN(G225));
endmodule


