//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n629, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n462));
  AND3_X1   g037(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(KEYINPUT3), .B1(new_n462), .B2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n461), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n471), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n470), .B1(new_n472), .B2(new_n461), .ZN(new_n473));
  AND2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(G125), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(KEYINPUT66), .A3(G2105), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n469), .B1(new_n473), .B2(new_n479), .ZN(G160));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n481), .B1(new_n466), .B2(KEYINPUT67), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n461), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(G2105), .B1(new_n482), .B2(new_n483), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(G136), .B2(new_n489), .ZN(G162));
  OAI211_X1 g065(.A(G138), .B(new_n461), .C1(new_n474), .C2(new_n475), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  OR2_X1    g067(.A1(new_n461), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n491), .A2(new_n492), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(KEYINPUT4), .A2(G138), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n461), .B(new_n497), .C1(new_n463), .C2(new_n464), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n482), .A2(new_n483), .ZN(new_n500));
  NAND2_X1  g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n499), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  AOI211_X1 g078(.A(KEYINPUT68), .B(new_n501), .C1(new_n482), .C2(new_n483), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n496), .B(new_n498), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G62), .ZN(new_n511));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n507), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  OAI21_X1  g094(.A(G543), .B1(new_n516), .B2(new_n517), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n513), .A2(new_n522), .ZN(G166));
  NOR2_X1   g098(.A1(new_n515), .A2(new_n514), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n516), .A2(new_n517), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n526), .A2(G89), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n510), .A2(KEYINPUT69), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT69), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n524), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n520), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G51), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n530), .A2(new_n535), .A3(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  AOI22_X1  g114(.A1(new_n526), .A2(G90), .B1(new_n536), .B2(G52), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n531), .A2(new_n533), .A3(G64), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n507), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n540), .B1(new_n543), .B2(KEYINPUT70), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT70), .ZN(new_n546));
  AOI211_X1 g121(.A(new_n546), .B(new_n507), .C1(new_n541), .C2(new_n542), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n545), .A2(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND3_X1  g125(.A1(new_n531), .A2(new_n533), .A3(G56), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  INV_X1    g130(.A(G43), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n518), .A2(new_n555), .B1(new_n520), .B2(new_n556), .ZN(new_n557));
  AND2_X1   g132(.A1(new_n557), .A2(KEYINPUT71), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n557), .A2(KEYINPUT71), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n554), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OR3_X1    g142(.A1(new_n520), .A2(KEYINPUT9), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT9), .B1(new_n520), .B2(new_n567), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n524), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(G651), .A2(new_n573), .B1(new_n526), .B2(G91), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(G299));
  OR2_X1    g150(.A1(new_n513), .A2(new_n522), .ZN(G303));
  INV_X1    g151(.A(G74), .ZN(new_n577));
  NOR3_X1   g152(.A1(new_n515), .A2(new_n514), .A3(KEYINPUT69), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n532), .B1(new_n508), .B2(new_n509), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT72), .ZN(new_n582));
  INV_X1    g157(.A(G87), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n518), .B2(new_n583), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n516), .A2(new_n517), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n585), .A2(KEYINPUT72), .A3(G87), .A4(new_n510), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n536), .A2(G49), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n581), .A2(new_n587), .A3(new_n588), .ZN(G288));
  INV_X1    g164(.A(G86), .ZN(new_n590));
  INV_X1    g165(.A(G48), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n518), .A2(new_n590), .B1(new_n520), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(G61), .B1(new_n515), .B2(new_n514), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n507), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G305));
  NAND3_X1  g172(.A1(new_n531), .A2(new_n533), .A3(G60), .ZN(new_n598));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n507), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n526), .A2(G85), .B1(new_n536), .B2(G47), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n526), .A2(KEYINPUT10), .A3(G92), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n518), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G54), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(new_n520), .B2(KEYINPUT73), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT73), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n585), .A2(new_n613), .A3(G543), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n524), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n612), .A2(new_n614), .B1(new_n617), .B2(G651), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n610), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT74), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n605), .B1(new_n622), .B2(G868), .ZN(G284));
  OAI21_X1  g198(.A(new_n605), .B1(new_n622), .B2(G868), .ZN(G321));
  NAND2_X1  g199(.A1(G286), .A2(G868), .ZN(new_n625));
  AND2_X1   g200(.A1(new_n570), .A2(new_n574), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(G297));
  OAI21_X1  g202(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n622), .B1(new_n629), .B2(G860), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT75), .ZN(G148));
  NAND2_X1  g206(.A1(new_n622), .A2(new_n629), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n561), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n484), .A2(G123), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n489), .A2(G135), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n461), .A2(G111), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  NAND3_X1  g216(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT12), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT13), .Z(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(G2100), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(G2100), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n641), .A2(new_n645), .A3(new_n646), .ZN(G156));
  INV_X1    g222(.A(KEYINPUT14), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(new_n651), .B2(new_n650), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n653), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(G14), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT76), .Z(G401));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT17), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n667), .B2(new_n664), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n668), .B1(KEYINPUT77), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(KEYINPUT77), .B2(new_n670), .ZN(new_n672));
  INV_X1    g247(.A(new_n664), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n673), .A2(new_n669), .A3(new_n666), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT18), .Z(new_n675));
  NAND3_X1  g250(.A1(new_n665), .A2(new_n669), .A3(new_n667), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n672), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2096), .B(G2100), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(G1971), .B(G1976), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  AND2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT20), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n682), .A2(new_n683), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n681), .A2(new_n684), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n681), .B2(new_n687), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT78), .Z(new_n691));
  XOR2_X1   g266(.A(G1981), .B(G1986), .Z(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n691), .B(new_n696), .ZN(G229));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G26), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT28), .Z(new_n700));
  NAND2_X1  g275(.A1(new_n484), .A2(G128), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n489), .A2(G140), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n461), .A2(G116), .ZN(new_n703));
  OAI21_X1  g278(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n701), .B(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT83), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n700), .B1(new_n706), .B2(G29), .ZN(new_n707));
  INV_X1    g282(.A(G2067), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n710), .A2(G4), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n621), .B2(G16), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT82), .B(G1348), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT93), .ZN(new_n715));
  NOR2_X1   g290(.A1(G29), .A2(G35), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G162), .B2(G29), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G2090), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI211_X1 g296(.A(new_n709), .B(new_n714), .C1(new_n715), .C2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT24), .ZN(new_n723));
  INV_X1    g298(.A(G34), .ZN(new_n724));
  AOI21_X1  g299(.A(G29), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(new_n723), .B2(new_n724), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G160), .B2(new_n698), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT88), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G2084), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n721), .B2(new_n715), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n710), .A2(G19), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n561), .B2(new_n710), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n732), .A2(G1341), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n698), .A2(G27), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G164), .B2(new_n698), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n732), .A2(G1341), .B1(G2078), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT30), .B(G28), .ZN(new_n738));
  OR2_X1    g313(.A1(KEYINPUT31), .A2(G11), .ZN(new_n739));
  NAND2_X1  g314(.A1(KEYINPUT31), .A2(G11), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n738), .A2(new_n698), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n710), .A2(G21), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G286), .B2(G16), .ZN(new_n743));
  INV_X1    g318(.A(G1966), .ZN(new_n744));
  OAI221_X1 g319(.A(new_n741), .B1(new_n698), .B2(new_n640), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT26), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n750), .A2(new_n751), .B1(G105), .B2(new_n467), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n489), .A2(G141), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n484), .A2(G129), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G29), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n757), .B(KEYINPUT89), .C1(G29), .C2(G32), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(KEYINPUT89), .B2(new_n757), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT27), .B(G1996), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  OAI22_X1  g336(.A1(new_n759), .A2(new_n761), .B1(G2078), .B2(new_n735), .ZN(new_n762));
  NOR4_X1   g337(.A1(new_n730), .A2(new_n737), .A3(new_n747), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n710), .A2(G20), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT23), .Z(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G299), .B2(G16), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1956), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n719), .B2(new_n720), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT94), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n710), .A2(G5), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G301), .B2(G16), .ZN(new_n771));
  INV_X1    g346(.A(G1961), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT90), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n722), .A2(new_n763), .A3(new_n769), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G29), .A2(G33), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT84), .B(KEYINPUT25), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G139), .B2(new_n489), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n471), .A2(G127), .ZN(new_n781));
  INV_X1    g356(.A(G115), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(new_n466), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(KEYINPUT85), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(G2105), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n783), .A2(KEYINPUT85), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n780), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT86), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(KEYINPUT87), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n787), .B(KEYINPUT86), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT87), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n776), .B1(new_n794), .B2(G29), .ZN(new_n795));
  INV_X1    g370(.A(G2072), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n771), .A2(new_n772), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n759), .A2(new_n761), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n798), .B(new_n799), .C1(new_n728), .C2(G2084), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT91), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n775), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n710), .A2(G24), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT80), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n603), .B2(new_n710), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(G1986), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n484), .A2(G119), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n489), .A2(G131), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n461), .A2(G107), .ZN(new_n810));
  OAI21_X1  g385(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n808), .B(new_n809), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  MUX2_X1   g387(.A(G25), .B(new_n812), .S(G29), .Z(new_n813));
  XOR2_X1   g388(.A(KEYINPUT35), .B(G1991), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT79), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n813), .B(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n806), .A2(G1986), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AND3_X1   g393(.A1(new_n581), .A2(new_n587), .A3(new_n588), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(new_n710), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(new_n710), .B2(G23), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT33), .B(G1976), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(G6), .A2(G16), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n596), .B2(G16), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT32), .B(G1981), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n821), .B2(new_n822), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n710), .A2(G22), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(G166), .B2(new_n710), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G1971), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT81), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n823), .A2(new_n828), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n807), .B(new_n818), .C1(new_n835), .C2(KEYINPUT34), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n835), .A2(KEYINPUT34), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT36), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  AND3_X1   g415(.A1(new_n803), .A2(new_n840), .A3(KEYINPUT95), .ZN(new_n841));
  AOI21_X1  g416(.A(KEYINPUT95), .B1(new_n803), .B2(new_n840), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(G311));
  AND3_X1   g418(.A1(new_n803), .A2(new_n840), .A3(KEYINPUT96), .ZN(new_n844));
  AOI21_X1  g419(.A(KEYINPUT96), .B1(new_n803), .B2(new_n840), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(G150));
  INV_X1    g421(.A(KEYINPUT97), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT71), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n557), .B(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n507), .B1(new_n551), .B2(new_n552), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n531), .A2(new_n533), .A3(G67), .ZN(new_n852));
  NAND2_X1  g427(.A1(G80), .A2(G543), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n507), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(G93), .ZN(new_n855));
  INV_X1    g430(.A(G55), .ZN(new_n856));
  OAI22_X1  g431(.A1(new_n518), .A2(new_n855), .B1(new_n520), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n554), .B(KEYINPUT97), .C1(new_n558), .C2(new_n559), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n851), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n560), .B(new_n847), .C1(new_n854), .C2(new_n857), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT38), .Z(new_n863));
  NOR2_X1   g438(.A1(new_n621), .A2(new_n629), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n866));
  AOI21_X1  g441(.A(G860), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n866), .B2(new_n865), .ZN(new_n868));
  OAI21_X1  g443(.A(G860), .B1(new_n854), .B2(new_n857), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT37), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(G145));
  NAND2_X1  g446(.A1(new_n484), .A2(G130), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n461), .A2(G118), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(G142), .B2(new_n489), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(new_n643), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n812), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n706), .A2(G164), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n706), .A2(G164), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n755), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n881), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n883), .A2(new_n756), .A3(new_n879), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n884), .A3(new_n791), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI22_X1  g461(.A1(new_n882), .A2(new_n884), .B1(new_n790), .B2(new_n793), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n878), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n882), .A2(new_n884), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n794), .ZN(new_n890));
  INV_X1    g465(.A(new_n878), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(new_n891), .A3(new_n885), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(G162), .B(new_n640), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(G160), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT98), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT98), .ZN(new_n897));
  INV_X1    g472(.A(new_n895), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n888), .A2(new_n892), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(G37), .B1(new_n893), .B2(new_n895), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT40), .ZN(G395));
  AND2_X1   g478(.A1(new_n610), .A2(new_n618), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n626), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n619), .A2(G299), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n908), .A2(KEYINPUT99), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n619), .A2(G299), .ZN(new_n910));
  AOI22_X1  g485(.A1(new_n610), .A2(new_n618), .B1(new_n570), .B2(new_n574), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT41), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n912), .A2(new_n908), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n909), .B1(new_n913), .B2(KEYINPUT99), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n910), .A2(new_n911), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n632), .B(new_n862), .ZN(new_n916));
  MUX2_X1   g491(.A(new_n914), .B(new_n915), .S(new_n916), .Z(new_n917));
  NAND2_X1  g492(.A1(new_n598), .A2(new_n599), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(G651), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n919), .A2(G303), .A3(new_n601), .ZN(new_n920));
  OAI21_X1  g495(.A(G166), .B1(new_n600), .B2(new_n602), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(G288), .A2(new_n596), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(G288), .A2(new_n596), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n819), .A2(G305), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n927), .A2(new_n921), .A3(new_n920), .A4(new_n923), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT42), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n926), .A2(KEYINPUT100), .A3(new_n928), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT100), .B1(new_n926), .B2(new_n928), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n929), .B1(new_n933), .B2(KEYINPUT42), .ZN(new_n934));
  XOR2_X1   g509(.A(new_n917), .B(new_n934), .Z(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(G868), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(G868), .B2(new_n858), .ZN(G295));
  OAI21_X1  g512(.A(new_n936), .B1(G868), .B2(new_n858), .ZN(G331));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT101), .ZN(new_n941));
  NAND2_X1  g516(.A1(G286), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n530), .A2(KEYINPUT101), .A3(new_n535), .A4(new_n537), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n944), .A2(new_n545), .A3(new_n548), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n942), .B(new_n943), .C1(new_n544), .C2(new_n547), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n862), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n860), .A2(new_n945), .A3(new_n861), .A4(new_n946), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n914), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n915), .A3(new_n949), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n932), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G37), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n912), .A2(new_n908), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n950), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n957), .A2(KEYINPUT104), .A3(new_n952), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT104), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n913), .B1(new_n948), .B2(new_n949), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n932), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n958), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n962), .B1(new_n958), .B2(new_n961), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n940), .B(new_n955), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT99), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n915), .A2(new_n966), .A3(new_n906), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(new_n956), .B2(new_n966), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n968), .B1(new_n949), .B2(new_n948), .ZN(new_n969));
  INV_X1    g544(.A(new_n952), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT102), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT102), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n951), .A2(new_n972), .A3(new_n952), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(new_n933), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n940), .B1(new_n974), .B2(new_n955), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT103), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n965), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI211_X1 g552(.A(KEYINPUT103), .B(new_n940), .C1(new_n974), .C2(new_n955), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n939), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n955), .B1(new_n963), .B2(new_n964), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(new_n940), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT43), .B1(new_n974), .B2(new_n955), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT44), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n979), .A2(new_n983), .ZN(G397));
  INV_X1    g559(.A(G1384), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n503), .A2(new_n504), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n491), .A2(new_n492), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n493), .A2(new_n495), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(new_n498), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n985), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n489), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT66), .B1(new_n478), .B2(G2105), .ZN(new_n994));
  AOI211_X1 g569(.A(new_n470), .B(new_n461), .C1(new_n476), .C2(new_n477), .ZN(new_n995));
  OAI211_X1 g570(.A(G40), .B(new_n993), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n706), .B(new_n708), .ZN(new_n998));
  XOR2_X1   g573(.A(new_n755), .B(G1996), .Z(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n812), .A2(new_n815), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n812), .A2(new_n815), .ZN(new_n1002));
  OR3_X1    g577(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1986), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n603), .B(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n997), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n505), .A2(new_n1007), .A3(new_n985), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1007), .B1(new_n505), .B2(new_n985), .ZN(new_n1010));
  NOR4_X1   g585(.A1(new_n1009), .A2(new_n1010), .A3(G2084), .A4(new_n996), .ZN(new_n1011));
  INV_X1    g586(.A(new_n996), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n992), .A2(KEYINPUT118), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT118), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT45), .B1(new_n505), .B2(new_n985), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1014), .B1(new_n1015), .B2(new_n996), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n985), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1013), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1011), .B1(new_n1018), .B2(new_n744), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT108), .B(G8), .Z(new_n1020));
  NOR3_X1   g595(.A1(new_n1019), .A2(G286), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G8), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n992), .A2(new_n1012), .A3(new_n1017), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT106), .ZN(new_n1025));
  INV_X1    g600(.A(G1971), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT106), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n992), .A2(new_n1012), .A3(new_n1027), .A4(new_n1017), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1025), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n996), .B1(KEYINPUT50), .B2(new_n990), .ZN(new_n1030));
  XOR2_X1   g605(.A(KEYINPUT107), .B(G2090), .Z(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(new_n1008), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1023), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G303), .A2(G8), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1034), .B(KEYINPUT55), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1022), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT63), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1020), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n990), .B2(new_n996), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n581), .A2(new_n587), .A3(G1976), .A4(new_n588), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT52), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT109), .B(G1976), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT52), .B1(G288), .B2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(G160), .A2(G40), .A3(new_n985), .A4(new_n505), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1047), .A2(new_n1048), .A3(new_n1041), .A4(new_n1043), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(G1981), .B1(new_n592), .B2(new_n595), .ZN(new_n1051));
  INV_X1    g626(.A(G61), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n508), .B2(new_n509), .ZN(new_n1053));
  INV_X1    g628(.A(new_n594), .ZN(new_n1054));
  OAI21_X1  g629(.A(G651), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n585), .A2(G86), .A3(new_n510), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n585), .A2(G48), .A3(G543), .ZN(new_n1057));
  INV_X1    g632(.A(G1981), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1051), .A2(KEYINPUT110), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT111), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT49), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT110), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(KEYINPUT111), .B2(KEYINPUT49), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(new_n1051), .B2(new_n1059), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1042), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1040), .B1(new_n1050), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT49), .B1(new_n1060), .B2(KEYINPUT111), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1041), .B(new_n1048), .C1(new_n1070), .C2(new_n1066), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1071), .A2(KEYINPUT112), .A3(new_n1049), .A4(new_n1045), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1039), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1074), .A2(G8), .A3(new_n1036), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1038), .A2(KEYINPUT119), .A3(new_n1073), .A4(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT117), .B1(new_n1050), .B2(new_n1068), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1071), .A2(new_n1078), .A3(new_n1049), .A4(new_n1045), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1009), .B1(new_n1030), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT116), .B1(new_n1010), .B2(new_n996), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n1031), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1020), .B1(new_n1029), .B2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1075), .B(new_n1080), .C1(new_n1036), .C2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1039), .B1(new_n1086), .B2(new_n1022), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1021), .B1(new_n1036), .B2(new_n1033), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1076), .A2(new_n1087), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1075), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1042), .B(KEYINPUT113), .ZN(new_n1094));
  NOR2_X1   g669(.A1(G288), .A2(G1976), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1095), .B(KEYINPUT115), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n1071), .ZN(new_n1097));
  XOR2_X1   g672(.A(new_n1059), .B(KEYINPUT114), .Z(new_n1098));
  AOI21_X1  g673(.A(new_n1094), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1093), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(G168), .A2(new_n1020), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT51), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1101), .A2(KEYINPUT51), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1019), .A2(new_n1102), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT124), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(new_n1019), .B2(new_n1102), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1086), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1114), .A2(G2078), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1013), .A2(new_n1016), .A3(new_n1017), .A4(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n990), .A2(KEYINPUT50), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1117), .A2(new_n1012), .A3(new_n1008), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n772), .ZN(new_n1119));
  AOI21_X1  g694(.A(G2078), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1116), .B(new_n1119), .C1(new_n1120), .C2(KEYINPUT53), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1121), .A2(G171), .ZN(new_n1122));
  OAI211_X1 g697(.A(G40), .B(new_n1115), .C1(new_n472), .C2(new_n461), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1123), .A2(new_n469), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n992), .A2(new_n1124), .A3(new_n1017), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1119), .B(new_n1125), .C1(new_n1120), .C2(KEYINPUT53), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1126), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT125), .B1(new_n1126), .B2(G171), .ZN(new_n1128));
  OAI211_X1 g703(.A(KEYINPUT54), .B(new_n1122), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT54), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1121), .A2(G171), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1126), .A2(G171), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1113), .A2(new_n1129), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(G1956), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n626), .B(KEYINPUT57), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(KEYINPUT56), .B(G2072), .ZN(new_n1138));
  AND4_X1   g713(.A1(new_n1012), .A2(new_n992), .A3(new_n1017), .A4(new_n1138), .ZN(new_n1139));
  NOR4_X1   g714(.A1(new_n1135), .A2(KEYINPUT120), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT120), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1117), .A2(new_n1081), .A3(new_n1012), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1142), .A2(new_n1083), .A3(new_n1008), .ZN(new_n1143));
  INV_X1    g718(.A(G1956), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1139), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1141), .B1(new_n1145), .B2(new_n1136), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1140), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1137), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1148));
  INV_X1    g723(.A(G1348), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1118), .A2(new_n1149), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n1048), .A2(G2067), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n619), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1148), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1147), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1145), .B2(new_n1136), .ZN(new_n1158));
  OAI211_X1 g733(.A(KEYINPUT123), .B(new_n1137), .C1(new_n1135), .C2(new_n1139), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1156), .B1(new_n1147), .B2(new_n1160), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1150), .A2(new_n1151), .A3(new_n619), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT60), .B1(new_n1162), .B2(new_n1152), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n619), .A2(KEYINPUT60), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1150), .A2(new_n1151), .A3(new_n1164), .ZN(new_n1165));
  XOR2_X1   g740(.A(KEYINPUT121), .B(G1996), .Z(new_n1166));
  NAND4_X1  g741(.A1(new_n992), .A2(new_n1012), .A3(new_n1017), .A4(new_n1166), .ZN(new_n1167));
  XOR2_X1   g742(.A(KEYINPUT58), .B(G1341), .Z(new_n1168));
  AOI22_X1  g743(.A1(new_n1167), .A2(KEYINPUT122), .B1(new_n1048), .B2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1015), .A2(new_n996), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT122), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1170), .A2(new_n1171), .A3(new_n1017), .A4(new_n1166), .ZN(new_n1172));
  AOI211_X1 g747(.A(KEYINPUT59), .B(new_n560), .C1(new_n1169), .C2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT59), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1167), .A2(KEYINPUT122), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1048), .A2(new_n1168), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1175), .A2(new_n1172), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1174), .B1(new_n1177), .B2(new_n561), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1163), .B(new_n1165), .C1(new_n1173), .C2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1145), .A2(new_n1136), .ZN(new_n1180));
  AND3_X1   g755(.A1(new_n1148), .A2(new_n1180), .A3(KEYINPUT61), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1155), .B1(new_n1161), .B2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g758(.A(new_n1092), .B(new_n1100), .C1(new_n1134), .C2(new_n1183), .ZN(new_n1184));
  OR2_X1    g759(.A1(new_n1085), .A2(new_n1036), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1033), .A2(new_n1036), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1131), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n1188));
  AOI22_X1  g763(.A1(new_n1104), .A2(new_n1106), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1191), .A2(new_n1192), .A3(KEYINPUT62), .ZN(new_n1193));
  OAI21_X1  g768(.A(KEYINPUT126), .B1(new_n1189), .B2(new_n1188), .ZN(new_n1194));
  AND3_X1   g769(.A1(new_n1190), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1006), .B1(new_n1184), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(new_n997), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1197), .B1(new_n998), .B2(new_n756), .ZN(new_n1198));
  OAI21_X1  g773(.A(KEYINPUT46), .B1(new_n1197), .B2(G1996), .ZN(new_n1199));
  OR3_X1    g774(.A1(new_n1197), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1198), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT47), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n706), .A2(G2067), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1000), .A2(new_n997), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1203), .B1(new_n1204), .B2(new_n1002), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n1206));
  AND2_X1   g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1208));
  NOR3_X1   g783(.A1(new_n1207), .A2(new_n1208), .A3(new_n1197), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1003), .A2(new_n997), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n997), .A2(new_n1004), .A3(new_n603), .ZN(new_n1211));
  XNOR2_X1  g786(.A(new_n1211), .B(KEYINPUT48), .ZN(new_n1212));
  AOI211_X1 g787(.A(new_n1202), .B(new_n1209), .C1(new_n1210), .C2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1196), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g789(.A1(G401), .A2(G229), .A3(new_n459), .A4(G227), .ZN(new_n1216));
  OAI211_X1 g790(.A(new_n902), .B(new_n1216), .C1(new_n977), .C2(new_n978), .ZN(G225));
  INV_X1    g791(.A(G225), .ZN(G308));
endmodule


