

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585;

  XOR2_X1 U325 ( .A(n317), .B(n316), .Z(n293) );
  XNOR2_X1 U326 ( .A(KEYINPUT45), .B(KEYINPUT65), .ZN(n347) );
  XNOR2_X1 U327 ( .A(n348), .B(n347), .ZN(n368) );
  XNOR2_X1 U328 ( .A(n318), .B(n293), .ZN(n319) );
  XNOR2_X1 U329 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U330 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U331 ( .A(n328), .B(n327), .ZN(n370) );
  INV_X1 U332 ( .A(G169GAT), .ZN(n457) );
  XNOR2_X1 U333 ( .A(n457), .B(KEYINPUT124), .ZN(n458) );
  XNOR2_X1 U334 ( .A(n459), .B(n458), .ZN(G1348GAT) );
  XOR2_X1 U335 ( .A(G22GAT), .B(G197GAT), .Z(n295) );
  XNOR2_X1 U336 ( .A(G43GAT), .B(G141GAT), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U338 ( .A(n296), .B(G36GAT), .Z(n298) );
  XOR2_X1 U339 ( .A(G1GAT), .B(KEYINPUT73), .Z(n344) );
  XNOR2_X1 U340 ( .A(n344), .B(G50GAT), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n298), .B(n297), .ZN(n304) );
  XOR2_X1 U342 ( .A(G29GAT), .B(KEYINPUT7), .Z(n300) );
  XNOR2_X1 U343 ( .A(KEYINPUT72), .B(KEYINPUT8), .ZN(n299) );
  XNOR2_X1 U344 ( .A(n300), .B(n299), .ZN(n313) );
  XOR2_X1 U345 ( .A(G113GAT), .B(G15GAT), .Z(n451) );
  XOR2_X1 U346 ( .A(n313), .B(n451), .Z(n302) );
  NAND2_X1 U347 ( .A1(G229GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U349 ( .A(n304), .B(n303), .Z(n312) );
  XOR2_X1 U350 ( .A(KEYINPUT71), .B(KEYINPUT74), .Z(n306) );
  XNOR2_X1 U351 ( .A(G169GAT), .B(G8GAT), .ZN(n305) );
  XNOR2_X1 U352 ( .A(n306), .B(n305), .ZN(n310) );
  XOR2_X1 U353 ( .A(KEYINPUT29), .B(KEYINPUT70), .Z(n308) );
  XNOR2_X1 U354 ( .A(KEYINPUT69), .B(KEYINPUT30), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U356 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U357 ( .A(n312), .B(n311), .Z(n507) );
  INV_X1 U358 ( .A(n507), .ZN(n571) );
  XOR2_X1 U359 ( .A(G85GAT), .B(G92GAT), .Z(n352) );
  XNOR2_X1 U360 ( .A(n313), .B(n352), .ZN(n315) );
  AND2_X1 U361 ( .A1(G232GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U362 ( .A(n315), .B(n314), .ZN(n320) );
  XOR2_X1 U363 ( .A(G43GAT), .B(G134GAT), .Z(n440) );
  XOR2_X1 U364 ( .A(G36GAT), .B(G190GAT), .Z(n383) );
  XNOR2_X1 U365 ( .A(n440), .B(n383), .ZN(n318) );
  XOR2_X1 U366 ( .A(KEYINPUT81), .B(KEYINPUT66), .Z(n317) );
  XNOR2_X1 U367 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n316) );
  XOR2_X1 U368 ( .A(n321), .B(G106GAT), .Z(n328) );
  XNOR2_X1 U369 ( .A(G50GAT), .B(KEYINPUT80), .ZN(n322) );
  XNOR2_X1 U370 ( .A(n322), .B(G162GAT), .ZN(n433) );
  XNOR2_X1 U371 ( .A(G99GAT), .B(n433), .ZN(n326) );
  XOR2_X1 U372 ( .A(KEYINPUT82), .B(KEYINPUT9), .Z(n324) );
  XNOR2_X1 U373 ( .A(KEYINPUT67), .B(KEYINPUT11), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U375 ( .A(n370), .B(KEYINPUT36), .Z(n583) );
  XOR2_X1 U376 ( .A(G8GAT), .B(KEYINPUT83), .Z(n380) );
  XOR2_X1 U377 ( .A(n380), .B(KEYINPUT86), .Z(n330) );
  NAND2_X1 U378 ( .A1(G231GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U379 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U380 ( .A(KEYINPUT12), .B(KEYINPUT85), .Z(n332) );
  XNOR2_X1 U381 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U383 ( .A(n334), .B(n333), .Z(n339) );
  XOR2_X1 U384 ( .A(G22GAT), .B(G155GAT), .Z(n423) );
  XOR2_X1 U385 ( .A(KEYINPUT84), .B(G64GAT), .Z(n336) );
  XNOR2_X1 U386 ( .A(G15GAT), .B(G71GAT), .ZN(n335) );
  XNOR2_X1 U387 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U388 ( .A(n423), .B(n337), .ZN(n338) );
  XNOR2_X1 U389 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U390 ( .A(G78GAT), .B(G211GAT), .Z(n341) );
  XNOR2_X1 U391 ( .A(G183GAT), .B(G127GAT), .ZN(n340) );
  XNOR2_X1 U392 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U393 ( .A(n343), .B(n342), .Z(n346) );
  XOR2_X1 U394 ( .A(G57GAT), .B(KEYINPUT13), .Z(n353) );
  XNOR2_X1 U395 ( .A(n344), .B(n353), .ZN(n345) );
  XOR2_X1 U396 ( .A(n346), .B(n345), .Z(n560) );
  INV_X1 U397 ( .A(n560), .ZN(n580) );
  NAND2_X1 U398 ( .A1(n583), .A2(n580), .ZN(n348) );
  XOR2_X1 U399 ( .A(G78GAT), .B(G148GAT), .Z(n350) );
  XNOR2_X1 U400 ( .A(G106GAT), .B(G204GAT), .ZN(n349) );
  XNOR2_X1 U401 ( .A(n350), .B(n349), .ZN(n424) );
  XOR2_X1 U402 ( .A(G99GAT), .B(G71GAT), .Z(n351) );
  XOR2_X1 U403 ( .A(G120GAT), .B(n351), .Z(n444) );
  XOR2_X1 U404 ( .A(n424), .B(n444), .Z(n366) );
  XOR2_X1 U405 ( .A(n353), .B(n352), .Z(n355) );
  NAND2_X1 U406 ( .A1(G230GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U407 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U408 ( .A(KEYINPUT77), .B(KEYINPUT31), .Z(n357) );
  XNOR2_X1 U409 ( .A(KEYINPUT78), .B(KEYINPUT75), .ZN(n356) );
  XNOR2_X1 U410 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U411 ( .A(n359), .B(n358), .Z(n364) );
  XOR2_X1 U412 ( .A(G176GAT), .B(G64GAT), .Z(n390) );
  XOR2_X1 U413 ( .A(KEYINPUT32), .B(KEYINPUT79), .Z(n361) );
  XNOR2_X1 U414 ( .A(KEYINPUT76), .B(KEYINPUT33), .ZN(n360) );
  XNOR2_X1 U415 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U416 ( .A(n390), .B(n362), .ZN(n363) );
  XNOR2_X1 U417 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U418 ( .A(n366), .B(n365), .ZN(n577) );
  NOR2_X1 U419 ( .A1(n577), .A2(n507), .ZN(n367) );
  AND2_X1 U420 ( .A1(n368), .A2(n367), .ZN(n369) );
  XOR2_X1 U421 ( .A(n369), .B(KEYINPUT119), .Z(n378) );
  XNOR2_X1 U422 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n371) );
  XNOR2_X1 U423 ( .A(n371), .B(n577), .ZN(n556) );
  NOR2_X1 U424 ( .A1(n571), .A2(n556), .ZN(n372) );
  XNOR2_X1 U425 ( .A(n372), .B(KEYINPUT46), .ZN(n373) );
  NOR2_X1 U426 ( .A1(n580), .A2(n373), .ZN(n374) );
  NAND2_X1 U427 ( .A1(n370), .A2(n374), .ZN(n375) );
  XNOR2_X1 U428 ( .A(n375), .B(KEYINPUT47), .ZN(n376) );
  XNOR2_X1 U429 ( .A(KEYINPUT118), .B(n376), .ZN(n377) );
  NOR2_X1 U430 ( .A1(n378), .A2(n377), .ZN(n379) );
  XNOR2_X1 U431 ( .A(KEYINPUT48), .B(n379), .ZN(n544) );
  XOR2_X1 U432 ( .A(n380), .B(KEYINPUT104), .Z(n382) );
  NAND2_X1 U433 ( .A1(G226GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U434 ( .A(n382), .B(n381), .ZN(n384) );
  XOR2_X1 U435 ( .A(n384), .B(n383), .Z(n394) );
  XOR2_X1 U436 ( .A(KEYINPUT96), .B(KEYINPUT21), .Z(n386) );
  XNOR2_X1 U437 ( .A(G218GAT), .B(KEYINPUT94), .ZN(n385) );
  XNOR2_X1 U438 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U439 ( .A(n387), .B(KEYINPUT95), .Z(n389) );
  XNOR2_X1 U440 ( .A(G197GAT), .B(G211GAT), .ZN(n388) );
  XNOR2_X1 U441 ( .A(n389), .B(n388), .ZN(n428) );
  XNOR2_X1 U442 ( .A(G204GAT), .B(G92GAT), .ZN(n391) );
  XNOR2_X1 U443 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U444 ( .A(n428), .B(n392), .ZN(n393) );
  XNOR2_X1 U445 ( .A(n394), .B(n393), .ZN(n399) );
  XOR2_X1 U446 ( .A(KEYINPUT92), .B(G183GAT), .Z(n396) );
  XNOR2_X1 U447 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n395) );
  XNOR2_X1 U448 ( .A(n396), .B(n395), .ZN(n398) );
  XOR2_X1 U449 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n397) );
  XOR2_X1 U450 ( .A(n398), .B(n397), .Z(n455) );
  XOR2_X1 U451 ( .A(n399), .B(n455), .Z(n522) );
  NOR2_X1 U452 ( .A1(n544), .A2(n522), .ZN(n400) );
  XNOR2_X1 U453 ( .A(n400), .B(KEYINPUT54), .ZN(n568) );
  XOR2_X1 U454 ( .A(KEYINPUT0), .B(G127GAT), .Z(n441) );
  XOR2_X1 U455 ( .A(G85GAT), .B(G162GAT), .Z(n402) );
  XNOR2_X1 U456 ( .A(G29GAT), .B(G134GAT), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U458 ( .A(n441), .B(n403), .Z(n405) );
  NAND2_X1 U459 ( .A1(G225GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U461 ( .A(n406), .B(KEYINPUT103), .Z(n410) );
  XOR2_X1 U462 ( .A(KEYINPUT97), .B(KEYINPUT3), .Z(n408) );
  XNOR2_X1 U463 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n432) );
  XNOR2_X1 U465 ( .A(G1GAT), .B(n432), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U467 ( .A(G155GAT), .B(G148GAT), .Z(n412) );
  XNOR2_X1 U468 ( .A(G113GAT), .B(G120GAT), .ZN(n411) );
  XNOR2_X1 U469 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U470 ( .A(n414), .B(n413), .Z(n422) );
  XOR2_X1 U471 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n416) );
  XNOR2_X1 U472 ( .A(KEYINPUT1), .B(G57GAT), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U474 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n418) );
  XNOR2_X1 U475 ( .A(KEYINPUT100), .B(KEYINPUT5), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U478 ( .A(n422), .B(n421), .Z(n567) );
  XOR2_X1 U479 ( .A(n423), .B(KEYINPUT22), .Z(n426) );
  XNOR2_X1 U480 ( .A(n424), .B(KEYINPUT98), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U482 ( .A(n428), .B(n427), .ZN(n437) );
  XOR2_X1 U483 ( .A(KEYINPUT24), .B(KEYINPUT99), .Z(n430) );
  NAND2_X1 U484 ( .A1(G228GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U486 ( .A(n431), .B(KEYINPUT23), .Z(n435) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U489 ( .A(n437), .B(n436), .ZN(n467) );
  AND2_X1 U490 ( .A1(n567), .A2(n467), .ZN(n438) );
  NAND2_X1 U491 ( .A1(n568), .A2(n438), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n439), .B(KEYINPUT55), .ZN(n456) );
  XOR2_X1 U493 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U495 ( .A(n443), .B(n442), .ZN(n447) );
  XNOR2_X1 U496 ( .A(n444), .B(KEYINPUT91), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n445), .B(KEYINPUT89), .ZN(n446) );
  XOR2_X1 U498 ( .A(n447), .B(n446), .Z(n453) );
  XOR2_X1 U499 ( .A(KEYINPUT90), .B(KEYINPUT20), .Z(n449) );
  XNOR2_X1 U500 ( .A(G190GAT), .B(G176GAT), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U502 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U503 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U504 ( .A(n455), .B(n454), .Z(n524) );
  INV_X1 U505 ( .A(n524), .ZN(n531) );
  NAND2_X1 U506 ( .A1(n456), .A2(n531), .ZN(n563) );
  NOR2_X1 U507 ( .A1(n571), .A2(n563), .ZN(n459) );
  NOR2_X1 U508 ( .A1(n571), .A2(n577), .ZN(n491) );
  XOR2_X1 U509 ( .A(n524), .B(KEYINPUT93), .Z(n463) );
  INV_X1 U510 ( .A(n522), .ZN(n496) );
  XOR2_X1 U511 ( .A(n496), .B(KEYINPUT105), .Z(n460) );
  XNOR2_X1 U512 ( .A(n460), .B(KEYINPUT27), .ZN(n465) );
  INV_X1 U513 ( .A(n567), .ZN(n493) );
  NAND2_X1 U514 ( .A1(n465), .A2(n493), .ZN(n461) );
  XNOR2_X1 U515 ( .A(n461), .B(KEYINPUT106), .ZN(n545) );
  XOR2_X1 U516 ( .A(n467), .B(KEYINPUT68), .Z(n462) );
  XOR2_X1 U517 ( .A(KEYINPUT28), .B(n462), .Z(n527) );
  INV_X1 U518 ( .A(n527), .ZN(n504) );
  NOR2_X1 U519 ( .A1(n545), .A2(n504), .ZN(n532) );
  NAND2_X1 U520 ( .A1(n463), .A2(n532), .ZN(n473) );
  NOR2_X1 U521 ( .A1(n531), .A2(n467), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n464), .B(KEYINPUT26), .ZN(n569) );
  NAND2_X1 U523 ( .A1(n569), .A2(n465), .ZN(n470) );
  NAND2_X1 U524 ( .A1(n531), .A2(n496), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n467), .A2(n466), .ZN(n468) );
  XOR2_X1 U526 ( .A(KEYINPUT25), .B(n468), .Z(n469) );
  NAND2_X1 U527 ( .A1(n470), .A2(n469), .ZN(n471) );
  NAND2_X1 U528 ( .A1(n471), .A2(n567), .ZN(n472) );
  NAND2_X1 U529 ( .A1(n473), .A2(n472), .ZN(n488) );
  XOR2_X1 U530 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n475) );
  NAND2_X1 U531 ( .A1(n580), .A2(n370), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U533 ( .A(KEYINPUT16), .B(n476), .Z(n477) );
  AND2_X1 U534 ( .A1(n488), .A2(n477), .ZN(n508) );
  NAND2_X1 U535 ( .A1(n491), .A2(n508), .ZN(n485) );
  NOR2_X1 U536 ( .A1(n567), .A2(n485), .ZN(n479) );
  XNOR2_X1 U537 ( .A(KEYINPUT107), .B(KEYINPUT34), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(n480), .ZN(G1324GAT) );
  NOR2_X1 U540 ( .A1(n522), .A2(n485), .ZN(n481) );
  XOR2_X1 U541 ( .A(KEYINPUT108), .B(n481), .Z(n482) );
  XNOR2_X1 U542 ( .A(G8GAT), .B(n482), .ZN(G1325GAT) );
  NOR2_X1 U543 ( .A1(n524), .A2(n485), .ZN(n484) );
  XNOR2_X1 U544 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n484), .B(n483), .ZN(G1326GAT) );
  NOR2_X1 U546 ( .A1(n527), .A2(n485), .ZN(n487) );
  XNOR2_X1 U547 ( .A(G22GAT), .B(KEYINPUT109), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n487), .B(n486), .ZN(G1327GAT) );
  XOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT39), .Z(n495) );
  NAND2_X1 U550 ( .A1(n583), .A2(n488), .ZN(n489) );
  NOR2_X1 U551 ( .A1(n580), .A2(n489), .ZN(n490) );
  XOR2_X1 U552 ( .A(KEYINPUT37), .B(n490), .Z(n520) );
  NAND2_X1 U553 ( .A1(n491), .A2(n520), .ZN(n492) );
  XOR2_X1 U554 ( .A(KEYINPUT38), .B(n492), .Z(n505) );
  NAND2_X1 U555 ( .A1(n493), .A2(n505), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(G1328GAT) );
  NAND2_X1 U557 ( .A1(n505), .A2(n496), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n497), .B(KEYINPUT110), .ZN(n498) );
  XNOR2_X1 U559 ( .A(G36GAT), .B(n498), .ZN(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT40), .B(KEYINPUT113), .Z(n500) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(KEYINPUT112), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U563 ( .A(KEYINPUT111), .B(n501), .Z(n503) );
  NAND2_X1 U564 ( .A1(n505), .A2(n531), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(G1330GAT) );
  NAND2_X1 U566 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n506), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U568 ( .A1(n507), .A2(n556), .ZN(n519) );
  NAND2_X1 U569 ( .A1(n519), .A2(n508), .ZN(n515) );
  NOR2_X1 U570 ( .A1(n567), .A2(n515), .ZN(n510) );
  XNOR2_X1 U571 ( .A(KEYINPUT114), .B(KEYINPUT42), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n511), .Z(G1332GAT) );
  NOR2_X1 U574 ( .A1(n522), .A2(n515), .ZN(n513) );
  XNOR2_X1 U575 ( .A(G64GAT), .B(KEYINPUT115), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n513), .B(n512), .ZN(G1333GAT) );
  NOR2_X1 U577 ( .A1(n524), .A2(n515), .ZN(n514) );
  XOR2_X1 U578 ( .A(G71GAT), .B(n514), .Z(G1334GAT) );
  NOR2_X1 U579 ( .A1(n527), .A2(n515), .ZN(n517) );
  XNOR2_X1 U580 ( .A(KEYINPUT116), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(n518), .ZN(G1335GAT) );
  NAND2_X1 U583 ( .A1(n520), .A2(n519), .ZN(n526) );
  NOR2_X1 U584 ( .A1(n567), .A2(n526), .ZN(n521) );
  XOR2_X1 U585 ( .A(G85GAT), .B(n521), .Z(G1336GAT) );
  NOR2_X1 U586 ( .A1(n522), .A2(n526), .ZN(n523) );
  XOR2_X1 U587 ( .A(G92GAT), .B(n523), .Z(G1337GAT) );
  NOR2_X1 U588 ( .A1(n524), .A2(n526), .ZN(n525) );
  XOR2_X1 U589 ( .A(G99GAT), .B(n525), .Z(G1338GAT) );
  NOR2_X1 U590 ( .A1(n527), .A2(n526), .ZN(n529) );
  XNOR2_X1 U591 ( .A(KEYINPUT44), .B(KEYINPUT117), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(KEYINPUT121), .ZN(n536) );
  NAND2_X1 U595 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U596 ( .A1(n544), .A2(n533), .ZN(n534) );
  XOR2_X1 U597 ( .A(KEYINPUT120), .B(n534), .Z(n541) );
  NOR2_X1 U598 ( .A1(n571), .A2(n541), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n536), .B(n535), .ZN(G1340GAT) );
  NOR2_X1 U600 ( .A1(n541), .A2(n556), .ZN(n538) );
  XNOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  NOR2_X1 U603 ( .A1(n541), .A2(n560), .ZN(n539) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(n539), .Z(n540) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  NOR2_X1 U606 ( .A1(n541), .A2(n370), .ZN(n543) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  NOR2_X1 U609 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U610 ( .A1(n546), .A2(n569), .ZN(n554) );
  NOR2_X1 U611 ( .A1(n571), .A2(n554), .ZN(n547) );
  XOR2_X1 U612 ( .A(KEYINPUT122), .B(n547), .Z(n548) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(n548), .ZN(G1344GAT) );
  NOR2_X1 U614 ( .A1(n556), .A2(n554), .ZN(n550) );
  XNOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(n551), .ZN(G1345GAT) );
  NOR2_X1 U618 ( .A1(n560), .A2(n554), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G155GAT), .B(KEYINPUT123), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1346GAT) );
  NOR2_X1 U621 ( .A1(n370), .A2(n554), .ZN(n555) );
  XOR2_X1 U622 ( .A(G162GAT), .B(n555), .Z(G1347GAT) );
  NOR2_X1 U623 ( .A1(n556), .A2(n563), .ZN(n558) );
  XNOR2_X1 U624 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(n559), .ZN(G1349GAT) );
  NOR2_X1 U627 ( .A1(n560), .A2(n563), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G183GAT), .B(KEYINPUT125), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1350GAT) );
  NOR2_X1 U630 ( .A1(n563), .A2(n370), .ZN(n565) );
  XNOR2_X1 U631 ( .A(KEYINPUT58), .B(KEYINPUT126), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n566) );
  XOR2_X1 U633 ( .A(G190GAT), .B(n566), .Z(G1351GAT) );
  AND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n576) );
  NOR2_X1 U636 ( .A1(n576), .A2(n571), .ZN(n575) );
  XOR2_X1 U637 ( .A(KEYINPUT127), .B(KEYINPUT60), .Z(n573) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .Z(n579) );
  INV_X1 U642 ( .A(n576), .ZN(n582) );
  NAND2_X1 U643 ( .A1(n582), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n582), .A2(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(n584), .B(KEYINPUT62), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

