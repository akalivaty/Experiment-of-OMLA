//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1240, new_n1241, new_n1242, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT65), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n202), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(new_n210), .A2(KEYINPUT0), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n217), .B1(KEYINPUT0), .B2(new_n210), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n225));
  INV_X1    g0025(.A(G50), .ZN(new_n226));
  INV_X1    g0026(.A(G226), .ZN(new_n227));
  INV_X1    g0027(.A(G58), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n225), .B1(new_n226), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n207), .B1(new_n224), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n218), .A2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n211), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(new_n226), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n212), .A2(G33), .ZN(new_n254));
  OAI22_X1  g0054(.A1(new_n254), .A2(new_n222), .B1(new_n212), .B2(G68), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n250), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT11), .ZN(new_n257));
  OR2_X1    g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n260));
  AOI211_X1 g0060(.A(G68), .B(new_n260), .C1(KEYINPUT69), .C2(KEYINPUT12), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n262));
  XNOR2_X1  g0062(.A(new_n261), .B(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n256), .A2(new_n257), .ZN(new_n264));
  INV_X1    g0064(.A(new_n260), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n250), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n266), .B(G68), .C1(G1), .C2(new_n212), .ZN(new_n267));
  AND4_X1   g0067(.A1(new_n258), .A2(new_n263), .A3(new_n264), .A4(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n229), .A2(G1698), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n269), .B1(G226), .B2(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G97), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT13), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G1), .A3(G13), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  INV_X1    g0083(.A(new_n211), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n283), .B1(new_n284), .B2(new_n278), .ZN(new_n285));
  INV_X1    g0085(.A(G41), .ZN(new_n286));
  INV_X1    g0086(.A(G45), .ZN(new_n287));
  AOI21_X1  g0087(.A(G1), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n282), .A2(G238), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n276), .A2(new_n277), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n279), .B1(new_n272), .B2(new_n273), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n288), .A2(new_n279), .A3(G274), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(new_n281), .B2(new_n221), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT13), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G169), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT14), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT14), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n295), .A2(new_n298), .A3(G169), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n290), .A2(new_n294), .A3(G179), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT70), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n290), .A2(new_n294), .A3(KEYINPUT70), .A4(G179), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT71), .B1(new_n300), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n298), .B1(new_n295), .B2(G169), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  AOI211_X1 g0108(.A(KEYINPUT14), .B(new_n308), .C1(new_n290), .C2(new_n294), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT71), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n303), .A2(new_n304), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n268), .B1(new_n306), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n295), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G190), .ZN(new_n316));
  INV_X1    g0116(.A(G200), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n316), .B(new_n268), .C1(new_n317), .C2(new_n315), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT8), .B(G58), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n321), .B(KEYINPUT67), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(new_n252), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT15), .B(G87), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n324), .A2(new_n254), .B1(new_n212), .B2(new_n222), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n250), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n222), .B1(new_n259), .B2(G20), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n266), .A2(new_n327), .B1(new_n222), .B2(new_n265), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n270), .A2(new_n271), .ZN(new_n330));
  INV_X1    g0130(.A(G1698), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n229), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n221), .A2(G1698), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n330), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT3), .B(G33), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n275), .B1(new_n335), .B2(G107), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n292), .B1(new_n223), .B2(new_n281), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n308), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n329), .A2(new_n341), .ZN(new_n342));
  OR2_X1    g0142(.A1(new_n342), .A2(KEYINPUT68), .ZN(new_n343));
  INV_X1    g0143(.A(G179), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n342), .A2(KEYINPUT68), .B1(new_n344), .B2(new_n339), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G150), .ZN(new_n347));
  OAI22_X1  g0147(.A1(new_n321), .A2(new_n254), .B1(new_n347), .B2(new_n252), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT66), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n348), .A2(new_n349), .B1(new_n203), .B2(G20), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n349), .B2(new_n348), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n250), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n226), .B1(new_n259), .B2(G20), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n266), .A2(new_n353), .B1(new_n226), .B2(new_n265), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n335), .A2(G222), .A3(new_n331), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n335), .A2(G223), .A3(G1698), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n356), .B(new_n357), .C1(new_n222), .C2(new_n335), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n275), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n282), .A2(G226), .B1(new_n285), .B2(new_n288), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n361), .A2(G179), .ZN(new_n362));
  AOI21_X1  g0162(.A(G169), .B1(new_n359), .B2(new_n360), .ZN(new_n363));
  OR3_X1    g0163(.A1(new_n355), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n329), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n339), .A2(G190), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n340), .A2(G200), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n346), .A2(new_n364), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n361), .A2(G200), .ZN(new_n371));
  INV_X1    g0171(.A(G190), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(new_n372), .B2(new_n361), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(KEYINPUT9), .B2(new_n355), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n355), .A2(KEYINPUT9), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT10), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT10), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n374), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n320), .A2(new_n370), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G58), .A2(G68), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n212), .B1(new_n214), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n251), .A2(G159), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT73), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n382), .ZN(new_n387));
  OAI21_X1  g0187(.A(G20), .B1(new_n387), .B2(new_n202), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT73), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(new_n384), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT72), .ZN(new_n392));
  OR2_X1    g0192(.A1(KEYINPUT3), .A2(G33), .ZN(new_n393));
  NAND2_X1  g0193(.A1(KEYINPUT3), .A2(G33), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(new_n212), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT7), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n393), .A2(KEYINPUT7), .A3(new_n212), .A4(new_n394), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n392), .B1(new_n399), .B2(G68), .ZN(new_n400));
  AOI211_X1 g0200(.A(KEYINPUT72), .B(new_n220), .C1(new_n397), .C2(new_n398), .ZN(new_n401));
  OAI211_X1 g0201(.A(KEYINPUT16), .B(new_n391), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  XOR2_X1   g0202(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n403));
  NAND2_X1  g0203(.A1(new_n386), .A2(new_n390), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n220), .B1(new_n397), .B2(new_n398), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n402), .A2(new_n406), .A3(new_n250), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n321), .B1(new_n259), .B2(G20), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(new_n266), .B1(new_n265), .B2(new_n321), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n292), .B1(new_n281), .B2(new_n229), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n227), .A2(G1698), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(G223), .B2(G1698), .ZN(new_n413));
  INV_X1    g0213(.A(G33), .ZN(new_n414));
  INV_X1    g0214(.A(G87), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n413), .A2(new_n330), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n411), .B1(new_n416), .B2(new_n275), .ZN(new_n417));
  OR2_X1    g0217(.A1(new_n417), .A2(new_n308), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(G179), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n410), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT18), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT18), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n410), .A2(new_n423), .A3(new_n420), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n372), .A2(KEYINPUT75), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n372), .A2(KEYINPUT75), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n417), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(G200), .B2(new_n417), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n407), .A2(new_n409), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT17), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n407), .A2(new_n430), .A3(KEYINPUT17), .A4(new_n409), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n422), .A2(new_n424), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n381), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g0236(.A(KEYINPUT5), .B(G41), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n287), .A2(G1), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n437), .A2(new_n438), .B1(new_n284), .B2(new_n278), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n259), .A2(G45), .ZN(new_n440));
  NOR2_X1   g0240(.A1(KEYINPUT5), .A2(G41), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(KEYINPUT5), .A2(G41), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n440), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n439), .A2(G270), .B1(new_n285), .B2(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(G264), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n446));
  OAI211_X1 g0246(.A(G257), .B(new_n331), .C1(new_n270), .C2(new_n271), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n393), .A2(G303), .A3(new_n394), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n275), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G116), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n265), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n250), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n259), .A2(G33), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n454), .A2(G116), .A3(new_n260), .A4(new_n455), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n249), .A2(new_n211), .B1(G20), .B2(new_n452), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G283), .ZN(new_n458));
  INV_X1    g0258(.A(G97), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n458), .B(new_n212), .C1(G33), .C2(new_n459), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n457), .A2(KEYINPUT20), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT20), .B1(new_n457), .B2(new_n460), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n453), .B(new_n456), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n451), .A2(G169), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT21), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n451), .A2(new_n463), .A3(KEYINPUT21), .A4(G169), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n445), .A2(G179), .A3(new_n450), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n463), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n463), .B1(new_n451), .B2(G200), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n428), .B2(new_n451), .ZN(new_n472));
  OAI211_X1 g0272(.A(G257), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n473));
  OAI211_X1 g0273(.A(G250), .B(new_n331), .C1(new_n270), .C2(new_n271), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G294), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n275), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n444), .A2(new_n285), .ZN(new_n478));
  INV_X1    g0278(.A(new_n443), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n438), .B1(new_n479), .B2(new_n441), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n480), .A2(G264), .A3(new_n279), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n477), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G169), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n439), .A2(KEYINPUT80), .A3(G264), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT80), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n476), .A2(new_n275), .B1(new_n285), .B2(new_n444), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n487), .A2(G179), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G107), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n491), .A2(KEYINPUT23), .A3(G20), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT23), .B1(new_n491), .B2(G20), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G116), .ZN(new_n494));
  OAI22_X1  g0294(.A1(new_n492), .A2(new_n493), .B1(G20), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT79), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT22), .ZN(new_n498));
  AOI21_X1  g0298(.A(G20), .B1(new_n393), .B2(new_n394), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n498), .B1(new_n499), .B2(G87), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n212), .B(G87), .C1(new_n270), .C2(new_n271), .ZN(new_n501));
  INV_X1    g0301(.A(new_n498), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n496), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT24), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n501), .A2(new_n502), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n335), .A2(new_n212), .A3(G87), .A4(new_n498), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT24), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n508), .A2(new_n509), .A3(new_n496), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n454), .B1(new_n505), .B2(new_n510), .ZN(new_n511));
  AND4_X1   g0311(.A1(new_n211), .A2(new_n260), .A3(new_n249), .A4(new_n455), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n265), .A2(KEYINPUT25), .A3(new_n491), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT25), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n260), .B2(G107), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n512), .A2(G107), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n490), .B1(new_n511), .B2(new_n517), .ZN(new_n518));
  AOI211_X1 g0318(.A(KEYINPUT24), .B(new_n495), .C1(new_n507), .C2(new_n506), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n509), .B1(new_n508), .B2(new_n496), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n250), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n482), .A2(G190), .ZN(new_n522));
  AOI21_X1  g0322(.A(G200), .B1(new_n487), .B2(new_n488), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n521), .B(new_n516), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n470), .A2(new_n472), .A3(new_n518), .A4(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n480), .A2(G257), .A3(new_n279), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n478), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(G250), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n393), .B2(new_n394), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT4), .ZN(new_n530));
  OAI21_X1  g0330(.A(G1698), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n458), .ZN(new_n532));
  OAI21_X1  g0332(.A(G244), .B1(new_n270), .B2(new_n271), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n532), .B1(new_n533), .B2(new_n530), .ZN(new_n534));
  AND2_X1   g0334(.A1(KEYINPUT4), .A2(G244), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n331), .B(new_n535), .C1(new_n270), .C2(new_n271), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n531), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n527), .B1(new_n537), .B2(new_n275), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G190), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT7), .B1(new_n330), .B2(new_n212), .ZN(new_n540));
  INV_X1    g0340(.A(new_n398), .ZN(new_n541));
  OAI21_X1  g0341(.A(G107), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT6), .ZN(new_n543));
  AND2_X1   g0343(.A1(G97), .A2(G107), .ZN(new_n544));
  NOR2_X1   g0344(.A1(G97), .A2(G107), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n491), .A2(KEYINPUT6), .A3(G97), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n548), .A2(G20), .B1(G77), .B2(new_n251), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n454), .B1(new_n542), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n260), .A2(G97), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n512), .B2(G97), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(G200), .B1(new_n538), .B2(KEYINPUT76), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n223), .B1(new_n393), .B2(new_n394), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n536), .B(new_n458), .C1(new_n556), .C2(KEYINPUT4), .ZN(new_n557));
  OAI21_X1  g0357(.A(G250), .B1(new_n270), .B2(new_n271), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n331), .B1(new_n558), .B2(KEYINPUT4), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n275), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n527), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT76), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n539), .B(new_n554), .C1(new_n555), .C2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n560), .A2(new_n561), .A3(G179), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n538), .B2(new_n308), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT77), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n550), .A2(new_n568), .A3(new_n553), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n491), .A2(KEYINPUT6), .A3(G97), .ZN(new_n570));
  XNOR2_X1  g0370(.A(G97), .B(G107), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n570), .B1(new_n571), .B2(new_n543), .ZN(new_n572));
  OAI22_X1  g0372(.A1(new_n572), .A2(new_n212), .B1(new_n222), .B2(new_n252), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n491), .B1(new_n397), .B2(new_n398), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n250), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT77), .B1(new_n575), .B2(new_n552), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n567), .B1(new_n569), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n221), .A2(G1698), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n270), .B2(new_n271), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT78), .ZN(new_n580));
  OAI211_X1 g0380(.A(G244), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT78), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n578), .B(new_n582), .C1(new_n271), .C2(new_n270), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n580), .A2(new_n494), .A3(new_n581), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n275), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n438), .A2(new_n283), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n440), .A2(new_n528), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n279), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(new_n344), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT19), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n212), .B1(new_n273), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n545), .A2(new_n415), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n212), .B(G68), .C1(new_n270), .C2(new_n271), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n590), .B1(new_n254), .B2(new_n459), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n250), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n324), .A2(new_n265), .ZN(new_n598));
  INV_X1    g0398(.A(new_n512), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n597), .B(new_n598), .C1(new_n324), .C2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n588), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n584), .B2(new_n275), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n589), .B(new_n600), .C1(G169), .C2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n585), .A2(G190), .A3(new_n588), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n512), .A2(G87), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n597), .A2(new_n598), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n604), .B(new_n607), .C1(new_n317), .C2(new_n602), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n565), .A2(new_n577), .A3(new_n603), .A4(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n525), .A2(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n436), .A2(new_n610), .ZN(G372));
  INV_X1    g0411(.A(new_n364), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT81), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n380), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT81), .B1(new_n377), .B2(new_n379), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n268), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n311), .B1(new_n310), .B2(new_n312), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n319), .B2(new_n346), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n622), .A2(new_n433), .A3(new_n434), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n422), .A2(new_n424), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n612), .B1(new_n617), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(G169), .B1(new_n585), .B2(new_n588), .ZN(new_n628));
  AOI211_X1 g0428(.A(G179), .B(new_n601), .C1(new_n584), .C2(new_n275), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n585), .A2(new_n588), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G200), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n606), .B1(new_n602), .B2(G190), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n630), .A2(new_n600), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n634), .A2(new_n565), .A3(new_n577), .A4(new_n524), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n521), .A2(new_n516), .B1(new_n483), .B2(new_n489), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n603), .A2(new_n608), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT26), .B1(new_n640), .B2(new_n577), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n562), .A2(G169), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n554), .B1(new_n642), .B2(new_n566), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n643), .A2(new_n644), .A3(new_n603), .A4(new_n608), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n641), .A2(new_n645), .A3(new_n603), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n639), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n436), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n627), .A2(new_n648), .ZN(G369));
  INV_X1    g0449(.A(G330), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n259), .A2(new_n212), .A3(G13), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT27), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n653), .A2(new_n259), .A3(new_n212), .A4(G13), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n652), .A2(G213), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT82), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(G343), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n636), .A2(new_n463), .A3(new_n658), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n464), .A2(new_n465), .B1(new_n468), .B2(new_n463), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n463), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n660), .A2(new_n472), .A3(new_n661), .A4(new_n467), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n650), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n658), .B1(new_n511), .B2(new_n517), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n518), .A2(new_n664), .A3(new_n524), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n637), .A2(new_n658), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n636), .A2(new_n518), .A3(new_n524), .A4(new_n657), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n637), .A2(new_n657), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n668), .A2(new_n671), .ZN(G399));
  INV_X1    g0472(.A(new_n208), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(G41), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n592), .A2(G116), .ZN(new_n676));
  XOR2_X1   g0476(.A(new_n676), .B(KEYINPUT83), .Z(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n675), .A2(new_n678), .A3(G1), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n215), .B2(new_n675), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT28), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT29), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT85), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n568), .B1(new_n550), .B2(new_n553), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n575), .A2(KEYINPUT77), .A3(new_n552), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n686), .A2(new_n603), .A3(new_n608), .A4(new_n567), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n603), .B1(new_n687), .B2(KEYINPUT26), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n644), .B1(new_n634), .B2(new_n643), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n683), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n575), .B(new_n552), .C1(new_n562), .C2(new_n372), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n538), .A2(KEYINPUT76), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n317), .B1(new_n562), .B2(new_n563), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n684), .A2(new_n685), .B1(new_n642), .B2(new_n566), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n694), .A2(new_n640), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT86), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n636), .B2(new_n637), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n470), .A2(KEYINPUT86), .A3(new_n518), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n696), .A2(new_n524), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n634), .A2(new_n644), .A3(new_n695), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n575), .A2(new_n552), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n567), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT26), .B1(new_n640), .B2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n701), .A2(new_n704), .A3(KEYINPUT85), .A4(new_n603), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n690), .A2(new_n700), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n682), .B1(new_n706), .B2(new_n657), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n682), .B(new_n657), .C1(new_n639), .C2(new_n646), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n487), .A2(new_n488), .ZN(new_n711));
  AOI21_X1  g0511(.A(G179), .B1(new_n445), .B2(new_n450), .ZN(new_n712));
  AND4_X1   g0512(.A1(new_n562), .A2(new_n631), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n484), .A2(new_n486), .B1(new_n275), .B2(new_n476), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n468), .A2(new_n538), .A3(new_n602), .A4(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT84), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n713), .B1(new_n717), .B2(KEYINPUT30), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n715), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n657), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n610), .A2(new_n657), .B1(new_n721), .B2(KEYINPUT31), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n718), .A2(new_n720), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n658), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G330), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n710), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n681), .B1(new_n730), .B2(G1), .ZN(G364));
  AND2_X1   g0531(.A1(new_n212), .A2(G13), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n259), .B1(new_n732), .B2(G45), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n675), .A2(KEYINPUT87), .A3(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT87), .ZN(new_n735));
  INV_X1    g0535(.A(new_n733), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n735), .B1(new_n674), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n208), .A2(new_n335), .ZN(new_n740));
  INV_X1    g0540(.A(G355), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n740), .A2(new_n741), .B1(G116), .B2(new_n208), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n673), .A2(new_n335), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(new_n287), .B2(new_n216), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n244), .A2(G45), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n742), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT88), .Z(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n211), .B1(G20), .B2(new_n308), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n739), .B1(new_n747), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n344), .A2(new_n317), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT91), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n756), .A2(new_n212), .A3(G190), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G159), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT32), .Z(new_n759));
  NOR2_X1   g0559(.A1(new_n212), .A2(G179), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(G190), .A3(G200), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n335), .B1(new_n761), .B2(new_n415), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT92), .Z(new_n763));
  NOR3_X1   g0563(.A1(new_n212), .A2(new_n344), .A3(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n427), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n760), .A2(new_n372), .A3(G200), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n765), .A2(new_n228), .B1(new_n491), .B2(new_n766), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n212), .A2(new_n344), .A3(new_n317), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n768), .A2(KEYINPUT90), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(KEYINPUT90), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n769), .A2(new_n427), .A3(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n767), .B1(G50), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n759), .A2(new_n763), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n764), .A2(new_n372), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n775), .A2(KEYINPUT89), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(KEYINPUT89), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AND3_X1   g0579(.A1(new_n769), .A2(new_n372), .A3(new_n770), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n779), .A2(G77), .B1(G68), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(G20), .B1(new_n756), .B2(new_n372), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n781), .B1(new_n459), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n765), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n335), .B1(new_n785), .B2(G322), .ZN(new_n786));
  INV_X1    g0586(.A(new_n761), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G303), .ZN(new_n788));
  INV_X1    g0588(.A(new_n775), .ZN(new_n789));
  INV_X1    g0589(.A(new_n766), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n789), .A2(G311), .B1(new_n790), .B2(G283), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n757), .A2(G329), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n786), .A2(new_n788), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n772), .A2(G326), .B1(G294), .B2(new_n782), .ZN(new_n794));
  INV_X1    g0594(.A(new_n780), .ZN(new_n795));
  XOR2_X1   g0595(.A(KEYINPUT33), .B(G317), .Z(new_n796));
  OAI21_X1  g0596(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n774), .A2(new_n784), .B1(new_n793), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n754), .B1(new_n798), .B2(new_n751), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n659), .A2(new_n662), .ZN(new_n800));
  INV_X1    g0600(.A(new_n750), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n663), .A2(new_n739), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(G330), .B2(new_n800), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  AND2_X1   g0606(.A1(new_n647), .A2(new_n657), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n365), .A2(new_n657), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(new_n343), .B2(new_n345), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n346), .A2(new_n368), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n810), .B1(new_n811), .B2(new_n809), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n807), .B(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n739), .B1(new_n813), .B2(new_n728), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(new_n728), .B2(new_n813), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n751), .A2(new_n748), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n738), .B1(new_n222), .B2(new_n816), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G97), .A2(new_n782), .B1(new_n785), .B2(G294), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT93), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G303), .A2(new_n772), .B1(new_n780), .B2(G283), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n330), .B1(new_n761), .B2(new_n491), .C1(new_n415), .C2(new_n766), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(G311), .B2(new_n757), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n820), .B(new_n822), .C1(new_n452), .C2(new_n778), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n780), .A2(G150), .B1(G143), .B2(new_n785), .ZN(new_n825));
  INV_X1    g0625(.A(G137), .ZN(new_n826));
  INV_X1    g0626(.A(G159), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n825), .B1(new_n826), .B2(new_n771), .C1(new_n827), .C2(new_n778), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT34), .Z(new_n829));
  OR2_X1    g0629(.A1(new_n829), .A2(KEYINPUT94), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n335), .B1(new_n766), .B2(new_n220), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(G50), .B2(new_n787), .ZN(new_n832));
  INV_X1    g0632(.A(G132), .ZN(new_n833));
  INV_X1    g0633(.A(new_n757), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n832), .B1(new_n783), .B2(new_n228), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(new_n829), .B2(KEYINPUT94), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n824), .B1(new_n830), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n751), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n817), .B1(new_n749), .B2(new_n812), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n815), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G384));
  OR2_X1    g0641(.A1(new_n548), .A2(KEYINPUT35), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n548), .A2(KEYINPUT35), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n842), .A2(new_n843), .A3(G116), .A4(new_n213), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT36), .Z(new_n845));
  NAND3_X1  g0645(.A1(new_n216), .A2(G77), .A3(new_n382), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n201), .A2(G68), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n259), .B(G13), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT38), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n410), .A2(new_n656), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n421), .A2(new_n851), .A3(new_n431), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT37), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT37), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n421), .A2(new_n851), .A3(new_n854), .A4(new_n431), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n853), .A2(KEYINPUT96), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n851), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n435), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT96), .B1(new_n853), .B2(new_n855), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n850), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT39), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n399), .A2(G68), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT72), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n405), .A2(new_n392), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n404), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n403), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n250), .B(new_n402), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n868), .A2(new_n409), .B1(new_n418), .B2(new_n419), .ZN(new_n869));
  INV_X1    g0669(.A(new_n656), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n868), .B2(new_n409), .ZN(new_n871));
  INV_X1    g0671(.A(new_n431), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n869), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n855), .B1(new_n873), .B2(new_n854), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n435), .A2(new_n871), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(new_n875), .A3(KEYINPUT38), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n861), .A2(new_n862), .A3(new_n876), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n874), .A2(new_n875), .A3(KEYINPUT38), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT38), .B1(new_n874), .B2(new_n875), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT39), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT97), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n314), .A2(new_n657), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT95), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT97), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n877), .A2(new_n885), .A3(new_n880), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n882), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n343), .A2(new_n345), .A3(new_n657), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n807), .B2(new_n812), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n618), .A2(new_n658), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n621), .A2(new_n318), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n306), .A2(new_n313), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n618), .B(new_n658), .C1(new_n893), .C2(new_n319), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n878), .A2(new_n879), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n896), .A2(new_n897), .B1(new_n624), .B2(new_n870), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n887), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n436), .B1(new_n707), .B2(new_n709), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n627), .A2(new_n900), .ZN(new_n901));
  XOR2_X1   g0701(.A(new_n899), .B(new_n901), .Z(new_n902));
  NAND2_X1  g0702(.A1(new_n861), .A2(new_n876), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n724), .A2(KEYINPUT98), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT98), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n721), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n904), .A2(new_n725), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n722), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n342), .A2(KEYINPUT68), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n329), .A2(KEYINPUT68), .A3(new_n341), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(G179), .B2(new_n340), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n808), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n368), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n343), .B2(new_n345), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n912), .B1(new_n914), .B2(new_n808), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n892), .B2(new_n894), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n903), .A2(KEYINPUT40), .A3(new_n908), .A4(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n908), .B(new_n916), .C1(new_n878), .C2(new_n879), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT99), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n919), .B1(new_n918), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n436), .A2(new_n908), .ZN(new_n924));
  OAI21_X1  g0724(.A(G330), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n924), .B2(new_n923), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n902), .A2(new_n926), .B1(new_n259), .B2(new_n732), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n902), .A2(new_n926), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n849), .B1(new_n927), .B2(new_n928), .ZN(G367));
  NOR2_X1   g0729(.A1(new_n744), .A2(new_n240), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n752), .B1(new_n208), .B2(new_n324), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n739), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n772), .A2(G143), .B1(G68), .B2(new_n782), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n933), .B1(new_n827), .B2(new_n795), .C1(new_n201), .C2(new_n778), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n765), .A2(new_n347), .B1(new_n228), .B2(new_n761), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n766), .A2(new_n222), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n935), .A2(new_n330), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n826), .B2(new_n834), .ZN(new_n938));
  AOI22_X1  g0738(.A1(G311), .A2(new_n772), .B1(new_n780), .B2(G294), .ZN(new_n939));
  INV_X1    g0739(.A(G283), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n939), .B1(new_n940), .B2(new_n778), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT46), .B1(new_n787), .B2(G116), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n757), .B2(G317), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n787), .A2(KEYINPUT46), .A3(G116), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n330), .B1(new_n766), .B2(new_n459), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n785), .B2(G303), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n782), .A2(G107), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n943), .A2(new_n944), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n934), .A2(new_n938), .B1(new_n941), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT47), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n932), .B1(new_n950), .B2(new_n751), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n657), .A2(new_n607), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(new_n603), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n634), .B2(new_n953), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n750), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n951), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n658), .A2(new_n702), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n565), .A2(new_n577), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n643), .A2(new_n658), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n669), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT100), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n966), .A2(KEYINPUT42), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n962), .A2(new_n637), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n658), .B1(new_n968), .B2(new_n577), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n966), .B2(KEYINPUT42), .ZN(new_n970));
  INV_X1    g0770(.A(new_n955), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n967), .A2(new_n970), .B1(KEYINPUT43), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(KEYINPUT43), .B2(new_n971), .ZN(new_n973));
  INV_X1    g0773(.A(new_n691), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n693), .A2(new_n692), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n974), .A2(new_n975), .B1(new_n686), .B2(new_n567), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n976), .A2(new_n959), .B1(new_n643), .B2(new_n658), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n668), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT43), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n967), .A2(new_n970), .A3(new_n979), .A4(new_n955), .ZN(new_n980));
  AND3_X1   g0780(.A1(new_n973), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n978), .B1(new_n973), .B2(new_n980), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n674), .B(KEYINPUT41), .Z(new_n984));
  NAND2_X1  g0784(.A1(new_n706), .A2(new_n657), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(KEYINPUT29), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n636), .A2(new_n657), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n665), .A2(new_n666), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n669), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n800), .A2(G330), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n986), .A2(new_n728), .A3(new_n708), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(KEYINPUT102), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT102), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n710), .A2(new_n995), .A3(new_n728), .A4(new_n992), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT44), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n671), .B2(new_n962), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n669), .A2(new_n670), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n977), .A2(KEYINPUT44), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT45), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n977), .B2(new_n999), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n671), .A2(KEYINPUT45), .A3(new_n962), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n668), .A2(KEYINPUT101), .ZN(new_n1006));
  AND3_X1   g0806(.A1(new_n1001), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1006), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n994), .A2(new_n996), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n984), .B1(new_n1011), .B2(new_n730), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n733), .B1(new_n1012), .B2(KEYINPUT103), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n650), .B1(new_n722), .B2(new_n726), .ZN(new_n1014));
  NOR4_X1   g0814(.A1(new_n707), .A2(new_n1014), .A3(new_n991), .A4(new_n709), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1009), .B1(new_n1015), .B2(new_n995), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n729), .B1(new_n1016), .B2(new_n994), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT103), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n1017), .A2(new_n1018), .A3(new_n984), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n983), .B1(new_n1013), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT104), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT104), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1022), .B(new_n983), .C1(new_n1013), .C2(new_n1019), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n958), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT105), .ZN(G387));
  NAND2_X1  g0825(.A1(new_n729), .A2(new_n991), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1026), .A2(new_n674), .A3(new_n993), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n765), .A2(new_n226), .B1(new_n222), .B2(new_n761), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n335), .B1(new_n459), .B2(new_n766), .C1(new_n834), .C2(new_n347), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(G68), .C2(new_n789), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n795), .A2(new_n321), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n783), .A2(new_n324), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n772), .A2(G159), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n757), .A2(G326), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n335), .B1(new_n790), .B2(G116), .ZN(new_n1036));
  INV_X1    g0836(.A(G294), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n783), .A2(new_n940), .B1(new_n1037), .B2(new_n761), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n780), .A2(G311), .B1(G317), .B2(new_n785), .ZN(new_n1039));
  INV_X1    g0839(.A(G303), .ZN(new_n1040));
  INV_X1    g0840(.A(G322), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1039), .B1(new_n1040), .B2(new_n778), .C1(new_n1041), .C2(new_n771), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT48), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1038), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n1043), .B2(new_n1042), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT49), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1035), .B(new_n1036), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1034), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n751), .ZN(new_n1050));
  AOI21_X1  g0850(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n322), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n226), .ZN(new_n1053));
  XOR2_X1   g0853(.A(KEYINPUT106), .B(KEYINPUT50), .Z(new_n1054));
  OAI211_X1 g0854(.A(new_n678), .B(new_n1051), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n743), .B1(new_n287), .B2(new_n237), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(G107), .B2(new_n208), .C1(new_n678), .C2(new_n740), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n738), .B1(new_n1058), .B2(new_n752), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1050), .B(new_n1059), .C1(new_n667), .C2(new_n801), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1027), .B(new_n1060), .C1(new_n733), .C2(new_n991), .ZN(G393));
  INV_X1    g0861(.A(KEYINPUT107), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1001), .A2(new_n1005), .B1(new_n1062), .B2(new_n668), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n668), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(KEYINPUT107), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1063), .B(new_n1065), .Z(new_n1066));
  AOI21_X1  g0866(.A(new_n675), .B1(new_n1066), .B2(new_n993), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1067), .A2(new_n1011), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n752), .B1(new_n459), .B2(new_n208), .C1(new_n744), .C2(new_n247), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n739), .A2(new_n1069), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n335), .B1(new_n761), .B2(new_n220), .C1(new_n415), .C2(new_n766), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n201), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n779), .A2(new_n1052), .B1(new_n1072), .B2(new_n780), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n222), .B2(new_n783), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1071), .B(new_n1074), .C1(G143), .C2(new_n757), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n771), .A2(new_n347), .B1(new_n765), .B2(new_n827), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT51), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n782), .A2(G116), .B1(G294), .B2(new_n789), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n795), .B2(new_n1040), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT109), .Z(new_n1080));
  AOI22_X1  g0880(.A1(new_n772), .A2(G317), .B1(new_n785), .B2(G311), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(KEYINPUT108), .B(KEYINPUT52), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n335), .B1(new_n790), .B2(G107), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n940), .B2(new_n761), .C1(new_n834), .C2(new_n1041), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1075), .A2(new_n1077), .B1(new_n1080), .B2(new_n1087), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1070), .B1(new_n801), .B2(new_n962), .C1(new_n1088), .C2(new_n838), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n1066), .B2(new_n733), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1068), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(G390));
  NAND3_X1  g0892(.A1(new_n812), .A2(new_n706), .A3(new_n657), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1093), .A2(new_n888), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n892), .A2(new_n894), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1014), .A2(new_n812), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n650), .B1(new_n907), .B2(new_n722), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1095), .B1(new_n1099), .B2(new_n812), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1014), .A2(new_n812), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n895), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1099), .A2(new_n916), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n890), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1098), .A2(new_n1101), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n436), .A2(new_n1099), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n627), .A2(new_n900), .A3(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT110), .Z(new_n1111));
  INV_X1    g0911(.A(new_n884), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n890), .B2(new_n895), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n877), .A2(new_n885), .A3(new_n880), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n885), .B1(new_n877), .B2(new_n880), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n903), .B(new_n1112), .C1(new_n1094), .C2(new_n895), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n1117), .A3(new_n1096), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1117), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n882), .A2(new_n886), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1119), .B1(new_n1120), .B2(new_n1113), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1118), .B1(new_n1121), .B2(new_n1104), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n675), .B1(new_n1111), .B2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1118), .B(new_n1110), .C1(new_n1121), .C2(new_n1104), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  OR2_X1    g0925(.A1(new_n1122), .A2(new_n733), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n749), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1120), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n738), .B1(new_n321), .B2(new_n816), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n780), .A2(G107), .B1(new_n782), .B2(G77), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1130), .B1(new_n459), .B2(new_n778), .C1(new_n940), .C2(new_n771), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n834), .A2(new_n1037), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n330), .B1(new_n761), .B2(new_n415), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n765), .A2(new_n452), .B1(new_n220), .B2(new_n766), .ZN(new_n1134));
  NOR4_X1   g0934(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  OR2_X1    g0936(.A1(new_n1136), .A2(KEYINPUT111), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n335), .B1(new_n201), .B2(new_n766), .C1(new_n765), .C2(new_n833), .ZN(new_n1138));
  OR3_X1    g0938(.A1(new_n761), .A2(KEYINPUT53), .A3(new_n347), .ZN(new_n1139));
  OAI21_X1  g0939(.A(KEYINPUT53), .B1(new_n761), .B2(new_n347), .ZN(new_n1140));
  INV_X1    g0940(.A(G125), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1139), .B(new_n1140), .C1(new_n834), .C2(new_n1141), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1138), .B(new_n1142), .C1(G137), .C2(new_n780), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n772), .A2(G128), .B1(G159), .B2(new_n782), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(KEYINPUT54), .B(G143), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1143), .B(new_n1144), .C1(new_n778), .C2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1136), .A2(KEYINPUT111), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1137), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1128), .B(new_n1129), .C1(new_n838), .C2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1125), .A2(new_n1126), .A3(new_n1149), .ZN(G378));
  OAI211_X1 g0950(.A(G330), .B(new_n917), .C1(new_n921), .C2(new_n922), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n899), .A2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n355), .A2(new_n870), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT55), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n617), .A2(new_n364), .A3(new_n1156), .ZN(new_n1157));
  XOR2_X1   g0957(.A(KEYINPUT113), .B(KEYINPUT56), .Z(new_n1158));
  OAI21_X1  g0958(.A(new_n1155), .B1(new_n616), .B2(new_n612), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1158), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1151), .A2(new_n887), .A3(new_n898), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1153), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1162), .B1(new_n1153), .B2(new_n1163), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1127), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n816), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n739), .B1(new_n1072), .B2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT112), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n783), .A2(new_n347), .B1(new_n771), .B2(new_n1141), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n785), .A2(G128), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1172), .B1(new_n826), .B2(new_n775), .C1(new_n761), .C2(new_n1145), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(G132), .C2(new_n780), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n414), .B(new_n286), .C1(new_n766), .C2(new_n827), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n757), .B2(G124), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n780), .A2(G97), .B1(new_n782), .B2(G68), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n452), .B2(new_n771), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n335), .A2(G41), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(new_n222), .B2(new_n761), .C1(new_n834), .C2(new_n940), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n785), .A2(G107), .B1(G58), .B2(new_n790), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n324), .B2(new_n775), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1182), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1187), .A2(KEYINPUT58), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(KEYINPUT58), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1183), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1190), .B(new_n226), .C1(G33), .C2(G41), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1180), .A2(new_n1188), .A3(new_n1189), .A4(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1170), .B1(new_n1192), .B2(new_n751), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1166), .A2(new_n736), .B1(new_n1167), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT114), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n627), .A2(new_n900), .A3(new_n1108), .ZN(new_n1196));
  AND3_X1   g0996(.A1(new_n1124), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1195), .B1(new_n1124), .B2(new_n1196), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1166), .B(KEYINPUT57), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n674), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1124), .A2(new_n1196), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(KEYINPUT114), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1124), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(KEYINPUT57), .B1(new_n1204), .B2(new_n1166), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1194), .B1(new_n1200), .B2(new_n1205), .ZN(G375));
  INV_X1    g1006(.A(new_n984), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1102), .A2(new_n895), .B1(new_n1099), .B2(new_n916), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n1097), .A2(new_n1100), .B1(new_n1208), .B2(new_n890), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1111), .B(new_n1207), .C1(new_n1196), .C2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n895), .A2(new_n748), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n739), .B1(G68), .B2(new_n1168), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n771), .A2(new_n833), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT117), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n765), .A2(new_n826), .B1(new_n827), .B2(new_n761), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G150), .B2(new_n789), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n335), .B1(new_n766), .B2(new_n228), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n757), .B2(G128), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1145), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n780), .A2(new_n1219), .B1(new_n782), .B2(G50), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1214), .A2(new_n1216), .A3(new_n1218), .A4(new_n1220), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n779), .A2(G107), .B1(G116), .B2(new_n780), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n1037), .B2(new_n771), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT115), .Z(new_n1224));
  AOI22_X1  g1024(.A1(new_n757), .A2(G303), .B1(G97), .B2(new_n787), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT116), .Z(new_n1226));
  AOI211_X1 g1026(.A(new_n335), .B(new_n936), .C1(new_n785), .C2(G283), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1226), .A2(new_n1032), .A3(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1221), .B1(new_n1224), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1212), .B1(new_n1229), .B2(new_n751), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1209), .A2(new_n736), .B1(new_n1211), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1210), .A2(new_n1231), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT118), .Z(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(G381));
  NAND2_X1  g1034(.A1(new_n1126), .A2(new_n1149), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n1124), .B2(new_n1123), .ZN(new_n1236));
  NOR4_X1   g1036(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1233), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  OR3_X1    g1038(.A1(new_n1238), .A2(G387), .A3(G375), .ZN(G407));
  INV_X1    g1039(.A(G343), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(G213), .ZN(new_n1241));
  OR3_X1    g1041(.A1(G375), .A2(G378), .A3(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(G407), .A2(G213), .A3(new_n1242), .ZN(G409));
  INV_X1    g1043(.A(KEYINPUT126), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(G393), .B(new_n805), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT122), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n1024), .B2(G390), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  XOR2_X1   g1048(.A(new_n1091), .B(KEYINPUT125), .Z(new_n1249));
  AOI21_X1  g1049(.A(new_n1248), .B1(G387), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT123), .B1(new_n1024), .B2(G390), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1023), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1018), .B1(new_n1017), .B2(new_n984), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1011), .A2(new_n730), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1254), .A2(KEYINPUT103), .A3(new_n1207), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(new_n733), .A3(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1022), .B1(new_n1256), .B2(new_n983), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n957), .B1(new_n1252), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT123), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n1259), .A3(new_n1091), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1024), .A2(G390), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1251), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1246), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(KEYINPUT124), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT124), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1262), .A2(new_n1265), .A3(new_n1246), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1250), .B1(new_n1264), .B2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1244), .B1(new_n1267), .B2(KEYINPUT61), .ZN(new_n1268));
  OAI211_X1 g1068(.A(G378), .B(new_n1194), .C1(new_n1200), .C2(new_n1205), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1204), .A2(new_n1207), .A3(new_n1166), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1194), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1236), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1269), .A2(new_n1272), .B1(G213), .B2(new_n1240), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1101), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1274), .A2(new_n1275), .A3(new_n1109), .A4(KEYINPUT60), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(KEYINPUT119), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT119), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1107), .A2(new_n1278), .A3(KEYINPUT60), .A4(new_n1109), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT60), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1209), .B2(new_n1196), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n675), .B1(new_n1209), .B2(new_n1196), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1280), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G384), .B1(new_n1285), .B2(new_n1231), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1231), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n840), .B(new_n1287), .C1(new_n1280), .C2(new_n1284), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1273), .A2(KEYINPUT63), .A3(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1273), .A2(new_n1289), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1240), .A2(G213), .A3(G2897), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT120), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1292), .B1(new_n1289), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT121), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(new_n1279), .B2(new_n1277), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n840), .B1(new_n1297), .B2(new_n1287), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1285), .A2(G384), .A3(new_n1231), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1295), .B1(new_n1300), .B2(KEYINPUT120), .ZN(new_n1301));
  AOI211_X1 g1101(.A(new_n1293), .B(KEYINPUT121), .C1(new_n1298), .C2(new_n1299), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1294), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(KEYINPUT121), .B1(new_n1289), .B2(new_n1293), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1292), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1305), .B1(new_n1300), .B2(KEYINPUT120), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1300), .A2(KEYINPUT120), .A3(new_n1295), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1304), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1303), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1269), .A2(new_n1272), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1309), .B1(new_n1310), .B2(new_n1241), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT63), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1291), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(G387), .A2(new_n1249), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1247), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1262), .A2(new_n1265), .A3(new_n1246), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1265), .B1(new_n1262), .B2(new_n1246), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1315), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT61), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1318), .A2(KEYINPUT126), .A3(new_n1319), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1268), .A2(new_n1290), .A3(new_n1313), .A4(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT62), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1310), .A2(new_n1322), .A3(new_n1241), .A4(new_n1289), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1323), .B(new_n1319), .C1(new_n1273), .C2(new_n1309), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1322), .B1(new_n1273), .B2(new_n1289), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1267), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1321), .A2(new_n1326), .ZN(G405));
  NAND2_X1  g1127(.A1(G375), .A2(new_n1236), .ZN(new_n1328));
  OR2_X1    g1128(.A1(new_n1300), .A2(KEYINPUT127), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1328), .A2(new_n1269), .A3(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1329), .B1(new_n1328), .B2(new_n1269), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(new_n1332), .B(new_n1318), .ZN(G402));
endmodule


