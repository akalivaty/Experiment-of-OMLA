//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n585, new_n586, new_n587, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1262,
    new_n1263, new_n1264, new_n1265;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G108), .Z(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT67), .ZN(G234));
  NAND2_X1  g027(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT68), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n461), .A2(KEYINPUT69), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n457), .A2(G567), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(KEYINPUT69), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT70), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n470), .A2(new_n467), .A3(G101), .A4(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  OAI211_X1 g049(.A(G137), .B(new_n467), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g051(.A(G125), .B1(new_n473), .B2(new_n474), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n467), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n476), .A2(new_n479), .ZN(G160));
  OR2_X1    g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n473), .A2(new_n474), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT71), .ZN(new_n487));
  AOI21_X1  g062(.A(G2105), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n467), .B1(new_n485), .B2(new_n487), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  OR2_X1    g066(.A1(G100), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n489), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  NAND2_X1  g070(.A1(G126), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT73), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n467), .A2(G138), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n496), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(new_n483), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n503), .B1(new_n473), .B2(new_n474), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(new_n498), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT72), .A2(G114), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT72), .A2(G114), .ZN(new_n507));
  OAI21_X1  g082(.A(G2105), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g083(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n501), .A2(new_n505), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G62), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n514), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  OAI211_X1 g097(.A(G50), .B(G543), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  AND2_X1   g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n524), .A2(new_n525), .B1(new_n521), .B2(new_n522), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT74), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT6), .B(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n517), .A2(new_n531), .A3(G88), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n532), .A2(KEYINPUT74), .A3(new_n523), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n520), .B1(new_n530), .B2(new_n533), .ZN(G166));
  INV_X1    g109(.A(new_n517), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n531), .A2(G89), .ZN(new_n536));
  NAND2_X1  g111(.A1(G63), .A2(G651), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n531), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G51), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n538), .A2(new_n543), .ZN(G168));
  AOI22_X1  g119(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n514), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT75), .B(G90), .Z(new_n548));
  OAI22_X1  g123(.A1(new_n541), .A2(new_n547), .B1(new_n526), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(G171));
  AOI22_X1  g125(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n514), .ZN(new_n552));
  INV_X1    g127(.A(G43), .ZN(new_n553));
  XNOR2_X1  g128(.A(KEYINPUT76), .B(G81), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n541), .A2(new_n553), .B1(new_n526), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n558));
  XOR2_X1   g133(.A(new_n558), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT79), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n563), .B(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(new_n515), .B2(new_n516), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  OR2_X1    g143(.A1(KEYINPUT6), .A2(G651), .ZN(new_n569));
  NAND2_X1  g144(.A1(KEYINPUT6), .A2(G651), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n515), .A2(new_n516), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G91), .ZN(new_n572));
  AND2_X1   g147(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(G543), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n569), .B2(new_n570), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n575), .A2(new_n576), .A3(G53), .ZN(new_n577));
  OAI211_X1 g152(.A(G53), .B(G543), .C1(new_n521), .C2(new_n522), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT9), .ZN(new_n579));
  AND3_X1   g154(.A1(new_n577), .A2(KEYINPUT78), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(KEYINPUT78), .B1(new_n577), .B2(new_n579), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n573), .B1(new_n580), .B2(new_n581), .ZN(G299));
  INV_X1    g157(.A(G171), .ZN(G301));
  XNOR2_X1  g158(.A(G168), .B(KEYINPUT80), .ZN(G286));
  INV_X1    g159(.A(new_n520), .ZN(new_n585));
  AND3_X1   g160(.A1(new_n532), .A2(KEYINPUT74), .A3(new_n523), .ZN(new_n586));
  AOI21_X1  g161(.A(KEYINPUT74), .B1(new_n532), .B2(new_n523), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(G303));
  INV_X1    g163(.A(G74), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n515), .A2(new_n589), .A3(new_n516), .ZN(new_n590));
  AOI22_X1  g165(.A1(G49), .A2(new_n575), .B1(new_n590), .B2(G651), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT81), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n571), .B2(G87), .ZN(new_n593));
  INV_X1    g168(.A(G87), .ZN(new_n594));
  NOR3_X1   g169(.A1(new_n526), .A2(KEYINPUT81), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n591), .B1(new_n593), .B2(new_n595), .ZN(G288));
  AOI22_X1  g171(.A1(new_n571), .A2(G86), .B1(new_n575), .B2(G48), .ZN(new_n597));
  OAI21_X1  g172(.A(G61), .B1(new_n525), .B2(new_n524), .ZN(new_n598));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n514), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n597), .A2(new_n601), .ZN(G305));
  AOI22_X1  g177(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(new_n514), .ZN(new_n604));
  INV_X1    g179(.A(G47), .ZN(new_n605));
  INV_X1    g180(.A(G85), .ZN(new_n606));
  OAI22_X1  g181(.A1(new_n541), .A2(new_n605), .B1(new_n526), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  AND3_X1   g185(.A1(new_n517), .A2(new_n531), .A3(G92), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g187(.A1(G79), .A2(G543), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT82), .ZN(new_n614));
  INV_X1    g189(.A(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n535), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n616), .A2(G651), .B1(G54), .B2(new_n575), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n610), .B1(new_n619), .B2(G868), .ZN(G284));
  OAI21_X1  g195(.A(new_n610), .B1(new_n619), .B2(G868), .ZN(G321));
  MUX2_X1   g196(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g197(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n619), .B1(new_n624), .B2(G860), .ZN(G148));
  INV_X1    g200(.A(new_n556), .ZN(new_n626));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n618), .A2(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(new_n627), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT83), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G111), .ZN(new_n635));
  AOI22_X1  g210(.A1(new_n632), .A2(new_n633), .B1(new_n635), .B2(G2105), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n490), .A2(G123), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n488), .A2(G135), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND3_X1  g215(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT12), .Z(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT13), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n644), .ZN(G156));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n649), .B2(new_n648), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n651), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(G14), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n660), .B1(new_n659), .B2(new_n657), .ZN(G401));
  XOR2_X1   g236(.A(G2067), .B(G2678), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT84), .ZN(new_n663));
  NOR2_X1   g238(.A1(G2072), .A2(G2078), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n442), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n663), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT18), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n663), .A2(new_n665), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n665), .B(KEYINPUT17), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n670), .B(new_n667), .C1(new_n663), .C2(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n663), .A2(new_n666), .A3(new_n671), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2096), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(KEYINPUT85), .B(KEYINPUT19), .Z(new_n677));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1956), .B(G2474), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT20), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n679), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n679), .B2(new_n685), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G229));
  NAND2_X1  g269(.A1(new_n490), .A2(G129), .ZN(new_n695));
  NAND3_X1  g270(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT26), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n467), .A2(G2104), .ZN(new_n700));
  AOI22_X1  g275(.A1(new_n698), .A2(new_n699), .B1(G105), .B2(new_n700), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n488), .A2(G141), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n704), .A2(KEYINPUT94), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT94), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n702), .B2(new_n703), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G29), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G29), .B2(G32), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT27), .B(G1996), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G21), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G168), .B2(new_n713), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(G1966), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT96), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G33), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT25), .Z(new_n721));
  AOI22_X1  g296(.A1(new_n483), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n467), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n488), .B2(G139), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n719), .B1(new_n724), .B2(new_n718), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G2072), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n713), .A2(G4), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n619), .B2(new_n713), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G1348), .ZN(new_n729));
  NOR4_X1   g304(.A1(new_n712), .A2(new_n717), .A3(new_n726), .A4(new_n729), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT97), .B(KEYINPUT23), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n713), .A2(G20), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n568), .A2(new_n572), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n577), .A2(new_n579), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT78), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n577), .A2(new_n579), .A3(KEYINPUT78), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n734), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n733), .B1(new_n739), .B2(new_n713), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1956), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n710), .B2(new_n711), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n718), .A2(G35), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G162), .B2(new_n718), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT29), .ZN(new_n745));
  INV_X1    g320(.A(G2090), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G34), .ZN(new_n748));
  AOI21_X1  g323(.A(G29), .B1(new_n748), .B2(KEYINPUT24), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(KEYINPUT24), .B2(new_n748), .ZN(new_n750));
  INV_X1    g325(.A(G160), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(new_n718), .ZN(new_n752));
  INV_X1    g327(.A(G2084), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n755), .A2(KEYINPUT93), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(KEYINPUT93), .ZN(new_n757));
  NOR2_X1   g332(.A1(G5), .A2(G16), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G171), .B2(G16), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G1961), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT31), .B(G11), .Z(new_n761));
  INV_X1    g336(.A(KEYINPUT30), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n718), .B1(new_n762), .B2(G28), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(KEYINPUT95), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n762), .B2(G28), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(KEYINPUT95), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n761), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n756), .A2(new_n757), .A3(new_n760), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n718), .A2(G26), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT28), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n488), .A2(G140), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n490), .A2(G128), .ZN(new_n772));
  OR2_X1    g347(.A1(G104), .A2(G2105), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n773), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n771), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n770), .B1(new_n775), .B2(G29), .ZN(new_n776));
  INV_X1    g351(.A(G2067), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n718), .A2(G27), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G164), .B2(new_n718), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(G2078), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n556), .A2(G16), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G16), .B2(G19), .ZN(new_n783));
  INV_X1    g358(.A(G1341), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n781), .B(new_n785), .C1(new_n718), .C2(new_n639), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n753), .A2(new_n752), .B1(new_n715), .B2(G1966), .ZN(new_n787));
  OAI221_X1 g362(.A(new_n787), .B1(G1961), .B2(new_n759), .C1(new_n784), .C2(new_n783), .ZN(new_n788));
  NOR4_X1   g363(.A1(new_n768), .A2(new_n778), .A3(new_n786), .A4(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n730), .A2(new_n742), .A3(new_n747), .A4(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G48), .ZN(new_n791));
  INV_X1    g366(.A(G86), .ZN(new_n792));
  OAI22_X1  g367(.A1(new_n541), .A2(new_n791), .B1(new_n526), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(new_n600), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(G16), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G6), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT32), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(G1981), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n796), .A2(KEYINPUT32), .ZN(new_n799));
  INV_X1    g374(.A(G1981), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n796), .A2(KEYINPUT32), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n713), .A2(G22), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G166), .B2(new_n713), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT90), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(G1971), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(G1971), .ZN(new_n808));
  NOR2_X1   g383(.A1(G16), .A2(G23), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT89), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G288), .B2(new_n713), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT33), .B(G1976), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n803), .A2(new_n807), .A3(new_n808), .A4(new_n813), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT88), .B(KEYINPUT34), .Z(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n718), .A2(G25), .ZN(new_n818));
  OAI21_X1  g393(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n819));
  INV_X1    g394(.A(G107), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(G2105), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n488), .B2(G131), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n490), .A2(KEYINPUT86), .A3(G119), .ZN(new_n823));
  AOI21_X1  g398(.A(KEYINPUT86), .B1(new_n490), .B2(G119), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n818), .B1(new_n825), .B2(G29), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT35), .B(G1991), .Z(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n826), .A2(new_n828), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT87), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n829), .B2(new_n830), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n713), .A2(G24), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n608), .B2(new_n713), .ZN(new_n835));
  INV_X1    g410(.A(G1986), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  NOR3_X1   g413(.A1(new_n817), .A2(new_n832), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n814), .A2(new_n816), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n840), .A2(KEYINPUT91), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(KEYINPUT91), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT92), .B(KEYINPUT36), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n839), .B(new_n844), .C1(new_n841), .C2(new_n842), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n790), .B1(new_n846), .B2(new_n847), .ZN(G311));
  INV_X1    g423(.A(new_n790), .ZN(new_n849));
  INV_X1    g424(.A(new_n847), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n840), .B(KEYINPUT91), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n844), .B1(new_n851), .B2(new_n839), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n849), .B1(new_n850), .B2(new_n852), .ZN(G150));
  INV_X1    g428(.A(G55), .ZN(new_n854));
  XOR2_X1   g429(.A(KEYINPUT98), .B(G93), .Z(new_n855));
  OAI22_X1  g430(.A1(new_n541), .A2(new_n854), .B1(new_n526), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(KEYINPUT99), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n575), .A2(G55), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n858), .B(new_n859), .C1(new_n526), .C2(new_n855), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n862), .A2(new_n514), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n863), .B1(new_n857), .B2(new_n860), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT100), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n867), .A2(new_n626), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(KEYINPUT100), .A3(new_n556), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT38), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n619), .A2(G559), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT39), .ZN(new_n876));
  AOI21_X1  g451(.A(G860), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n876), .B2(new_n875), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n865), .A2(G860), .ZN(new_n879));
  XOR2_X1   g454(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n878), .A2(new_n881), .ZN(G145));
  OR2_X1    g457(.A1(new_n775), .A2(G164), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n775), .A2(G164), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n488), .A2(G142), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n490), .A2(G130), .ZN(new_n887));
  OR2_X1    g462(.A1(G106), .A2(G2105), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n888), .B(G2104), .C1(G118), .C2(new_n467), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n885), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n825), .A2(new_n642), .ZN(new_n893));
  INV_X1    g468(.A(new_n825), .ZN(new_n894));
  INV_X1    g469(.A(new_n642), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n883), .A2(new_n884), .A3(new_n890), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n892), .A2(new_n893), .A3(new_n896), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n893), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n883), .A2(new_n884), .A3(new_n890), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n890), .B1(new_n883), .B2(new_n884), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n724), .B1(new_n705), .B2(new_n707), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n704), .A2(new_n724), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n639), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n639), .A2(new_n909), .ZN(new_n912));
  OAI21_X1  g487(.A(G160), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n912), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(new_n751), .A3(new_n910), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n913), .A2(new_n915), .A3(G162), .ZN(new_n916));
  AOI21_X1  g491(.A(G162), .B1(new_n913), .B2(new_n915), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n898), .A2(new_n902), .A3(new_n906), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n908), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n908), .A2(new_n918), .A3(KEYINPUT103), .A4(new_n919), .ZN(new_n923));
  AOI21_X1  g498(.A(G37), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n918), .ZN(new_n925));
  INV_X1    g500(.A(new_n919), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n906), .B1(new_n898), .B2(new_n902), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT104), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n925), .B(new_n930), .C1(new_n926), .C2(new_n927), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n924), .A2(new_n932), .A3(KEYINPUT40), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT40), .B1(new_n924), .B2(new_n932), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(G395));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n618), .A2(G299), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n618), .A2(G299), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n870), .A2(new_n629), .A3(new_n871), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n629), .B1(new_n870), .B2(new_n871), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT42), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT41), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n938), .A2(new_n946), .A3(new_n939), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n618), .A2(G299), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT41), .B1(new_n948), .B2(new_n937), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n629), .ZN(new_n951));
  INV_X1    g526(.A(new_n869), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n626), .B1(new_n868), .B2(KEYINPUT100), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n871), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n951), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n870), .A2(new_n629), .A3(new_n871), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n950), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n944), .A2(new_n945), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n945), .B1(new_n944), .B2(new_n958), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n794), .A2(KEYINPUT105), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n794), .A2(KEYINPUT105), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n963), .A3(G288), .ZN(new_n964));
  XNOR2_X1  g539(.A(G166), .B(new_n608), .ZN(new_n965));
  INV_X1    g540(.A(G288), .ZN(new_n966));
  INV_X1    g541(.A(new_n961), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n966), .B1(new_n962), .B2(new_n967), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n964), .A2(new_n965), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n965), .B1(new_n964), .B2(new_n968), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n959), .A2(new_n960), .A3(new_n972), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n950), .A2(new_n956), .A3(new_n957), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n940), .B1(new_n956), .B2(new_n957), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT42), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n944), .A2(new_n958), .A3(new_n945), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n971), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(G868), .B1(new_n973), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n868), .A2(G868), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n936), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n972), .B1(new_n959), .B2(new_n960), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n976), .A2(new_n971), .A3(new_n977), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n627), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n985), .A2(KEYINPUT106), .A3(new_n980), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n982), .A2(new_n986), .ZN(G295));
  NAND2_X1  g562(.A1(new_n979), .A2(new_n981), .ZN(G331));
  NOR2_X1   g563(.A1(G171), .A2(G168), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(G286), .B2(G301), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n991), .A2(new_n870), .A3(new_n871), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n991), .B1(new_n871), .B2(new_n870), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n941), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n991), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n872), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n997), .A2(new_n950), .A3(new_n992), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n995), .A2(new_n971), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G37), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n971), .B1(new_n995), .B2(new_n998), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT43), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n947), .A2(new_n949), .A3(KEYINPUT107), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT107), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n940), .A2(new_n1005), .A3(KEYINPUT41), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1004), .A2(new_n997), .A3(new_n992), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n995), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n972), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1009), .A2(new_n1010), .A3(new_n1000), .A4(new_n999), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n1003), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1002), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1014), .A2(new_n1010), .A3(new_n1000), .A4(new_n999), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT108), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1001), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT108), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1017), .A2(new_n1018), .A3(new_n1010), .A4(new_n1014), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1009), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT43), .B1(new_n1020), .B2(new_n1001), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1016), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1013), .B1(new_n1022), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g598(.A(G1384), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n512), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G40), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n476), .A2(new_n479), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1025), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1996), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n708), .A2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n775), .B(new_n777), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1029), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n704), .A2(new_n1034), .A3(G1996), .ZN(new_n1035));
  XOR2_X1   g610(.A(new_n1035), .B(KEYINPUT110), .Z(new_n1036));
  NOR2_X1   g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n894), .A2(new_n827), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n894), .A2(new_n827), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1034), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1037), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n608), .A2(new_n836), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1043), .B(KEYINPUT109), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n836), .B2(new_n608), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1042), .B1(new_n1034), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n483), .A2(new_n500), .B1(new_n504), .B2(new_n498), .ZN(new_n1049));
  AOI21_X1  g624(.A(G1384), .B1(new_n1049), .B2(new_n511), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1027), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n512), .A2(new_n1051), .A3(new_n1024), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1048), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1961), .ZN(new_n1055));
  INV_X1    g630(.A(G125), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1056), .B1(new_n481), .B2(new_n482), .ZN(new_n1057));
  INV_X1    g632(.A(new_n478), .ZN(new_n1058));
  OAI21_X1  g633(.A(G2105), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1059), .A2(G40), .A3(new_n472), .A4(new_n475), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1060), .B1(new_n1025), .B2(KEYINPUT50), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(KEYINPUT121), .A3(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1054), .A2(new_n1055), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT123), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1060), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n512), .A2(KEYINPUT45), .A3(new_n1024), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT116), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n512), .A2(new_n1069), .A3(KEYINPUT45), .A4(new_n1024), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(G2078), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1066), .A2(new_n1068), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1064), .A2(new_n1065), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1075), .A2(new_n1027), .A3(new_n1067), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1071), .B1(new_n1077), .B2(G2078), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1074), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1065), .B1(new_n1064), .B2(new_n1073), .ZN(new_n1080));
  OAI21_X1  g655(.A(G171), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1076), .A2(new_n1072), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT124), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n1082), .B(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1084), .A2(G301), .A3(new_n1064), .A4(new_n1078), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT54), .B1(new_n1081), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1976), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT114), .B1(G288), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT52), .B1(G288), .B2(new_n1087), .ZN(new_n1089));
  INV_X1    g664(.A(G8), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n1050), .B2(new_n1027), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n571), .A2(new_n592), .A3(G87), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT81), .B1(new_n526), .B2(new_n594), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1094), .A2(new_n1095), .A3(G1976), .A4(new_n591), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1088), .A2(new_n1089), .A3(new_n1091), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT49), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n793), .A2(G1981), .A3(new_n600), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n800), .B1(new_n597), .B2(new_n601), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(G1981), .B1(new_n793), .B2(new_n600), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n597), .A2(new_n601), .A3(new_n800), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n1103), .A3(KEYINPUT49), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1101), .A2(new_n1091), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1097), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1088), .A2(new_n1091), .A3(new_n1096), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1107), .A2(KEYINPUT115), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT52), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(new_n1107), .B2(KEYINPUT115), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1106), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1052), .A2(G2090), .A3(new_n1053), .ZN(new_n1112));
  AOI21_X1  g687(.A(G1971), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1113));
  OAI21_X1  g688(.A(G8), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n1115));
  NOR3_X1   g690(.A1(G166), .A2(new_n1090), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT55), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1117), .A2(KEYINPUT112), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1118), .B1(G303), .B2(G8), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1114), .A2(new_n1120), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1111), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT113), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1115), .ZN(new_n1125));
  NAND3_X1  g700(.A1(G303), .A2(G8), .A3(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(G166), .A2(new_n1090), .ZN(new_n1127));
  OAI211_X1 g702(.A(KEYINPUT113), .B(new_n1126), .C1(new_n1127), .C2(new_n1118), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT111), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1061), .A2(new_n746), .A3(new_n1062), .ZN(new_n1132));
  OAI211_X1 g707(.A(KEYINPUT111), .B(new_n1132), .C1(new_n1076), .C2(G1971), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1129), .A2(new_n1131), .A3(G8), .A4(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT51), .ZN(new_n1135));
  INV_X1    g710(.A(G1966), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1066), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1051), .B1(new_n512), .B2(new_n1024), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1053), .A2(new_n1138), .A3(new_n1060), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1136), .A2(new_n1137), .B1(new_n1139), .B2(new_n753), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1090), .B1(new_n1140), .B2(G168), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1137), .A2(new_n1136), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1139), .A2(new_n753), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(G168), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1135), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1147));
  AOI211_X1 g722(.A(KEYINPUT51), .B(new_n1090), .C1(new_n1140), .C2(G168), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1122), .B(new_n1134), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1086), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1064), .A2(new_n1073), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT123), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1152), .A2(G301), .A3(new_n1078), .A4(new_n1074), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT125), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1074), .A2(new_n1078), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1155), .A2(new_n1156), .A3(G301), .A4(new_n1152), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1084), .A2(new_n1064), .A3(new_n1078), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1159), .B1(new_n1160), .B2(G171), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT57), .ZN(new_n1163));
  AND4_X1   g738(.A1(new_n1163), .A2(new_n735), .A3(new_n572), .A4(new_n568), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(new_n739), .B2(new_n1163), .ZN(new_n1166));
  XNOR2_X1  g741(.A(KEYINPUT56), .B(G2072), .ZN(new_n1167));
  AND4_X1   g742(.A1(new_n1027), .A2(new_n1075), .A3(new_n1067), .A4(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(G1956), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1166), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(KEYINPUT119), .B1(new_n1025), .B2(new_n1060), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT119), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1050), .A2(new_n1027), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n777), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(KEYINPUT120), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT120), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1175), .A2(new_n1178), .A3(new_n777), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(G1348), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1054), .A2(new_n1181), .A3(new_n1063), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1164), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1066), .A2(new_n1067), .A3(new_n1167), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1184), .B(new_n1185), .C1(new_n1139), .C2(G1956), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1186), .A2(new_n619), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1171), .B1(new_n1183), .B2(new_n1187), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1170), .A2(new_n1186), .A3(KEYINPUT61), .ZN(new_n1189));
  AOI21_X1  g764(.A(KEYINPUT61), .B1(new_n1170), .B2(new_n1186), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1180), .A2(KEYINPUT60), .A3(new_n618), .A4(new_n1182), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT59), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT122), .ZN(new_n1194));
  XOR2_X1   g769(.A(KEYINPUT58), .B(G1341), .Z(new_n1195));
  NAND3_X1  g770(.A1(new_n1172), .A2(new_n1174), .A3(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1066), .A2(new_n1030), .A3(new_n1067), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1194), .B1(new_n1198), .B2(new_n556), .ZN(new_n1199));
  AOI211_X1 g774(.A(KEYINPUT122), .B(new_n626), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1193), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1199), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1198), .A2(new_n1194), .A3(new_n556), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1202), .A2(KEYINPUT59), .A3(new_n1203), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1191), .A2(new_n1192), .A3(new_n1201), .A4(new_n1204), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1177), .A2(new_n1182), .A3(KEYINPUT60), .A4(new_n1179), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1206), .A2(new_n619), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT60), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1207), .B1(new_n1208), .B2(new_n1183), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1188), .B1(new_n1205), .B2(new_n1209), .ZN(new_n1210));
  AND3_X1   g785(.A1(new_n1150), .A2(new_n1162), .A3(new_n1210), .ZN(new_n1211));
  AOI211_X1 g786(.A(new_n1090), .B(G286), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1134), .A2(new_n1111), .A3(new_n1121), .A4(new_n1212), .ZN(new_n1213));
  INV_X1    g788(.A(KEYINPUT63), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT117), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  AND3_X1   g792(.A1(new_n1111), .A2(new_n1212), .A3(KEYINPUT63), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n1131), .A2(new_n1133), .A3(G8), .ZN(new_n1219));
  INV_X1    g794(.A(KEYINPUT118), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1221), .A2(new_n1120), .ZN(new_n1222));
  NOR2_X1   g797(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1223));
  OAI211_X1 g798(.A(new_n1134), .B(new_n1218), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g799(.A1(new_n1213), .A2(KEYINPUT117), .A3(new_n1214), .ZN(new_n1225));
  NAND3_X1  g800(.A1(new_n1217), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  AND2_X1   g801(.A1(new_n1122), .A2(new_n1134), .ZN(new_n1227));
  INV_X1    g802(.A(KEYINPUT62), .ZN(new_n1228));
  INV_X1    g803(.A(new_n1148), .ZN(new_n1229));
  AND2_X1   g804(.A1(new_n1141), .A2(new_n1146), .ZN(new_n1230));
  OAI211_X1 g805(.A(new_n1228), .B(new_n1229), .C1(new_n1230), .C2(new_n1135), .ZN(new_n1231));
  INV_X1    g806(.A(new_n1081), .ZN(new_n1232));
  OAI21_X1  g807(.A(KEYINPUT62), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1233));
  NAND4_X1  g808(.A1(new_n1227), .A2(new_n1231), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  INV_X1    g809(.A(new_n1134), .ZN(new_n1235));
  NAND3_X1  g810(.A1(new_n1105), .A2(new_n1087), .A3(new_n966), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1236), .A2(new_n1103), .ZN(new_n1237));
  AOI22_X1  g812(.A1(new_n1235), .A2(new_n1111), .B1(new_n1091), .B2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g813(.A1(new_n1226), .A2(new_n1234), .A3(new_n1238), .ZN(new_n1239));
  OAI21_X1  g814(.A(new_n1047), .B1(new_n1211), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g815(.A(new_n704), .ZN(new_n1241));
  AOI21_X1  g816(.A(new_n1029), .B1(new_n1032), .B2(new_n1241), .ZN(new_n1242));
  NOR2_X1   g817(.A1(new_n1029), .A2(G1996), .ZN(new_n1243));
  XNOR2_X1  g818(.A(new_n1243), .B(KEYINPUT46), .ZN(new_n1244));
  NOR2_X1   g819(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  XNOR2_X1  g820(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n1246));
  XNOR2_X1  g821(.A(new_n1245), .B(new_n1246), .ZN(new_n1247));
  INV_X1    g822(.A(new_n1042), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n1044), .A2(new_n1034), .ZN(new_n1249));
  XNOR2_X1  g824(.A(new_n1249), .B(KEYINPUT48), .ZN(new_n1250));
  AOI21_X1  g825(.A(new_n1247), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1251));
  NOR3_X1   g826(.A1(new_n1033), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1252));
  NOR2_X1   g827(.A1(new_n775), .A2(G2067), .ZN(new_n1253));
  OAI21_X1  g828(.A(new_n1034), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g829(.A(KEYINPUT126), .ZN(new_n1255));
  NAND2_X1  g830(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g831(.A1(new_n1251), .A2(new_n1256), .ZN(new_n1257));
  NOR2_X1   g832(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1258));
  NOR2_X1   g833(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g834(.A1(new_n1240), .A2(new_n1259), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g835(.A1(new_n924), .A2(new_n932), .ZN(new_n1262));
  OR2_X1    g836(.A1(G227), .A2(new_n465), .ZN(new_n1263));
  NOR3_X1   g837(.A1(G229), .A2(G401), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g838(.A1(new_n1003), .A2(new_n1011), .ZN(new_n1265));
  AND3_X1   g839(.A1(new_n1262), .A2(new_n1264), .A3(new_n1265), .ZN(G308));
  NAND3_X1  g840(.A1(new_n1262), .A2(new_n1264), .A3(new_n1265), .ZN(G225));
endmodule


