//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  XNOR2_X1  g000(.A(KEYINPUT2), .B(G113), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G116), .B(G119), .ZN(new_n189));
  OR2_X1    g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n189), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT30), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT69), .ZN(new_n195));
  INV_X1    g009(.A(G134), .ZN(new_n196));
  OAI22_X1  g010(.A1(new_n195), .A2(KEYINPUT11), .B1(new_n196), .B2(G137), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  INV_X1    g012(.A(G137), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n198), .A2(new_n199), .A3(KEYINPUT69), .A4(G134), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  OAI22_X1  g015(.A1(KEYINPUT69), .A2(new_n198), .B1(new_n199), .B2(G134), .ZN(new_n202));
  OAI21_X1  g016(.A(G131), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n202), .B1(new_n197), .B2(new_n200), .ZN(new_n204));
  INV_X1    g018(.A(G131), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  OR2_X1    g022(.A1(new_n208), .A2(KEYINPUT65), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT0), .A2(G128), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n211), .B1(KEYINPUT65), .B2(new_n208), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n213), .B1(new_n214), .B2(G146), .ZN(new_n215));
  AND2_X1   g029(.A1(KEYINPUT66), .A2(G143), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT66), .A2(G143), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n215), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NOR4_X1   g034(.A1(new_n216), .A2(new_n217), .A3(new_n213), .A4(G146), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n209), .B(new_n212), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n214), .A2(G146), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(new_n218), .B2(new_n219), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT68), .B1(new_n225), .B2(new_n210), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT66), .B(G143), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n223), .B1(new_n227), .B2(G146), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n229), .A3(new_n211), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n207), .A2(new_n222), .A3(new_n226), .A4(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n196), .A2(G137), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n199), .A2(G134), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n205), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(new_n204), .B2(new_n205), .ZN(new_n235));
  INV_X1    g049(.A(G128), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n236), .B1(new_n224), .B2(KEYINPUT1), .ZN(new_n237));
  INV_X1    g051(.A(new_n215), .ZN(new_n238));
  OR2_X1    g052(.A1(KEYINPUT66), .A2(G143), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT66), .A2(G143), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n219), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n239), .A2(KEYINPUT67), .A3(new_n219), .A4(new_n240), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n237), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n236), .A2(KEYINPUT1), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n225), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n235), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  AOI211_X1 g062(.A(new_n193), .B(new_n194), .C1(new_n231), .C2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n222), .A2(new_n226), .A3(new_n230), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n204), .B(G131), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT30), .B1(new_n252), .B2(KEYINPUT64), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n192), .B1(new_n249), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n192), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n231), .A2(new_n255), .A3(new_n248), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n257), .B(G101), .ZN(new_n258));
  INV_X1    g072(.A(G237), .ZN(new_n259));
  INV_X1    g073(.A(G953), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n260), .A3(G210), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n258), .B(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n254), .A2(new_n256), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT31), .ZN(new_n264));
  INV_X1    g078(.A(new_n262), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT28), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n252), .A2(new_n192), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n266), .B1(new_n267), .B2(new_n256), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n256), .A2(new_n266), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n265), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n263), .A2(new_n264), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G472), .ZN(new_n273));
  INV_X1    g087(.A(G902), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n254), .A2(KEYINPUT31), .A3(new_n256), .A4(new_n262), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n272), .A2(new_n273), .A3(new_n274), .A4(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n276), .A2(KEYINPUT32), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(KEYINPUT32), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n231), .A2(new_n255), .A3(new_n248), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n255), .B1(new_n231), .B2(new_n248), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT28), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n281), .A2(KEYINPUT29), .A3(new_n262), .A4(new_n269), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n262), .A3(new_n269), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT29), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n262), .B1(new_n254), .B2(new_n256), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n274), .B(new_n282), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n287), .A2(KEYINPUT70), .A3(G472), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT70), .B1(new_n287), .B2(G472), .ZN(new_n289));
  OAI22_X1  g103(.A1(new_n277), .A2(new_n278), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G214), .B1(G237), .B2(G902), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT6), .ZN(new_n292));
  INV_X1    g106(.A(G116), .ZN(new_n293));
  NOR3_X1   g107(.A1(new_n293), .A2(KEYINPUT5), .A3(G119), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n294), .B1(new_n189), .B2(KEYINPUT5), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n295), .A2(G113), .B1(new_n189), .B2(new_n188), .ZN(new_n296));
  INV_X1    g110(.A(G104), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT3), .B1(new_n297), .B2(G107), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT3), .ZN(new_n299));
  INV_X1    g113(.A(G107), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n300), .A3(G104), .ZN(new_n301));
  INV_X1    g115(.A(G101), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n297), .A2(G107), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n298), .A2(new_n301), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n300), .A2(G104), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n297), .A2(G107), .ZN(new_n306));
  OAI21_X1  g120(.A(G101), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT78), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n304), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n308), .B1(new_n304), .B2(new_n307), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n296), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT82), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n298), .A2(new_n301), .A3(new_n303), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT4), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(G101), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(G101), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(KEYINPUT4), .A3(new_n304), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n192), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT82), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n296), .B(new_n319), .C1(new_n309), .C2(new_n310), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n312), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(G110), .B(G122), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n292), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n312), .A2(new_n322), .A3(new_n318), .A4(new_n320), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT83), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n325), .A2(new_n326), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n324), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n321), .A2(new_n292), .A3(new_n323), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n330), .A2(KEYINPUT84), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(KEYINPUT84), .ZN(new_n332));
  INV_X1    g146(.A(new_n237), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n216), .A2(new_n217), .A3(G146), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n243), .B1(new_n334), .B2(new_n215), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n228), .A2(new_n245), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G125), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n222), .A2(new_n226), .A3(G125), .A4(new_n230), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n260), .A2(G224), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n342), .B(new_n343), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n329), .A2(new_n331), .A3(new_n332), .A4(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(G210), .B1(G237), .B2(G902), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(KEYINPUT7), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n340), .A2(new_n341), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT85), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT85), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n340), .A2(new_n350), .A3(new_n341), .A4(new_n347), .ZN(new_n351));
  INV_X1    g165(.A(new_n347), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n342), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n296), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n304), .A2(new_n307), .ZN(new_n355));
  OR2_X1    g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n322), .B(KEYINPUT8), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n354), .A2(new_n355), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  AND4_X1   g173(.A1(new_n349), .A2(new_n351), .A3(new_n353), .A4(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n325), .B(new_n326), .ZN(new_n361));
  AOI21_X1  g175(.A(G902), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n345), .A2(new_n346), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n346), .B(KEYINPUT86), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(new_n345), .B2(new_n362), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n291), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(G475), .A2(G902), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(G125), .B(G140), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(KEYINPUT88), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G146), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n219), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT87), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n259), .A2(new_n260), .A3(G214), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n375), .B1(new_n218), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(G143), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n259), .A2(new_n260), .A3(G214), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n227), .A2(KEYINPUT87), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(KEYINPUT89), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT18), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(new_n205), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NOR4_X1   g199(.A1(new_n381), .A2(KEYINPUT89), .A3(new_n383), .A4(new_n205), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n374), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n381), .A2(G131), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT90), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n381), .A2(KEYINPUT90), .A3(G131), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n381), .A2(G131), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NOR3_X1   g207(.A1(new_n339), .A2(KEYINPUT16), .A3(G140), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n394), .B1(new_n370), .B2(KEYINPUT16), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G146), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n371), .A2(KEYINPUT19), .ZN(new_n397));
  INV_X1    g211(.A(new_n370), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n397), .B1(KEYINPUT19), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n396), .B1(new_n399), .B2(G146), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n387), .B1(new_n393), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G113), .B(G122), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n402), .B(new_n297), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT17), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n390), .A2(new_n392), .A3(new_n406), .A4(new_n391), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n381), .A2(KEYINPUT90), .A3(G131), .ZN(new_n408));
  AOI21_X1  g222(.A(KEYINPUT90), .B1(new_n381), .B2(G131), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT17), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n395), .B(new_n219), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n407), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(new_n403), .A3(new_n387), .ZN(new_n413));
  AOI211_X1 g227(.A(KEYINPUT20), .B(new_n369), .C1(new_n405), .C2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n405), .A2(new_n413), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n368), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT20), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n260), .A2(G952), .ZN(new_n420));
  NAND2_X1  g234(.A1(G234), .A2(G237), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  XOR2_X1   g237(.A(KEYINPUT21), .B(G898), .Z(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n421), .A2(G902), .A3(G953), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n423), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n227), .A2(G128), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n236), .A2(G143), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(new_n196), .A3(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G116), .B(G122), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(new_n300), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT13), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n431), .B1(new_n430), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT92), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n437), .B1(new_n430), .B2(new_n435), .ZN(new_n438));
  AOI211_X1 g252(.A(KEYINPUT92), .B(KEYINPUT13), .C1(new_n227), .C2(G128), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n432), .B(new_n434), .C1(new_n440), .C2(new_n196), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n293), .A2(KEYINPUT14), .A3(G122), .ZN(new_n442));
  INV_X1    g256(.A(new_n433), .ZN(new_n443));
  OAI211_X1 g257(.A(G107), .B(new_n442), .C1(new_n443), .C2(KEYINPUT14), .ZN(new_n444));
  INV_X1    g258(.A(new_n432), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n196), .B1(new_n430), .B2(new_n431), .ZN(new_n446));
  OAI221_X1 g260(.A(new_n444), .B1(G107), .B2(new_n443), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  XOR2_X1   g261(.A(KEYINPUT9), .B(G234), .Z(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(G217), .A3(new_n260), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n441), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n450), .B1(new_n441), .B2(new_n447), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n274), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G478), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(KEYINPUT15), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n441), .A2(new_n447), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n449), .ZN(new_n459));
  AOI21_X1  g273(.A(G902), .B1(new_n459), .B2(new_n451), .ZN(new_n460));
  INV_X1    g274(.A(new_n456), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n412), .A2(new_n403), .A3(new_n387), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n403), .B1(new_n412), .B2(new_n387), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n274), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  XOR2_X1   g281(.A(KEYINPUT91), .B(G475), .Z(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n419), .A2(new_n429), .A3(new_n464), .A4(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n367), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT23), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n473), .B1(G119), .B2(new_n236), .ZN(new_n474));
  INV_X1    g288(.A(G119), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n475), .A2(KEYINPUT23), .A3(G128), .ZN(new_n476));
  OAI22_X1  g290(.A1(new_n474), .A2(new_n476), .B1(G119), .B2(new_n236), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT71), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n478), .B1(new_n475), .B2(G128), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n236), .A2(KEYINPUT71), .A3(G119), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n479), .A2(new_n480), .B1(new_n475), .B2(G128), .ZN(new_n481));
  XOR2_X1   g295(.A(KEYINPUT24), .B(G110), .Z(new_n482));
  OAI22_X1  g296(.A1(new_n477), .A2(G110), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(new_n396), .A3(new_n373), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(KEYINPUT73), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n411), .B1(new_n481), .B2(new_n482), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n477), .B(KEYINPUT72), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(G110), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT22), .B(G137), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(KEYINPUT74), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n260), .A2(G221), .A3(G234), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n492), .B(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n485), .A2(new_n489), .A3(new_n494), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n274), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT25), .ZN(new_n499));
  INV_X1    g313(.A(G217), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(G234), .B2(new_n274), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT25), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n496), .A2(new_n502), .A3(new_n274), .A4(new_n497), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n499), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT75), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n496), .A2(new_n497), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n501), .A2(G902), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n505), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n496), .A2(KEYINPUT75), .A3(new_n497), .A4(new_n507), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n504), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G221), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n513), .B1(new_n448), .B2(new_n274), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n236), .B1(new_n241), .B2(KEYINPUT1), .ZN(new_n515));
  OAI21_X1  g329(.A(KEYINPUT77), .B1(new_n515), .B2(new_n228), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT77), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT1), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n518), .B1(new_n218), .B2(new_n219), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n517), .B(new_n225), .C1(new_n519), .C2(new_n236), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n516), .A2(new_n520), .A3(new_n337), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n355), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT10), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n317), .A2(new_n315), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n250), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n338), .B(KEYINPUT10), .C1(new_n310), .C2(new_n309), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT79), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n251), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n207), .A2(KEYINPUT79), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n524), .A2(new_n527), .A3(new_n528), .A4(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT10), .B1(new_n521), .B2(new_n355), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n309), .A2(new_n310), .ZN(new_n535));
  AOI22_X1  g349(.A1(new_n333), .A2(new_n335), .B1(new_n228), .B2(new_n245), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n535), .A2(new_n536), .A3(new_n523), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n534), .A2(new_n537), .A3(new_n526), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n533), .B1(new_n538), .B2(new_n251), .ZN(new_n539));
  XOR2_X1   g353(.A(G110), .B(G140), .Z(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(KEYINPUT76), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n260), .A2(G227), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n541), .B(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT81), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n522), .B1(new_n338), .B2(new_n355), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT12), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n547), .A2(KEYINPUT80), .A3(new_n548), .A4(new_n207), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(KEYINPUT80), .ZN(new_n550));
  OR2_X1    g364(.A1(new_n548), .A2(KEYINPUT80), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n244), .A2(new_n247), .A3(new_n355), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(new_n355), .B2(new_n521), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n550), .B(new_n551), .C1(new_n553), .C2(new_n251), .ZN(new_n554));
  AND4_X1   g368(.A1(new_n533), .A2(new_n549), .A3(new_n554), .A4(new_n543), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT81), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n539), .A2(new_n557), .A3(new_n544), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n546), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(G469), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n274), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n560), .A2(new_n274), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n549), .A2(new_n554), .A3(new_n533), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n544), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n544), .B1(new_n538), .B2(new_n532), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n524), .A2(new_n527), .A3(new_n528), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n207), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n562), .B1(new_n569), .B2(G469), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n514), .B1(new_n561), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n290), .A2(new_n472), .A3(new_n512), .A4(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT93), .B(G101), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(G3));
  INV_X1    g388(.A(KEYINPUT20), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(new_n416), .B2(new_n368), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n470), .B1(new_n576), .B2(new_n414), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n452), .A2(KEYINPUT33), .A3(new_n453), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT33), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n459), .B2(new_n451), .ZN(new_n580));
  OAI211_X1 g394(.A(G478), .B(new_n274), .C1(new_n578), .C2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT95), .B(G478), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n460), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(KEYINPUT96), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT96), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n587), .B1(new_n577), .B2(new_n584), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n586), .A2(new_n588), .A3(new_n428), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n345), .A2(KEYINPUT94), .A3(new_n362), .A4(new_n346), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT94), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n363), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n346), .B1(new_n345), .B2(new_n362), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n291), .B(new_n591), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n263), .A2(new_n264), .A3(new_n271), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n275), .A2(new_n274), .ZN(new_n598));
  OAI21_X1  g412(.A(G472), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n276), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(new_n511), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n596), .A2(new_n601), .A3(new_n571), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n590), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT34), .B(G104), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G6));
  NAND2_X1  g419(.A1(new_n470), .A2(new_n463), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT97), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n607), .B1(new_n576), .B2(new_n414), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n418), .A2(KEYINPUT97), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n602), .A2(new_n428), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT35), .B(G107), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G9));
  NOR2_X1   g428(.A1(new_n495), .A2(KEYINPUT36), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n490), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n507), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n504), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n599), .A2(new_n276), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT98), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n599), .A2(new_n621), .A3(new_n276), .A4(new_n618), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(new_n571), .A3(new_n472), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n624), .B(KEYINPUT37), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G110), .ZN(G12));
  INV_X1    g440(.A(KEYINPUT99), .ZN(new_n627));
  INV_X1    g441(.A(G900), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n423), .B1(new_n427), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n610), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n627), .B1(new_n610), .B2(new_n630), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n287), .A2(G472), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT70), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n287), .A2(KEYINPUT70), .A3(G472), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n276), .A2(KEYINPUT32), .ZN(new_n638));
  INV_X1    g452(.A(new_n598), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT32), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n639), .A2(new_n640), .A3(new_n273), .A4(new_n272), .ZN(new_n641));
  AOI22_X1  g455(.A1(new_n636), .A2(new_n637), .B1(new_n638), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n561), .A2(new_n570), .ZN(new_n643));
  INV_X1    g457(.A(new_n514), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n633), .A2(new_n646), .A3(new_n596), .A4(new_n618), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G128), .ZN(G30));
  XNOR2_X1  g462(.A(new_n629), .B(KEYINPUT39), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n571), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT100), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT40), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n638), .A2(new_n641), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n254), .A2(new_n256), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n265), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n279), .A2(new_n280), .ZN(new_n657));
  AOI21_X1  g471(.A(G902), .B1(new_n657), .B2(new_n265), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(G472), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n618), .B1(new_n654), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n291), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n364), .A2(new_n366), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT38), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n464), .B1(new_n419), .B2(new_n470), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n662), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n653), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(new_n218), .ZN(G45));
  NOR2_X1   g483(.A1(new_n585), .A2(new_n629), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n646), .A2(new_n596), .A3(new_n618), .A4(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT101), .B(G146), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G48));
  NAND2_X1  g487(.A1(new_n636), .A2(new_n637), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n511), .B1(new_n674), .B2(new_n654), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n560), .A2(KEYINPUT102), .ZN(new_n676));
  AOI211_X1 g490(.A(KEYINPUT81), .B(new_n543), .C1(new_n567), .C2(new_n533), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n557), .B1(new_n539), .B2(new_n544), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n677), .A2(new_n678), .A3(new_n555), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n676), .B1(new_n679), .B2(G902), .ZN(new_n680));
  INV_X1    g494(.A(new_n676), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n559), .A2(new_n274), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n680), .A2(new_n644), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n595), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n675), .A2(new_n589), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT41), .B(G113), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G15));
  NOR2_X1   g501(.A1(new_n611), .A2(new_n428), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n675), .A2(new_n684), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G116), .ZN(G18));
  NOR3_X1   g504(.A1(new_n577), .A2(new_n428), .A3(new_n463), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n684), .A2(new_n290), .A3(new_n691), .A4(new_n618), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G119), .ZN(G21));
  NOR2_X1   g507(.A1(new_n666), .A2(new_n595), .ZN(new_n694));
  INV_X1    g508(.A(new_n683), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n694), .A2(new_n429), .A3(new_n695), .A4(new_n601), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G122), .ZN(G24));
  INV_X1    g511(.A(new_n670), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n619), .A2(KEYINPUT103), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT103), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n599), .A2(new_n700), .A3(new_n276), .A4(new_n618), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n698), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n684), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(KEYINPUT104), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G125), .ZN(G27));
  NAND2_X1  g519(.A1(new_n345), .A2(new_n362), .ZN(new_n706));
  INV_X1    g520(.A(new_n365), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n291), .A3(new_n363), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n708), .A2(KEYINPUT105), .A3(new_n291), .A4(new_n363), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n571), .A3(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n711), .A2(new_n571), .A3(KEYINPUT106), .A4(new_n712), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n290), .A2(new_n512), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT107), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n675), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n717), .A2(new_n670), .A3(new_n719), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT42), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n698), .A2(KEYINPUT42), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n717), .A2(new_n675), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n205), .ZN(G33));
  NAND3_X1  g541(.A1(new_n717), .A2(new_n675), .A3(new_n633), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G134), .ZN(G36));
  INV_X1    g543(.A(KEYINPUT46), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n569), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(G469), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n730), .B1(new_n734), .B2(new_n562), .ZN(new_n735));
  INV_X1    g549(.A(new_n562), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n733), .A2(KEYINPUT46), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n735), .A2(new_n737), .A3(new_n561), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n644), .ZN(new_n739));
  INV_X1    g553(.A(new_n577), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n584), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n584), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n740), .A2(KEYINPUT109), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n740), .A2(KEYINPUT109), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT43), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n600), .A2(new_n618), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n752), .B(KEYINPUT110), .Z(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n739), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n711), .A2(new_n712), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n757), .A2(new_n649), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n756), .B(new_n758), .C1(new_n755), .C2(new_n754), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G137), .ZN(G39));
  INV_X1    g574(.A(KEYINPUT47), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n739), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n738), .A2(KEYINPUT47), .A3(new_n644), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n757), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n764), .A2(new_n511), .A3(new_n642), .A4(new_n670), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT111), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n766), .B(G140), .Z(G42));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n512), .A2(new_n276), .A3(new_n599), .ZN(new_n769));
  AOI211_X1 g583(.A(new_n422), .B(new_n769), .C1(new_n745), .C2(new_n750), .ZN(new_n770));
  INV_X1    g584(.A(new_n291), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n664), .A2(new_n695), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n757), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(new_n423), .A3(new_n695), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n654), .A2(new_n660), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n512), .ZN(new_n780));
  OR3_X1    g594(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n778), .B1(new_n777), .B2(new_n780), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n781), .A2(new_n740), .A3(new_n746), .A4(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(KEYINPUT50), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n770), .A2(new_n771), .A3(new_n785), .A4(new_n772), .ZN(new_n786));
  INV_X1    g600(.A(new_n777), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n699), .A2(new_n701), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n751), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n775), .A2(new_n783), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n682), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n681), .B1(new_n559), .B2(new_n274), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n514), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n762), .A2(new_n763), .A3(new_n794), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n795), .A2(new_n776), .A3(new_n770), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n768), .B1(new_n790), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n420), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n751), .A2(new_n787), .A3(new_n719), .A4(new_n721), .ZN(new_n799));
  XOR2_X1   g613(.A(new_n799), .B(KEYINPUT48), .Z(new_n800));
  NOR3_X1   g614(.A1(new_n790), .A2(new_n796), .A3(new_n768), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n798), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n694), .A2(new_n661), .A3(new_n571), .A4(new_n630), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n647), .A2(new_n671), .A3(new_n703), .A4(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AND4_X1   g620(.A1(new_n290), .A2(new_n596), .A3(new_n571), .A4(new_n618), .ZN(new_n807));
  AOI22_X1  g621(.A1(new_n807), .A2(new_n633), .B1(new_n702), .B2(new_n684), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n808), .A2(KEYINPUT52), .A3(new_n671), .A4(new_n803), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n740), .A2(new_n463), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n367), .B1(new_n812), .B2(new_n585), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n813), .A2(new_n571), .A3(new_n429), .A4(new_n601), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n624), .A2(new_n814), .A3(new_n572), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n685), .A2(new_n692), .A3(new_n689), .A4(new_n696), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n811), .B(new_n815), .C1(new_n816), .C2(KEYINPUT113), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n816), .A2(KEYINPUT113), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n810), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n585), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n788), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n716), .B2(new_n715), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n290), .A2(new_n571), .A3(new_n618), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n463), .B1(new_n608), .B2(new_n609), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n470), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n823), .A2(new_n757), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n630), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n723), .A2(new_n827), .A3(new_n725), .A4(new_n728), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n819), .A2(new_n828), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n723), .A2(new_n827), .A3(new_n725), .A4(new_n728), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n624), .A2(new_n814), .A3(new_n572), .ZN(new_n831));
  INV_X1    g645(.A(new_n346), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n706), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(new_n592), .A3(new_n363), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n591), .A2(new_n291), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n665), .A2(new_n834), .A3(new_n429), .A4(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n836), .A2(new_n769), .A3(new_n683), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n642), .A2(new_n683), .A3(new_n595), .A4(new_n511), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n837), .B1(new_n838), .B2(new_n688), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n831), .A2(new_n839), .A3(new_n685), .A4(new_n692), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n806), .B2(new_n809), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT53), .B1(new_n830), .B2(new_n841), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n829), .A2(new_n842), .A3(KEYINPUT54), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n830), .A2(new_n841), .A3(KEYINPUT53), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT112), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n840), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n810), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n811), .B1(new_n848), .B2(new_n828), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n830), .A2(new_n841), .A3(KEYINPUT112), .A4(KEYINPUT53), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n846), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n843), .B1(KEYINPUT54), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n586), .A2(new_n588), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n781), .A2(new_n853), .A3(new_n782), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n802), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n770), .A2(new_n684), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT116), .ZN(new_n857));
  OAI22_X1  g671(.A1(new_n855), .A2(new_n857), .B1(G952), .B2(G953), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n793), .B(KEYINPUT49), .Z(new_n859));
  NOR3_X1   g673(.A1(new_n859), .A2(new_n511), .A3(new_n771), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n749), .A2(new_n644), .A3(new_n779), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(new_n664), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n858), .A2(new_n862), .ZN(G75));
  NAND3_X1  g677(.A1(new_n329), .A2(new_n332), .A3(new_n331), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(new_n344), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT55), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n830), .A2(new_n810), .A3(new_n818), .A4(new_n817), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n274), .B1(new_n849), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(G210), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT56), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n260), .A2(G952), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n866), .A2(new_n870), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n873), .B1(new_n868), .B2(new_n707), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n871), .A2(new_n872), .A3(new_n874), .ZN(G51));
  OAI21_X1  g689(.A(KEYINPUT54), .B1(new_n829), .B2(new_n842), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n849), .A2(new_n877), .A3(new_n867), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n879), .B1(new_n880), .B2(new_n562), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n736), .A2(KEYINPUT57), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n559), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n868), .A2(new_n734), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n872), .B1(new_n883), .B2(new_n884), .ZN(G54));
  NAND4_X1  g699(.A1(new_n868), .A2(KEYINPUT58), .A3(G475), .A4(new_n416), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT117), .ZN(new_n887));
  INV_X1    g701(.A(new_n872), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n868), .A2(KEYINPUT58), .A3(G475), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n888), .B1(new_n889), .B2(new_n416), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n887), .A2(new_n890), .ZN(G60));
  INV_X1    g705(.A(KEYINPUT120), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n578), .A2(new_n580), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT118), .Z(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(G478), .A2(G902), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT59), .Z(new_n897));
  NOR2_X1   g711(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT119), .B1(new_n879), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n900));
  INV_X1    g714(.A(new_n898), .ZN(new_n901));
  AOI211_X1 g715(.A(new_n900), .B(new_n901), .C1(new_n876), .C2(new_n878), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n888), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n851), .A2(KEYINPUT54), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n878), .ZN(new_n905));
  INV_X1    g719(.A(new_n897), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n894), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n892), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n877), .B1(new_n849), .B2(new_n867), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n898), .B1(new_n843), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n900), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n879), .A2(KEYINPUT119), .A3(new_n898), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n895), .B1(new_n852), .B2(new_n897), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT120), .A4(new_n888), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n908), .A2(new_n915), .ZN(G63));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT121), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT60), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n829), .B2(new_n842), .ZN(new_n920));
  INV_X1    g734(.A(new_n616), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n888), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n506), .B2(new_n920), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT61), .ZN(G66));
  INV_X1    g738(.A(G224), .ZN(new_n925));
  OAI21_X1  g739(.A(G953), .B1(new_n425), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n847), .B2(G953), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n864), .B1(G898), .B2(new_n260), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(G69));
  OR2_X1    g743(.A1(new_n249), .A2(new_n253), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n399), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n931), .A2(G953), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n765), .A2(new_n759), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT122), .B1(new_n812), .B2(new_n585), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n718), .A2(new_n757), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n812), .A2(KEYINPUT122), .A3(new_n585), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n652), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n808), .A2(new_n671), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT62), .B1(new_n668), .B2(new_n939), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n668), .A2(KEYINPUT62), .A3(new_n939), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n933), .B(new_n937), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n932), .B1(new_n942), .B2(new_n260), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n943), .B1(new_n628), .B2(new_n931), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n723), .A2(new_n725), .A3(new_n728), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT124), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n719), .A2(new_n721), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n739), .A2(new_n649), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n938), .B1(new_n950), .B2(new_n694), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n933), .A2(new_n947), .A3(new_n948), .A4(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n932), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n260), .B1(G227), .B2(G900), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT123), .Z(new_n955));
  NAND3_X1  g769(.A1(new_n944), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n628), .A2(KEYINPUT125), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n628), .A2(KEYINPUT125), .ZN(new_n958));
  OR3_X1    g772(.A1(new_n931), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n954), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n956), .A2(new_n960), .ZN(G72));
  XNOR2_X1  g775(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n273), .A2(new_n274), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n942), .B2(new_n840), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n872), .B1(new_n965), .B2(new_n656), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n964), .B1(new_n952), .B2(new_n840), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n967), .A2(new_n655), .A3(new_n265), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n263), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n964), .B1(new_n970), .B2(new_n286), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT127), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n969), .B1(new_n851), .B2(new_n972), .ZN(G57));
endmodule


