//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G120gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G113gat), .ZN(new_n206));
  INV_X1    g005(.A(G113gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G120gat), .ZN(new_n208));
  AND2_X1   g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n204), .B1(new_n209), .B2(KEYINPUT1), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT73), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n206), .A2(new_n208), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n205), .A2(KEYINPUT73), .A3(G113gat), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n203), .A4(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT28), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(G190gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT68), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT27), .ZN(new_n225));
  INV_X1    g024(.A(G183gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT68), .B1(new_n227), .B2(new_n220), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n219), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT69), .ZN(new_n230));
  INV_X1    g029(.A(G190gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(new_n221), .B2(new_n222), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n218), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n223), .B1(new_n221), .B2(new_n222), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n227), .A2(KEYINPUT68), .A3(new_n220), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n237), .A3(new_n219), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n230), .A2(new_n233), .A3(new_n238), .ZN(new_n239));
  OR2_X1    g038(.A1(KEYINPUT71), .A2(KEYINPUT26), .ZN(new_n240));
  NOR2_X1   g039(.A1(G169gat), .A2(G176gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(KEYINPUT71), .A2(KEYINPUT26), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT26), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT70), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G169gat), .A2(G176gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n247), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n243), .A2(new_n245), .A3(new_n246), .A4(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(G183gat), .A2(G190gat), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT72), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(KEYINPUT72), .A3(new_n250), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n239), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT25), .ZN(new_n255));
  INV_X1    g054(.A(new_n246), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n256), .B1(KEYINPUT23), .B2(new_n241), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT24), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n250), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n226), .A2(new_n231), .ZN(new_n260));
  NAND3_X1  g059(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT65), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n257), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n259), .A2(new_n260), .A3(new_n263), .A4(new_n261), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n265), .B1(KEYINPUT23), .B2(new_n241), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n255), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G169gat), .ZN(new_n268));
  INV_X1    g067(.A(G176gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT23), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n246), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n272), .A2(new_n273), .B1(new_n271), .B2(new_n270), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n260), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT67), .B1(new_n226), .B2(new_n231), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n259), .B(new_n261), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n257), .A2(KEYINPUT66), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n274), .A2(new_n278), .A3(KEYINPUT25), .A4(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n267), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n217), .B1(new_n254), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n254), .A2(new_n217), .A3(new_n281), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G227gat), .A2(G233gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT64), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n285), .A2(KEYINPUT34), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n283), .A2(new_n284), .A3(new_n286), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n289), .B1(KEYINPUT34), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n288), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT32), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT33), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G15gat), .B(G43gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(G71gat), .B(G99gat), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n296), .B(new_n297), .Z(new_n298));
  NAND3_X1  g097(.A1(new_n293), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n298), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n292), .B(KEYINPUT32), .C1(new_n294), .C2(new_n300), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n291), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n291), .B1(new_n299), .B2(new_n301), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT85), .ZN(new_n306));
  INV_X1    g105(.A(G211gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT74), .B(G218gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT22), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G197gat), .B(G204gat), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n307), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(KEYINPUT22), .A3(new_n307), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(G218gat), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  OR2_X1    g114(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT22), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(G197gat), .B(G204gat), .Z(new_n319));
  OAI21_X1  g118(.A(G211gat), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G218gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(new_n321), .A3(new_n313), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n315), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(KEYINPUT75), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n325));
  XOR2_X1   g124(.A(G141gat), .B(G148gat), .Z(new_n326));
  INV_X1    g125(.A(G155gat), .ZN(new_n327));
  INV_X1    g126(.A(G162gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(KEYINPUT2), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n326), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G141gat), .B(G148gat), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n330), .B(new_n329), .C1(new_n334), .C2(KEYINPUT2), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n325), .B1(new_n336), .B2(KEYINPUT3), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(KEYINPUT84), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n324), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G228gat), .A2(G233gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n333), .A2(new_n335), .A3(KEYINPUT78), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT78), .B1(new_n333), .B2(new_n335), .ZN(new_n343));
  OR2_X1    g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n315), .A2(new_n325), .A3(new_n322), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n344), .B1(new_n346), .B2(KEYINPUT3), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n339), .A2(new_n341), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT82), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n315), .A2(KEYINPUT82), .A3(new_n325), .A4(new_n322), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n336), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT83), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n323), .A2(new_n337), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n345), .A2(new_n349), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n358), .A2(new_n352), .A3(new_n351), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n359), .A2(KEYINPUT83), .A3(new_n336), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n356), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n348), .B1(new_n361), .B2(new_n340), .ZN(new_n362));
  XNOR2_X1  g161(.A(G78gat), .B(G106gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT31), .B(G50gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n306), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(G22gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n361), .A2(new_n340), .ZN(new_n369));
  INV_X1    g168(.A(new_n348), .ZN(new_n370));
  AND4_X1   g169(.A1(new_n368), .A2(new_n369), .A3(new_n370), .A4(new_n366), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n368), .B1(new_n362), .B2(new_n366), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n367), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n359), .A2(KEYINPUT83), .A3(new_n336), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT83), .B1(new_n359), .B2(new_n336), .ZN(new_n375));
  INV_X1    g174(.A(new_n357), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n370), .B(new_n366), .C1(new_n377), .C2(new_n341), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(G22gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n369), .A2(new_n370), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n365), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n362), .A2(new_n368), .A3(new_n366), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n379), .A2(new_n381), .A3(new_n306), .A4(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n373), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n305), .A2(new_n384), .ZN(new_n385));
  XOR2_X1   g184(.A(KEYINPUT79), .B(KEYINPUT0), .Z(new_n386));
  XNOR2_X1  g185(.A(G1gat), .B(G29gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n386), .B(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G57gat), .B(G85gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n336), .A2(KEYINPUT3), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n392), .A2(new_n217), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT3), .B1(new_n342), .B2(new_n343), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n210), .A2(new_n215), .A3(new_n333), .A4(new_n335), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n396), .A2(KEYINPUT4), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(KEYINPUT4), .ZN(new_n398));
  NAND2_X1  g197(.A1(G225gat), .A2(G233gat), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n395), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n396), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n403), .B1(new_n344), .B2(new_n216), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n402), .B(KEYINPUT5), .C1(new_n399), .C2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT80), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n398), .B1(new_n397), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n396), .A2(KEYINPUT80), .A3(KEYINPUT4), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n407), .A2(new_n408), .B1(new_n394), .B2(new_n393), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT5), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(new_n399), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n391), .B1(new_n405), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT6), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT81), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n412), .A2(KEYINPUT81), .A3(KEYINPUT6), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n405), .A2(new_n411), .A3(new_n391), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT6), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n415), .B(new_n416), .C1(new_n412), .C2(new_n419), .ZN(new_n420));
  AND2_X1   g219(.A1(G226gat), .A2(G233gat), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n249), .A2(KEYINPUT72), .A3(new_n250), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(new_n251), .ZN(new_n423));
  AOI221_X4 g222(.A(KEYINPUT76), .B1(new_n267), .B2(new_n280), .C1(new_n423), .C2(new_n239), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT76), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n425), .B1(new_n254), .B2(new_n281), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n421), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n254), .A2(new_n281), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n421), .A2(KEYINPUT29), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n427), .A2(new_n430), .A3(new_n324), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT77), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n427), .A2(KEYINPUT77), .A3(new_n430), .A4(new_n324), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n428), .A2(KEYINPUT76), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n254), .A2(new_n425), .A3(new_n281), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n437), .A3(new_n429), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n254), .A2(new_n281), .A3(new_n421), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n323), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G8gat), .B(G36gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(G64gat), .B(G92gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n435), .A2(KEYINPUT30), .A3(new_n442), .A4(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n433), .A2(new_n442), .A3(new_n434), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n445), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n433), .A2(new_n442), .A3(new_n434), .A4(new_n446), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT30), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n420), .A2(new_n447), .A3(new_n449), .A4(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n202), .B1(new_n385), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT92), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n447), .A2(new_n449), .A3(new_n452), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT86), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT86), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n447), .A2(new_n460), .A3(new_n452), .A4(new_n449), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n405), .A2(new_n411), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n462), .B1(new_n405), .B2(new_n411), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n463), .A2(new_n464), .A3(new_n391), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n416), .B(new_n415), .C1(new_n465), .C2(new_n419), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n459), .A2(new_n461), .A3(new_n466), .ZN(new_n467));
  XOR2_X1   g266(.A(KEYINPUT91), .B(KEYINPUT35), .Z(new_n468));
  NAND4_X1  g267(.A1(new_n304), .A2(new_n383), .A3(new_n373), .A4(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n457), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n459), .A2(new_n461), .A3(new_n466), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n472), .A2(KEYINPUT92), .A3(new_n469), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n456), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n407), .A2(new_n408), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n395), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n476), .A2(KEYINPUT87), .A3(new_n400), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT87), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n478), .B1(new_n409), .B2(new_n399), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT39), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n480), .B1(new_n404), .B2(new_n399), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT87), .B1(new_n476), .B2(new_n400), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n409), .A2(new_n478), .A3(new_n399), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n480), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT88), .B1(new_n485), .B2(new_n391), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT39), .B1(new_n477), .B2(new_n479), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT88), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n487), .A2(new_n488), .A3(new_n390), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n482), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT40), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT40), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n492), .B(new_n482), .C1(new_n486), .C2(new_n489), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n465), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n450), .B(KEYINPUT30), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n460), .B1(new_n495), .B2(new_n449), .ZN(new_n496));
  INV_X1    g295(.A(new_n461), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n384), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n448), .A2(KEYINPUT37), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT37), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n433), .A2(new_n442), .A3(new_n501), .A4(new_n434), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(new_n445), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n466), .B1(new_n503), .B2(KEYINPUT38), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n440), .A2(new_n441), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n324), .B1(new_n427), .B2(new_n430), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT37), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT38), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n507), .A2(new_n502), .A3(new_n508), .A4(new_n445), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n509), .A2(KEYINPUT90), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(KEYINPUT90), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n504), .A2(new_n510), .A3(new_n450), .A4(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n498), .A2(new_n499), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n384), .A2(new_n453), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n304), .B(KEYINPUT36), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n474), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT93), .B(G36gat), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(G29gat), .ZN(new_n520));
  OR3_X1    g319(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT94), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G43gat), .B(G50gat), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n520), .B(new_n523), .C1(KEYINPUT15), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(KEYINPUT15), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G99gat), .A2(G106gat), .ZN(new_n529));
  INV_X1    g328(.A(G85gat), .ZN(new_n530));
  INV_X1    g329(.A(G92gat), .ZN(new_n531));
  AOI22_X1  g330(.A1(KEYINPUT8), .A2(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT100), .ZN(new_n533));
  XNOR2_X1  g332(.A(G99gat), .B(G106gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(G85gat), .A2(G92gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n534), .B1(new_n533), .B2(new_n536), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n528), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT41), .ZN(new_n542));
  NAND2_X1  g341(.A1(G232gat), .A2(G233gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n527), .B(KEYINPUT17), .ZN(new_n544));
  OAI221_X1 g343(.A(new_n541), .B1(new_n542), .B2(new_n543), .C1(new_n544), .C2(new_n540), .ZN(new_n545));
  XNOR2_X1  g344(.A(G190gat), .B(G218gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G134gat), .B(G162gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n543), .A2(new_n542), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n547), .B(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT9), .ZN(new_n553));
  INV_X1    g352(.A(G71gat), .ZN(new_n554));
  INV_X1    g353(.A(G78gat), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT98), .ZN(new_n557));
  XOR2_X1   g356(.A(G57gat), .B(G64gat), .Z(new_n558));
  XNOR2_X1  g357(.A(G71gat), .B(G78gat), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT98), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n560), .B(new_n553), .C1(new_n554), .C2(new_n555), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n557), .A2(new_n558), .A3(new_n559), .A4(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT99), .ZN(new_n563));
  INV_X1    g362(.A(new_n559), .ZN(new_n564));
  XNOR2_X1  g363(.A(G57gat), .B(G64gat), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n564), .B1(new_n553), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n562), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n563), .B1(new_n562), .B2(new_n566), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT21), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(new_n307), .ZN(new_n573));
  XOR2_X1   g372(.A(G15gat), .B(G22gat), .Z(new_n574));
  INV_X1    g373(.A(G1gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT96), .ZN(new_n577));
  XNOR2_X1  g376(.A(G15gat), .B(G22gat), .ZN(new_n578));
  XOR2_X1   g377(.A(KEYINPUT95), .B(G1gat), .Z(new_n579));
  INV_X1    g378(.A(KEYINPUT16), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OR3_X1    g380(.A1(new_n578), .A2(KEYINPUT96), .A3(G1gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n577), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(G8gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT97), .ZN(new_n585));
  INV_X1    g384(.A(G8gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n581), .A2(new_n586), .A3(new_n576), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n570), .A2(new_n571), .ZN(new_n589));
  OR3_X1    g388(.A1(new_n588), .A2(G183gat), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(G183gat), .B1(new_n588), .B2(new_n589), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n592), .B1(new_n590), .B2(new_n591), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n573), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n590), .A2(new_n591), .ZN(new_n597));
  INV_X1    g396(.A(new_n592), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n573), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n593), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G127gat), .B(G155gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n596), .A2(new_n601), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n604), .B1(new_n596), .B2(new_n601), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n552), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT101), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT101), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n552), .B(new_n609), .C1(new_n605), .C2(new_n606), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n588), .A2(new_n528), .ZN(new_n612));
  NAND2_X1  g411(.A1(G229gat), .A2(G233gat), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n612), .B(new_n613), .C1(new_n588), .C2(new_n544), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT18), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n585), .A2(new_n527), .A3(new_n587), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n613), .B(KEYINPUT13), .Z(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n527), .B(KEYINPUT17), .Z(new_n621));
  INV_X1    g420(.A(new_n588), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n623), .A2(new_n612), .A3(KEYINPUT18), .A4(new_n613), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n616), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G113gat), .B(G141gat), .ZN(new_n626));
  INV_X1    g425(.A(G197gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT11), .B(G169gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  NAND2_X1  g430(.A1(new_n625), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n631), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n616), .A2(new_n620), .A3(new_n624), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  OAI22_X1  g438(.A1(new_n538), .A2(new_n539), .B1(new_n568), .B2(new_n569), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n533), .A2(new_n536), .ZN(new_n641));
  INV_X1    g440(.A(new_n534), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n562), .A2(new_n566), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(new_n644), .A3(new_n537), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n640), .A2(G230gat), .A3(G233gat), .A4(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n643), .A2(new_n644), .A3(new_n537), .ZN(new_n651));
  INV_X1    g450(.A(new_n569), .ZN(new_n652));
  AOI22_X1  g451(.A1(new_n537), .A2(new_n643), .B1(new_n652), .B2(new_n567), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n650), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n540), .B(KEYINPUT10), .C1(new_n569), .C2(new_n568), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT10), .B1(new_n640), .B2(new_n645), .ZN(new_n658));
  NOR4_X1   g457(.A1(new_n570), .A2(new_n538), .A3(new_n650), .A4(new_n539), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT102), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(G230gat), .A2(G233gat), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n657), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n646), .ZN(new_n663));
  AOI211_X1 g462(.A(new_n639), .B(new_n649), .C1(new_n663), .C2(KEYINPUT103), .ZN(new_n664));
  INV_X1    g463(.A(new_n639), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n654), .A2(new_n656), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n661), .B(KEYINPUT104), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n665), .B1(new_n668), .B2(new_n646), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT105), .B1(new_n664), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n663), .A2(KEYINPUT103), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n671), .A2(new_n665), .A3(new_n648), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n673));
  INV_X1    g472(.A(new_n669), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n611), .A2(new_n636), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n517), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(new_n420), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(new_n575), .ZN(G1324gat));
  NOR2_X1   g479(.A1(new_n496), .A2(new_n497), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(KEYINPUT106), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(KEYINPUT106), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT16), .B(G8gat), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n683), .B(new_n684), .C1(KEYINPUT42), .C2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT42), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n688), .B2(G8gat), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n682), .A2(KEYINPUT42), .A3(new_n686), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(G1325gat));
  INV_X1    g490(.A(new_n678), .ZN(new_n692));
  AOI21_X1  g491(.A(G15gat), .B1(new_n692), .B2(new_n304), .ZN(new_n693));
  INV_X1    g492(.A(new_n515), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G15gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT107), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n693), .B1(new_n692), .B2(new_n696), .ZN(G1326gat));
  NOR2_X1   g496(.A1(new_n678), .A2(new_n499), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT43), .B(G22gat), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  AOI21_X1  g499(.A(new_n552), .B1(new_n474), .B2(new_n516), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n605), .A2(new_n606), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n703), .A2(new_n636), .A3(new_n676), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n705), .A2(G29gat), .A3(new_n420), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT45), .Z(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  INV_X1    g507(.A(new_n552), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n384), .A2(new_n710), .A3(new_n453), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n710), .B1(new_n384), .B2(new_n453), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n513), .A2(new_n515), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n467), .A2(new_n457), .A3(new_n470), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT92), .B1(new_n472), .B2(new_n469), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n455), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n708), .B(new_n709), .C1(new_n714), .C2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n718), .B1(new_n701), .B2(new_n708), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n704), .ZN(new_n720));
  OAI21_X1  g519(.A(G29gat), .B1(new_n720), .B2(new_n420), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n707), .A2(new_n721), .ZN(G1328gat));
  OAI21_X1  g521(.A(new_n519), .B1(new_n720), .B2(new_n681), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n705), .A2(new_n681), .A3(new_n519), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(KEYINPUT109), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n723), .B(new_n726), .C1(new_n727), .C2(new_n724), .ZN(G1329gat));
  NOR3_X1   g527(.A1(new_n705), .A2(G43gat), .A3(new_n305), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n719), .A2(new_n694), .A3(new_n704), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n729), .B1(new_n730), .B2(G43gat), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT47), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT110), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n732), .A2(KEYINPUT110), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1330gat));
  NAND2_X1  g535(.A1(new_n384), .A2(G50gat), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n705), .A2(new_n499), .ZN(new_n738));
  OAI22_X1  g537(.A1(new_n720), .A2(new_n737), .B1(new_n738), .B2(G50gat), .ZN(new_n739));
  XNOR2_X1  g538(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n739), .B(new_n740), .Z(G1331gat));
  NAND3_X1  g540(.A1(new_n513), .A2(new_n713), .A3(new_n515), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n635), .B1(new_n474), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n676), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n611), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n420), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g547(.A1(new_n746), .A2(new_n681), .ZN(new_n749));
  NOR2_X1   g548(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n750));
  AND2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n749), .B2(new_n750), .ZN(G1333gat));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n746), .B2(new_n305), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n743), .A2(KEYINPUT112), .A3(new_n304), .A4(new_n745), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n755), .A2(new_n554), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n694), .A2(G71gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n746), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g559(.A1(new_n746), .A2(new_n499), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(new_n555), .ZN(G1335gat));
  INV_X1    g561(.A(new_n420), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n703), .A2(new_n635), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n676), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n709), .B1(new_n767), .B2(new_n717), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT44), .ZN(new_n769));
  AOI211_X1 g568(.A(new_n764), .B(new_n766), .C1(new_n769), .C2(new_n718), .ZN(new_n770));
  INV_X1    g569(.A(new_n766), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT113), .B1(new_n719), .B2(new_n771), .ZN(new_n772));
  OAI211_X1 g571(.A(G85gat), .B(new_n763), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n709), .B(new_n765), .C1(new_n714), .C2(new_n717), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n474), .A2(new_n742), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n777), .A2(KEYINPUT51), .A3(new_n709), .A4(new_n765), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n779), .A2(new_n763), .A3(new_n676), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n530), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n773), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n773), .A2(KEYINPUT114), .A3(new_n781), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(G1336gat));
  NAND2_X1  g585(.A1(new_n719), .A2(new_n771), .ZN(new_n787));
  OAI21_X1  g586(.A(G92gat), .B1(new_n787), .B2(new_n681), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789));
  INV_X1    g588(.A(new_n779), .ZN(new_n790));
  INV_X1    g589(.A(new_n681), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n791), .A2(new_n531), .A3(new_n676), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n788), .B(new_n789), .C1(new_n790), .C2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n770), .B2(new_n772), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n792), .B(KEYINPUT115), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n794), .A2(G92gat), .B1(new_n779), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n793), .B1(new_n796), .B2(new_n789), .ZN(G1337gat));
  NOR3_X1   g596(.A1(new_n790), .A2(new_n305), .A3(new_n744), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n694), .B1(new_n770), .B2(new_n772), .ZN(new_n799));
  MUX2_X1   g598(.A(new_n798), .B(new_n799), .S(G99gat), .Z(G1338gat));
  INV_X1    g599(.A(G106gat), .ZN(new_n801));
  AND4_X1   g600(.A1(new_n801), .A2(new_n779), .A3(new_n384), .A4(new_n676), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n802), .A2(KEYINPUT53), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n787), .B2(new_n499), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n719), .A2(KEYINPUT116), .A3(new_n384), .A4(new_n771), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(G106gat), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n384), .B1(new_n770), .B2(new_n772), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n802), .B1(new_n809), .B2(G106gat), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(G1339gat));
  OAI211_X1 g611(.A(new_n662), .B(KEYINPUT54), .C1(new_n667), .C2(new_n666), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n666), .A2(new_n814), .A3(new_n667), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n815), .A2(KEYINPUT117), .A3(new_n639), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT117), .B1(new_n815), .B2(new_n639), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n813), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n813), .B(KEYINPUT55), .C1(new_n816), .C2(new_n817), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n635), .A2(new_n672), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n613), .B1(new_n623), .B2(new_n612), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n618), .A2(new_n619), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n630), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n634), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n826), .B1(new_n670), .B2(new_n675), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n822), .B1(new_n827), .B2(KEYINPUT118), .ZN(new_n828));
  INV_X1    g627(.A(new_n826), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n664), .A2(KEYINPUT105), .A3(new_n669), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n673), .B1(new_n672), .B2(new_n674), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n552), .B1(new_n828), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n552), .A2(new_n826), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n836), .A2(new_n672), .A3(new_n820), .A4(new_n821), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n703), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n611), .A2(new_n635), .A3(new_n676), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n763), .B(new_n681), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n385), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(new_n636), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(new_n207), .ZN(G1340gat));
  NOR2_X1   g643(.A1(new_n842), .A2(new_n744), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(new_n205), .ZN(G1341gat));
  NOR2_X1   g645(.A1(new_n842), .A2(new_n702), .ZN(new_n847));
  XOR2_X1   g646(.A(new_n847), .B(G127gat), .Z(G1342gat));
  NAND3_X1  g647(.A1(new_n841), .A2(new_n385), .A3(new_n709), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(G134gat), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT56), .ZN(new_n851));
  OR3_X1    g650(.A1(new_n850), .A2(KEYINPUT119), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT119), .B1(new_n850), .B2(new_n851), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n849), .A2(G134gat), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n852), .A2(new_n853), .A3(new_n854), .A4(new_n855), .ZN(G1343gat));
  OAI21_X1  g655(.A(new_n822), .B1(new_n827), .B2(KEYINPUT120), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n676), .A2(KEYINPUT120), .A3(new_n829), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n552), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n703), .B1(new_n859), .B2(new_n837), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n384), .B1(new_n860), .B2(new_n839), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT57), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n863), .B(new_n384), .C1(new_n838), .C2(new_n839), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n694), .A2(new_n791), .A3(new_n420), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n862), .A2(new_n635), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT122), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n864), .A2(new_n865), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT122), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n868), .A2(new_n869), .A3(new_n635), .A4(new_n862), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n867), .A2(new_n870), .A3(G141gat), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n694), .A2(new_n499), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n840), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(G141gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n876), .A3(new_n635), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n871), .A2(new_n872), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n866), .A2(G141gat), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n877), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT121), .B1(new_n880), .B2(KEYINPUT58), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n882));
  AOI211_X1 g681(.A(new_n882), .B(new_n872), .C1(new_n879), .C2(new_n877), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n878), .B1(new_n881), .B2(new_n883), .ZN(G1344gat));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n862), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n744), .ZN(new_n886));
  INV_X1    g685(.A(G148gat), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n886), .A2(KEYINPUT59), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g687(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n820), .A2(new_n672), .A3(new_n821), .ZN(new_n890));
  AOI22_X1  g689(.A1(new_n832), .A2(new_n833), .B1(new_n635), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n827), .A2(KEYINPUT118), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n709), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n837), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n702), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n839), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n863), .B1(new_n897), .B2(new_n384), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n863), .B(new_n384), .C1(new_n860), .C2(new_n839), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n901), .A2(G148gat), .A3(new_n676), .A4(new_n865), .ZN(new_n902));
  INV_X1    g701(.A(new_n875), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n887), .B1(new_n903), .B2(new_n744), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n889), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n888), .A2(new_n905), .ZN(G1345gat));
  OAI21_X1  g705(.A(G155gat), .B1(new_n885), .B2(new_n702), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n875), .A2(new_n327), .A3(new_n703), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n908), .B1(new_n907), .B2(new_n909), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(G1346gat));
  AOI21_X1  g711(.A(G162gat), .B1(new_n875), .B2(new_n709), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n885), .A2(new_n328), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n709), .ZN(G1347gat));
  NAND3_X1  g714(.A1(new_n897), .A2(new_n420), .A3(new_n791), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n385), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n918), .A2(new_n636), .ZN(new_n919));
  XNOR2_X1  g718(.A(KEYINPUT125), .B(G169gat), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n919), .B(new_n920), .ZN(G1348gat));
  NOR2_X1   g720(.A1(new_n918), .A2(new_n744), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(new_n269), .ZN(G1349gat));
  NAND3_X1  g722(.A1(new_n917), .A2(new_n385), .A3(new_n703), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G183gat), .ZN(new_n925));
  INV_X1    g724(.A(new_n236), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(new_n924), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT60), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n925), .B(new_n929), .C1(new_n926), .C2(new_n924), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1350gat));
  NOR2_X1   g730(.A1(new_n918), .A2(new_n552), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(new_n231), .ZN(new_n934));
  XOR2_X1   g733(.A(KEYINPUT61), .B(G190gat), .Z(new_n935));
  OAI21_X1  g734(.A(new_n934), .B1(new_n932), .B2(new_n935), .ZN(G1351gat));
  AOI21_X1  g735(.A(new_n499), .B1(new_n895), .B2(new_n896), .ZN(new_n937));
  OAI211_X1 g736(.A(KEYINPUT126), .B(new_n899), .C1(new_n937), .C2(new_n863), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n835), .A2(new_n837), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n839), .B1(new_n940), .B2(new_n702), .ZN(new_n941));
  OAI21_X1  g740(.A(KEYINPUT57), .B1(new_n941), .B2(new_n499), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT126), .B1(new_n942), .B2(new_n899), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n694), .A2(new_n681), .A3(new_n763), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n944), .A2(new_n945), .A3(new_n635), .A4(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT126), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n948), .B1(new_n898), .B2(new_n900), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n949), .A2(new_n635), .A3(new_n946), .A4(new_n938), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT127), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n947), .A2(G197gat), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n917), .A2(new_n873), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n954), .A2(new_n627), .A3(new_n635), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n952), .A2(new_n955), .ZN(G1352gat));
  NAND3_X1  g755(.A1(new_n944), .A2(new_n676), .A3(new_n946), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(G204gat), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n953), .A2(G204gat), .A3(new_n744), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n960), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n958), .A2(new_n961), .A3(new_n962), .ZN(G1353gat));
  NAND3_X1  g762(.A1(new_n954), .A2(new_n307), .A3(new_n703), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n901), .A2(new_n703), .A3(new_n946), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n965), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n966));
  AOI21_X1  g765(.A(KEYINPUT63), .B1(new_n965), .B2(G211gat), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(G1354gat));
  AOI21_X1  g767(.A(G218gat), .B1(new_n954), .B2(new_n709), .ZN(new_n969));
  AND4_X1   g768(.A1(new_n316), .A2(new_n944), .A3(new_n317), .A4(new_n946), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n969), .B1(new_n970), .B2(new_n709), .ZN(G1355gat));
endmodule


