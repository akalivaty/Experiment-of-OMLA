//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n212), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT64), .B(G244), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G77), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G50), .A2(G226), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n222), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n230));
  OR2_X1    g0030(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n218), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT66), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  AND2_X1   g0048(.A1(G1), .A2(G13), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G226), .ZN(new_n254));
  AND2_X1   g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  OAI21_X1  g0055(.A(G274), .B1(new_n255), .B2(new_n213), .ZN(new_n256));
  OAI22_X1  g0056(.A1(new_n253), .A2(new_n254), .B1(new_n256), .B2(new_n252), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G222), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n258), .A2(G223), .A3(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(G77), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n260), .B(new_n261), .C1(new_n262), .C2(new_n258), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n255), .A2(new_n213), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n257), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G190), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT9), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n213), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  XOR2_X1   g0070(.A(KEYINPUT8), .B(G58), .Z(new_n271));
  NAND2_X1  g0071(.A1(new_n207), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n271), .A2(new_n273), .B1(G150), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n203), .A2(G20), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n270), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(new_n269), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n206), .A2(G20), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G50), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n280), .A2(new_n283), .B1(new_n202), .B2(new_n279), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n267), .B1(new_n277), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  INV_X1    g0087(.A(G150), .ZN(new_n288));
  INV_X1    g0088(.A(new_n274), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n287), .A2(new_n272), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(G20), .B2(new_n203), .ZN(new_n291));
  OAI211_X1 g0091(.A(KEYINPUT9), .B(new_n284), .C1(new_n291), .C2(new_n270), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT69), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n266), .A2(new_n286), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT10), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n266), .A2(new_n286), .A3(new_n292), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n263), .A2(new_n264), .ZN(new_n298));
  INV_X1    g0098(.A(new_n257), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(KEYINPUT68), .B1(new_n300), .B2(G200), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT68), .ZN(new_n303));
  INV_X1    g0103(.A(G200), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n265), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n296), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n303), .B1(new_n265), .B2(new_n304), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n308), .A2(new_n266), .A3(new_n286), .A4(new_n292), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n295), .B(new_n294), .C1(new_n309), .C2(new_n305), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n284), .B1(new_n291), .B2(new_n270), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(G169), .B2(new_n265), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n300), .A2(G179), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AND3_X1   g0114(.A1(new_n307), .A2(new_n310), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G68), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n279), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n317), .B(KEYINPUT12), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n280), .A2(G68), .A3(new_n281), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT70), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT70), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n318), .A2(new_n322), .A3(new_n319), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n289), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n272), .A2(new_n262), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n269), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n326), .B(KEYINPUT11), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n321), .A2(new_n323), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n258), .A2(G232), .A3(G1698), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n258), .A2(G226), .A3(new_n259), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G97), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n264), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n256), .A2(new_n252), .ZN(new_n334));
  INV_X1    g0134(.A(G41), .ZN(new_n335));
  INV_X1    g0135(.A(G45), .ZN(new_n336));
  AOI21_X1  g0136(.A(G1), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n264), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n334), .B1(G238), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT13), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n333), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n340), .B1(new_n333), .B2(new_n339), .ZN(new_n342));
  OAI21_X1  g0142(.A(G200), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n333), .A2(new_n339), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT13), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n333), .A2(new_n339), .A3(new_n340), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(G190), .A3(new_n346), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n328), .A2(new_n343), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(KEYINPUT71), .A2(KEYINPUT14), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n341), .A2(new_n342), .ZN(new_n351));
  INV_X1    g0151(.A(G169), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n345), .A2(G179), .A3(new_n346), .ZN(new_n354));
  OAI211_X1 g0154(.A(G169), .B(new_n349), .C1(new_n341), .C2(new_n342), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n328), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n348), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI22_X1  g0158(.A1(new_n287), .A2(new_n289), .B1(new_n207), .B2(new_n262), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT15), .B(G87), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n359), .A2(KEYINPUT67), .B1(new_n273), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(KEYINPUT67), .B2(new_n359), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n269), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n262), .B1(new_n206), .B2(G20), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n280), .A2(new_n365), .B1(new_n262), .B2(new_n279), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n258), .A2(G232), .A3(new_n259), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n258), .A2(G238), .A3(G1698), .ZN(new_n369));
  INV_X1    g0169(.A(G107), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n368), .B(new_n369), .C1(new_n370), .C2(new_n258), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n264), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n334), .B1(new_n223), .B2(new_n338), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G200), .ZN(new_n375));
  INV_X1    g0175(.A(new_n374), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G190), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n367), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n364), .A2(new_n366), .B1(new_n352), .B2(new_n374), .ZN(new_n379));
  INV_X1    g0179(.A(G179), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n315), .A2(new_n358), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n280), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n271), .A2(new_n281), .ZN(new_n386));
  OAI22_X1  g0186(.A1(new_n385), .A2(new_n386), .B1(new_n278), .B2(new_n271), .ZN(new_n387));
  INV_X1    g0187(.A(G58), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(new_n316), .ZN(new_n389));
  OAI21_X1  g0189(.A(G20), .B1(new_n389), .B2(new_n201), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n274), .A2(G159), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G33), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT3), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT3), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G33), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT7), .B1(new_n397), .B2(new_n207), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  AOI211_X1 g0199(.A(new_n399), .B(G20), .C1(new_n394), .C2(new_n396), .ZN(new_n400));
  OAI21_X1  g0200(.A(G68), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n392), .B1(new_n401), .B2(KEYINPUT72), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n399), .B1(new_n258), .B2(G20), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n397), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n316), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT72), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT16), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n392), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n401), .A2(KEYINPUT16), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n269), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT73), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT16), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n409), .B1(new_n405), .B2(new_n406), .ZN(new_n414));
  AOI211_X1 g0214(.A(KEYINPUT72), .B(new_n316), .C1(new_n403), .C2(new_n404), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT73), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n405), .A2(new_n392), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n270), .B1(new_n418), .B2(KEYINPUT16), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n387), .B1(new_n412), .B2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n394), .A2(new_n396), .A3(G226), .A4(G1698), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n394), .A2(new_n396), .A3(G223), .A4(new_n259), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G33), .A2(G87), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n264), .ZN(new_n426));
  INV_X1    g0226(.A(G274), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n249), .B2(new_n250), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n338), .A2(G232), .B1(new_n337), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(new_n380), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(G169), .B2(new_n430), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT18), .B1(new_n421), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n387), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n417), .B1(new_n416), .B2(new_n419), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT18), .ZN(new_n438));
  INV_X1    g0238(.A(new_n432), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(G190), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n426), .A2(new_n429), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(G200), .B1(new_n426), .B2(new_n429), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT74), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n430), .A2(new_n304), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n426), .A2(new_n429), .A3(new_n441), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT74), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n449), .B(new_n434), .C1(new_n435), .C2(new_n436), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT17), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(KEYINPUT75), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g0253(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n454), .B1(new_n421), .B2(new_n449), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n433), .B(new_n440), .C1(new_n453), .C2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT76), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n384), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n421), .A2(KEYINPUT18), .A3(new_n432), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n438), .B1(new_n437), .B2(new_n439), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n454), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n450), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n450), .B2(new_n452), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n461), .A2(KEYINPUT76), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n458), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n394), .A2(new_n396), .A3(G257), .A4(G1698), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n394), .A2(new_n396), .A3(G250), .A4(new_n259), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G294), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g0270(.A(KEYINPUT5), .B(G41), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n336), .A2(G1), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n471), .A2(new_n472), .B1(new_n249), .B2(new_n250), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n470), .A2(new_n264), .B1(new_n473), .B2(G264), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT77), .ZN(new_n475));
  AND2_X1   g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  NOR2_X1   g0276(.A1(KEYINPUT5), .A2(G41), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n475), .B1(new_n478), .B2(new_n256), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n428), .A2(KEYINPUT77), .A3(new_n471), .A4(new_n472), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(G169), .B1(new_n474), .B2(new_n481), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n474), .A2(new_n380), .A3(new_n481), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT24), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n394), .A2(new_n396), .A3(new_n207), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT22), .ZN(new_n486));
  OAI21_X1  g0286(.A(G87), .B1(new_n486), .B2(KEYINPUT83), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT83), .ZN(new_n488));
  OAI22_X1  g0288(.A1(new_n485), .A2(new_n487), .B1(new_n488), .B2(KEYINPUT22), .ZN(new_n489));
  INV_X1    g0289(.A(G87), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n490), .B1(new_n488), .B2(KEYINPUT22), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n488), .A2(KEYINPUT22), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n258), .A2(new_n491), .A3(new_n207), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n370), .A2(KEYINPUT23), .A3(G20), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT23), .B1(new_n370), .B2(G20), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G116), .ZN(new_n497));
  OAI22_X1  g0297(.A1(new_n495), .A2(new_n496), .B1(G20), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n484), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  AOI211_X1 g0300(.A(KEYINPUT24), .B(new_n498), .C1(new_n489), .C2(new_n493), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n269), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n206), .A2(G33), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n280), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT25), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n278), .B2(G107), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n279), .A2(KEYINPUT25), .A3(new_n370), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n504), .A2(G107), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI211_X1 g0308(.A(new_n482), .B(new_n483), .C1(new_n502), .C2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n502), .A2(new_n508), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n474), .A2(new_n441), .A3(new_n481), .ZN(new_n511));
  AOI21_X1  g0311(.A(G200), .B1(new_n474), .B2(new_n481), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(KEYINPUT84), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n483), .A2(new_n482), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT84), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n502), .B(new_n508), .C1(new_n511), .C2(new_n512), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n479), .A2(new_n480), .B1(new_n473), .B2(G270), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n394), .A2(new_n396), .A3(G257), .A4(new_n259), .ZN(new_n523));
  INV_X1    g0323(.A(G303), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(new_n258), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n258), .A2(G264), .A3(G1698), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n264), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n280), .A2(G116), .A3(new_n503), .ZN(new_n529));
  INV_X1    g0329(.A(G116), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n279), .A2(new_n530), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n268), .A2(new_n213), .B1(G20), .B2(new_n530), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G283), .ZN(new_n533));
  INV_X1    g0333(.A(G97), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n533), .B(new_n207), .C1(G33), .C2(new_n534), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n532), .A2(KEYINPUT20), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT20), .B1(new_n532), .B2(new_n535), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n529), .B(new_n531), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n528), .A2(G169), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT82), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT21), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n352), .B1(new_n522), .B2(new_n527), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT82), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(new_n543), .A3(new_n538), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n540), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n528), .A2(KEYINPUT21), .A3(G169), .A4(new_n538), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT81), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT81), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n542), .A2(new_n548), .A3(KEYINPUT21), .A4(new_n538), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n522), .A2(new_n527), .A3(G179), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n538), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n538), .B1(new_n528), .B2(G200), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n441), .B2(new_n528), .ZN(new_n555));
  AND4_X1   g0355(.A1(new_n545), .A2(new_n550), .A3(new_n553), .A4(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT80), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n278), .A2(G97), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n280), .A2(new_n503), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(new_n560), .B2(new_n534), .ZN(new_n561));
  XNOR2_X1  g0361(.A(G97), .B(G107), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT6), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NOR3_X1   g0364(.A1(new_n563), .A2(new_n534), .A3(G107), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n567), .A2(G20), .B1(G77), .B2(new_n274), .ZN(new_n568));
  OAI21_X1  g0368(.A(G107), .B1(new_n398), .B2(new_n400), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n561), .B1(new_n570), .B2(new_n269), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n394), .A2(new_n396), .A3(G244), .A4(new_n259), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT4), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n258), .A2(KEYINPUT4), .A3(G244), .A4(new_n259), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n258), .A2(G250), .A3(G1698), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n533), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n264), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n479), .A2(new_n480), .B1(new_n473), .B2(G257), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n578), .A2(new_n441), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(G200), .B1(new_n578), .B2(new_n579), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n571), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n578), .A2(new_n579), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n352), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n565), .B1(new_n563), .B2(new_n562), .ZN(new_n585));
  OAI22_X1  g0385(.A1(new_n585), .A2(new_n207), .B1(new_n262), .B2(new_n289), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n370), .B1(new_n403), .B2(new_n404), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n269), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n561), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n578), .A2(new_n380), .A3(new_n579), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n584), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n582), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n206), .A2(G45), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G250), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n256), .A2(new_n594), .B1(new_n264), .B2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n394), .A2(new_n396), .A3(G244), .A4(G1698), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n394), .A2(new_n396), .A3(G238), .A4(new_n259), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n598), .A3(new_n497), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n596), .B1(new_n599), .B2(new_n264), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n380), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT78), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n394), .A2(new_n396), .A3(new_n207), .A4(G68), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT19), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n272), .B2(new_n534), .ZN(new_n606));
  NAND3_X1  g0406(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n607));
  NOR2_X1   g0407(.A1(G97), .A2(G107), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n207), .A2(new_n607), .B1(new_n608), .B2(new_n490), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n604), .B(new_n606), .C1(new_n609), .C2(KEYINPUT79), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n607), .A2(new_n207), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n608), .A2(new_n490), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT79), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n269), .B1(new_n610), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n504), .A2(new_n361), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n360), .A2(new_n279), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n599), .A2(new_n264), .ZN(new_n620));
  INV_X1    g0420(.A(new_n596), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n352), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n600), .A2(KEYINPUT78), .A3(new_n380), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n603), .A2(new_n619), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n622), .A2(G200), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n613), .A2(new_n614), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n609), .A2(KEYINPUT79), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n627), .A2(new_n628), .A3(new_n604), .A4(new_n606), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n629), .A2(new_n269), .B1(new_n279), .B2(new_n360), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n600), .A2(G190), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n504), .A2(G87), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n626), .A2(new_n630), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n625), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n557), .B1(new_n593), .B2(new_n634), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n622), .A2(new_n602), .A3(G179), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT78), .B1(new_n600), .B2(new_n380), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n619), .A2(new_n623), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n622), .A2(new_n441), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n600), .A2(new_n304), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n616), .A2(new_n632), .A3(new_n618), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n638), .A2(new_n639), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n644), .A2(KEYINPUT80), .A3(new_n592), .A4(new_n582), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n521), .A2(new_n556), .A3(new_n635), .A4(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n466), .A2(new_n646), .ZN(G372));
  INV_X1    g0447(.A(new_n314), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n433), .A2(new_n440), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT85), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n355), .A2(new_n354), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n345), .A2(new_n346), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n349), .B1(new_n653), .B2(G169), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n357), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n348), .B1(new_n655), .B2(new_n382), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(new_n455), .B2(new_n453), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n433), .A2(new_n440), .A3(KEYINPUT85), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n651), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n307), .A2(new_n310), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n648), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n584), .A2(new_n590), .A3(new_n591), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n662), .A2(KEYINPUT26), .A3(new_n625), .A4(new_n633), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n619), .A2(new_n623), .A3(new_n601), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n633), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n664), .B1(new_n666), .B2(new_n592), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  AND4_X1   g0468(.A1(new_n545), .A2(new_n550), .A3(new_n517), .A4(new_n553), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n519), .A2(new_n582), .A3(new_n592), .A4(new_n633), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n668), .B(new_n665), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n458), .A2(new_n465), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n661), .A2(new_n672), .ZN(G369));
  AND2_X1   g0473(.A1(new_n550), .A2(new_n553), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n545), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G213), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n538), .A2(new_n681), .ZN(new_n682));
  MUX2_X1   g0482(.A(new_n675), .B(new_n556), .S(new_n682), .Z(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n510), .A2(new_n681), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n521), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n509), .A2(new_n681), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n684), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n681), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n675), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT86), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n675), .A2(KEYINPUT86), .A3(new_n692), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n688), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n509), .A2(new_n692), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n691), .A2(new_n698), .A3(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n210), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n612), .A2(G116), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G1), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n216), .B2(new_n703), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  INV_X1    g0507(.A(G330), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n635), .A2(new_n645), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(new_n556), .A3(new_n521), .A4(new_n692), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT30), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n578), .A2(new_n474), .A3(new_n600), .A4(new_n579), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n711), .B1(new_n712), .B2(new_n551), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT87), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI211_X1 g0515(.A(KEYINPUT87), .B(new_n711), .C1(new_n712), .C2(new_n551), .ZN(new_n716));
  OR3_X1    g0516(.A1(new_n712), .A2(new_n711), .A3(new_n551), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n600), .A2(G179), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n474), .A2(new_n481), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n583), .A2(new_n718), .A3(new_n528), .A4(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n715), .A2(new_n716), .A3(new_n717), .A4(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT31), .B1(new_n721), .B2(new_n681), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n717), .A2(new_n713), .A3(new_n720), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n681), .A2(KEYINPUT31), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n708), .B1(new_n710), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n671), .A2(new_n692), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT29), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT88), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n732), .B(new_n664), .C1(new_n634), .C2(new_n592), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n662), .A2(KEYINPUT26), .A3(new_n633), .A4(new_n665), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n662), .A2(new_n625), .A3(new_n633), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n732), .B1(new_n736), .B2(new_n664), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n739));
  OAI211_X1 g0539(.A(KEYINPUT29), .B(new_n692), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n731), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n728), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n707), .B1(new_n743), .B2(G1), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT89), .Z(G364));
  NOR2_X1   g0545(.A1(new_n683), .A2(G330), .ZN(new_n746));
  XOR2_X1   g0546(.A(new_n746), .B(KEYINPUT90), .Z(new_n747));
  INV_X1    g0547(.A(G13), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n206), .B1(new_n749), .B2(G45), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n702), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n747), .A2(new_n684), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n701), .A2(new_n397), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G355), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(G116), .B2(new_n210), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n701), .A2(new_n258), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n759), .B1(new_n336), .B2(new_n217), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n244), .A2(new_n336), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G13), .A2(G33), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT91), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n213), .B1(G20), .B2(new_n352), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n752), .B1(new_n762), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n207), .A2(G179), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n772), .A2(G190), .A3(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n490), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n207), .A2(new_n380), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G190), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n775), .A2(G190), .A3(new_n304), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n258), .B1(new_n777), .B2(new_n262), .C1(new_n388), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n775), .A2(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n441), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n774), .B(new_n779), .C1(G50), .C2(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n772), .A2(new_n441), .A3(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n370), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n441), .A2(G179), .A3(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n207), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n534), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n780), .A2(G190), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n784), .B(new_n787), .C1(G68), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n772), .A2(new_n776), .ZN(new_n790));
  INV_X1    g0590(.A(G159), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT32), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n782), .A2(new_n789), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT92), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(KEYINPUT33), .B(G317), .ZN(new_n797));
  INV_X1    g0597(.A(new_n778), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n788), .A2(new_n797), .B1(new_n798), .B2(G322), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT93), .ZN(new_n800));
  INV_X1    g0600(.A(new_n777), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G311), .ZN(new_n802));
  INV_X1    g0602(.A(new_n790), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n258), .B1(new_n803), .B2(G329), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n773), .A2(new_n524), .ZN(new_n805));
  INV_X1    g0605(.A(G294), .ZN(new_n806));
  INV_X1    g0606(.A(G283), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n786), .A2(new_n806), .B1(new_n783), .B2(new_n807), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n805), .B(new_n808), .C1(G326), .C2(new_n781), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n800), .A2(new_n802), .A3(new_n804), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n794), .A2(new_n795), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n796), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n771), .B1(new_n812), .B2(new_n768), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n683), .B2(new_n766), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT94), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n754), .A2(new_n815), .ZN(G396));
  NOR2_X1   g0616(.A1(new_n768), .A2(new_n763), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n258), .B1(new_n803), .B2(G311), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n819), .B1(new_n530), .B2(new_n777), .C1(new_n806), .C2(new_n778), .ZN(new_n820));
  INV_X1    g0620(.A(new_n783), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n781), .A2(G303), .B1(new_n821), .B2(G87), .ZN(new_n822));
  INV_X1    g0622(.A(new_n788), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n807), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n773), .A2(new_n370), .ZN(new_n825));
  NOR4_X1   g0625(.A1(new_n820), .A2(new_n824), .A3(new_n787), .A4(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(G132), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n258), .B1(new_n790), .B2(new_n827), .C1(new_n202), .C2(new_n773), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n786), .A2(new_n388), .B1(new_n783), .B2(new_n316), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n798), .A2(G143), .B1(new_n801), .B2(G159), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G137), .A2(new_n781), .B1(new_n788), .B2(G150), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(KEYINPUT95), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n832), .A2(KEYINPUT95), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n830), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT34), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n828), .B(new_n829), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n826), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n768), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n752), .B1(G77), .B2(new_n818), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n378), .B1(new_n367), .B2(new_n692), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n382), .ZN(new_n844));
  INV_X1    g0644(.A(new_n382), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n692), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n842), .B1(new_n763), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT96), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n729), .A2(new_n847), .ZN(new_n850));
  INV_X1    g0650(.A(new_n847), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n851), .A2(new_n671), .A3(new_n692), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n728), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n752), .B1(new_n728), .B2(new_n853), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n849), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G384));
  NOR2_X1   g0658(.A1(new_n749), .A2(new_n206), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n418), .A2(KEYINPUT16), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n434), .B1(new_n411), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n679), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n861), .B1(new_n439), .B2(new_n862), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n450), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n437), .A2(new_n439), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n679), .B(KEYINPUT97), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n437), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n868), .A2(new_n870), .A3(new_n871), .A4(new_n450), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n456), .A2(new_n864), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT38), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n651), .A2(new_n464), .A3(new_n658), .ZN(new_n875));
  INV_X1    g0675(.A(new_n870), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n868), .A2(new_n870), .A3(new_n450), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT37), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n875), .A2(new_n876), .B1(new_n872), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n874), .B1(new_n879), .B2(KEYINPUT38), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n881), .A2(new_n722), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n646), .B2(new_n681), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n357), .A2(new_n681), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n358), .A2(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n357), .B(new_n681), .C1(new_n356), .C2(new_n348), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n847), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n880), .A2(new_n883), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT40), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n863), .B1(new_n461), .B2(new_n464), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n872), .A2(new_n867), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n453), .A2(new_n455), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n864), .B1(new_n894), .B2(new_n649), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT98), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n872), .A2(new_n867), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT38), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n896), .B1(new_n873), .B2(KEYINPUT38), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n883), .A2(new_n887), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n902), .A2(KEYINPUT40), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n889), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n466), .B1(new_n710), .B2(new_n882), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n708), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n906), .B2(new_n905), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n908), .B(KEYINPUT100), .Z(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT39), .B1(new_n899), .B2(new_n900), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT39), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n912), .B(new_n874), .C1(new_n879), .C2(KEYINPUT38), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n356), .A2(new_n357), .A3(new_n692), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT99), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n651), .A2(new_n658), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n918), .A2(new_n869), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n885), .A2(new_n886), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n852), .B2(new_n846), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n919), .B1(new_n901), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n458), .A2(new_n731), .A3(new_n740), .A4(new_n465), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n661), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n924), .B(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n859), .B1(new_n910), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n910), .B2(new_n927), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n567), .A2(KEYINPUT35), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n567), .A2(KEYINPUT35), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n930), .A2(G116), .A3(new_n214), .A4(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT36), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n216), .A2(new_n262), .A3(new_n389), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n316), .A2(G50), .ZN(new_n935));
  OAI211_X1 g0735(.A(G1), .B(new_n748), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n929), .A2(new_n933), .A3(new_n936), .ZN(G367));
  OAI211_X1 g0737(.A(new_n582), .B(new_n592), .C1(new_n571), .C2(new_n692), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT102), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n592), .B2(new_n692), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OR3_X1    g0741(.A1(new_n691), .A2(KEYINPUT101), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(KEYINPUT101), .B1(new_n691), .B2(new_n941), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n643), .A2(new_n692), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(new_n639), .A3(new_n601), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n666), .B2(new_n945), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n944), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n942), .A2(new_n948), .A3(new_n943), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n939), .A2(new_n517), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n681), .B1(new_n953), .B2(new_n592), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n697), .A2(new_n688), .A3(new_n940), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n954), .B1(new_n955), .B2(KEYINPUT42), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(KEYINPUT42), .B2(new_n955), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n952), .B(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n702), .B(KEYINPUT41), .Z(new_n961));
  NAND3_X1  g0761(.A1(new_n698), .A2(new_n699), .A3(new_n940), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT45), .Z(new_n963));
  NAND2_X1  g0763(.A1(new_n698), .A2(new_n699), .ZN(new_n964));
  XOR2_X1   g0764(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n965));
  NAND3_X1  g0765(.A1(new_n964), .A2(new_n941), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n940), .B1(new_n698), .B2(new_n699), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(new_n965), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n963), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n690), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n689), .A2(new_n695), .A3(new_n696), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n698), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT104), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n972), .A2(new_n973), .A3(new_n684), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n684), .A2(new_n973), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n976), .A2(new_n971), .A3(new_n698), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n743), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n963), .A2(new_n691), .A3(new_n966), .A4(new_n968), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n970), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n961), .B1(new_n983), .B2(new_n743), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n960), .B1(new_n984), .B2(new_n751), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n759), .A2(new_n240), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n769), .B1(new_n210), .B2(new_n360), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n778), .A2(new_n288), .B1(new_n777), .B2(new_n202), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n397), .B(new_n988), .C1(G137), .C2(new_n803), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n773), .A2(new_n388), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n786), .A2(new_n316), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n990), .B(new_n991), .C1(G159), .C2(new_n788), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n781), .A2(G143), .B1(new_n821), .B2(G77), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n989), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n258), .B1(new_n803), .B2(G317), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n534), .B2(new_n783), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(KEYINPUT107), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(KEYINPUT107), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n778), .A2(new_n524), .B1(new_n777), .B2(new_n807), .ZN(new_n999));
  XOR2_X1   g0799(.A(KEYINPUT105), .B(G311), .Z(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n999), .B1(new_n781), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n786), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G107), .A2(new_n1003), .B1(new_n788), .B2(G294), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n997), .A2(new_n998), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(KEYINPUT106), .B1(new_n773), .B2(new_n530), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT46), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n994), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT47), .Z(new_n1009));
  OAI221_X1 g0809(.A(new_n752), .B1(new_n986), .B2(new_n987), .C1(new_n1009), .C2(new_n841), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT108), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n766), .B2(new_n947), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n985), .A2(new_n1012), .ZN(G387));
  OAI21_X1  g0813(.A(new_n742), .B1(new_n975), .B2(new_n978), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n980), .A2(new_n702), .A3(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n788), .A2(new_n271), .B1(new_n801), .B2(G68), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT109), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n258), .B1(new_n790), .B2(new_n288), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G50), .B2(new_n798), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n786), .A2(new_n360), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n262), .A2(new_n773), .B1(new_n783), .B2(new_n534), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(G159), .C2(new_n781), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1017), .A2(new_n1019), .A3(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n798), .A2(G317), .B1(new_n801), .B2(G303), .ZN(new_n1024));
  INV_X1    g0824(.A(G322), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n781), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1024), .B1(new_n823), .B2(new_n1000), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT48), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n786), .A2(new_n807), .B1(new_n773), .B2(new_n806), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1029), .A2(KEYINPUT49), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n258), .B1(new_n803), .B2(G326), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(new_n530), .C2(new_n783), .ZN(new_n1034));
  AOI21_X1  g0834(.A(KEYINPUT49), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1023), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n768), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n704), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n755), .A2(new_n1038), .B1(new_n370), .B2(new_n701), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n237), .A2(new_n336), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n271), .A2(new_n202), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT50), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n704), .B(new_n336), .C1(new_n316), .C2(new_n262), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n758), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1039), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n753), .B1(new_n1045), .B2(new_n769), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1037), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n689), .B2(new_n767), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n979), .B2(new_n751), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1015), .A2(new_n1049), .ZN(G393));
  NAND2_X1  g0850(.A1(new_n970), .A2(new_n982), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n980), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1052), .A2(new_n702), .A3(new_n983), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n970), .A2(new_n751), .A3(new_n982), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n769), .B1(new_n534), .B2(new_n210), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n759), .A2(new_n247), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n752), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n258), .B(new_n784), .C1(G294), .C2(new_n801), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n773), .A2(new_n807), .B1(new_n790), .B2(new_n1025), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1059), .A2(KEYINPUT110), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(KEYINPUT110), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G116), .A2(new_n1003), .B1(new_n788), .B2(G303), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G317), .A2(new_n781), .B1(new_n798), .B2(G311), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT52), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G150), .A2(new_n781), .B1(new_n798), .B2(G159), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT51), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G77), .A2(new_n1003), .B1(new_n788), .B2(G50), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n801), .A2(new_n271), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n397), .B1(new_n803), .B2(G143), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n773), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1071), .A2(G68), .B1(new_n821), .B2(G87), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1063), .A2(new_n1065), .B1(new_n1067), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1057), .B1(new_n1074), .B2(new_n768), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n940), .B2(new_n766), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1053), .A2(new_n1054), .A3(new_n1076), .ZN(G390));
  NAND3_X1  g0877(.A1(new_n883), .A2(G330), .A3(new_n887), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT112), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n708), .B1(new_n710), .B2(new_n882), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(KEYINPUT112), .A3(new_n887), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(KEYINPUT111), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n922), .A2(new_n916), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n911), .A2(new_n913), .A3(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n692), .B1(new_n738), .B2(new_n739), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n844), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n846), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n916), .B1(new_n1089), .B2(new_n920), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n880), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1084), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(KEYINPUT111), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n518), .B1(new_n517), .B2(new_n519), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n635), .B(new_n645), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n556), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n1096), .A2(new_n1097), .A3(new_n681), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n726), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n887), .B(G330), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT113), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n727), .A2(KEYINPUT113), .A3(new_n887), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1093), .A2(new_n1104), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1086), .A2(new_n1091), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1092), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n911), .A2(new_n763), .A3(new_n913), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n752), .B1(new_n271), .B2(new_n818), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n370), .A2(new_n823), .B1(new_n1026), .B2(new_n807), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n783), .A2(new_n316), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n397), .B1(new_n790), .B2(new_n806), .C1(new_n534), .C2(new_n777), .ZN(new_n1112));
  OR4_X1    g0912(.A1(new_n774), .A2(new_n1110), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n786), .A2(new_n262), .B1(new_n778), .B2(new_n530), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT118), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT54), .B(G143), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n788), .A2(G137), .B1(new_n801), .B2(new_n1117), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT117), .Z(new_n1119));
  INV_X1    g0919(.A(G125), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n258), .B1(new_n790), .B2(new_n1120), .C1(new_n778), .C2(new_n827), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1071), .A2(G150), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1121), .B1(KEYINPUT53), .B2(new_n1122), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n786), .A2(new_n791), .B1(new_n783), .B2(new_n202), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(G128), .B2(new_n781), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1123), .B(new_n1125), .C1(KEYINPUT53), .C2(new_n1122), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n1113), .A2(new_n1115), .B1(new_n1119), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1109), .B1(new_n1127), .B2(new_n768), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1107), .A2(new_n751), .B1(new_n1108), .B2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n458), .A2(new_n883), .A3(G330), .A4(new_n465), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n925), .A2(new_n1130), .A3(new_n661), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(KEYINPUT114), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT114), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n925), .A2(new_n1130), .A3(new_n661), .A4(new_n1133), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(G330), .B(new_n851), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n921), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1080), .A2(new_n1137), .A3(new_n1082), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n852), .A2(new_n846), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n883), .A2(G330), .A3(new_n851), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1089), .B1(new_n921), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1104), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT115), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1135), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1138), .A2(new_n1139), .B1(new_n1104), .B2(new_n1142), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1148));
  OAI21_X1  g0948(.A(KEYINPUT115), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1146), .A2(new_n1149), .A3(KEYINPUT116), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT116), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n1150), .A2(new_n1151), .A3(new_n1107), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1105), .A2(new_n1086), .A3(new_n1091), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n1106), .B2(new_n1084), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n702), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1129), .B1(new_n1152), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(KEYINPUT119), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT119), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1159), .B(new_n1129), .C1(new_n1152), .C2(new_n1156), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1158), .A2(new_n1160), .ZN(G378));
  INV_X1    g0961(.A(KEYINPUT57), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n311), .A2(new_n862), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n315), .B(new_n1163), .Z(new_n1164));
  XOR2_X1   g0964(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1165));
  XNOR2_X1  g0965(.A(new_n1164), .B(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n917), .A2(new_n923), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n708), .B1(new_n889), .B2(new_n904), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n916), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n911), .B2(new_n913), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n922), .B1(new_n899), .B2(new_n900), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n918), .B2(new_n869), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1166), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1168), .A2(new_n1169), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1169), .B1(new_n1168), .B2(new_n1174), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1148), .B1(new_n1107), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1162), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1135), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n905), .A2(G330), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1167), .B1(new_n917), .B2(new_n923), .ZN(new_n1183));
  NOR3_X1   g0983(.A1(new_n1171), .A2(new_n1173), .A3(new_n1166), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1168), .A2(new_n1169), .A3(new_n1174), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1181), .A2(new_n1187), .A3(KEYINPUT57), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1180), .A2(new_n702), .A3(new_n1188), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n534), .A2(new_n823), .B1(new_n1026), .B2(new_n530), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n991), .B(new_n1190), .C1(G77), .C2(new_n1071), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n821), .A2(G58), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT120), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n397), .A2(new_n335), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G283), .B2(new_n803), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n798), .A2(G107), .B1(new_n801), .B2(new_n361), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1191), .A2(new_n1193), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT58), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1194), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n1120), .A2(new_n1026), .B1(new_n823), .B2(new_n827), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n798), .A2(G128), .B1(new_n801), .B2(G137), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n773), .B2(new_n1116), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1202), .B(new_n1204), .C1(G150), .C2(new_n1003), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n821), .A2(G159), .ZN(new_n1209));
  AOI211_X1 g1009(.A(G33), .B(G41), .C1(new_n803), .C2(G124), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1201), .B1(new_n1198), .B2(new_n1197), .C1(new_n1207), .C2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n768), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n753), .B1(new_n202), .B2(new_n817), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(new_n1167), .C2(new_n764), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1177), .B2(new_n750), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1189), .A2(new_n1217), .ZN(G375));
  NAND2_X1  g1018(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NOR4_X1   g1020(.A1(new_n1150), .A2(new_n1151), .A3(new_n961), .A4(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n752), .B1(G68), .B2(new_n818), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT121), .Z(new_n1223));
  OAI21_X1  g1023(.A(new_n397), .B1(new_n783), .B2(new_n262), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT122), .Z(new_n1225));
  OAI22_X1  g1025(.A1(new_n777), .A2(new_n370), .B1(new_n790), .B2(new_n524), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G283), .B2(new_n798), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1020), .B1(G116), .B2(new_n788), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n781), .A2(G294), .B1(new_n1071), .B2(G97), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1225), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT123), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(G128), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n777), .A2(new_n288), .B1(new_n790), .B2(new_n1233), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n397), .B(new_n1234), .C1(G137), .C2(new_n798), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G132), .A2(new_n781), .B1(new_n788), .B2(new_n1117), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1003), .A2(G50), .B1(new_n1071), .B2(G159), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1235), .A2(new_n1193), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1232), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1223), .B1(new_n841), .B2(new_n1240), .C1(new_n920), .C2(new_n764), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1147), .B2(new_n750), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1221), .A2(new_n1242), .ZN(G381));
  INV_X1    g1043(.A(new_n1157), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1189), .A2(new_n1244), .A3(new_n1217), .ZN(new_n1245));
  INV_X1    g1045(.A(G390), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(G393), .A2(G396), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1246), .A2(new_n857), .A3(new_n1247), .ZN(new_n1248));
  OR4_X1    g1048(.A1(G387), .A2(new_n1245), .A3(new_n1248), .A4(G381), .ZN(G407));
  OAI211_X1 g1049(.A(G407), .B(G213), .C1(G343), .C2(new_n1245), .ZN(G409));
  INV_X1    g1050(.A(KEYINPUT61), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n680), .A2(G213), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1158), .A2(new_n1189), .A3(new_n1160), .A4(new_n1217), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1177), .A2(new_n1179), .A3(new_n961), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1244), .B1(new_n1254), .B2(new_n1216), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1252), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1252), .A2(G2897), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1146), .A2(new_n1149), .A3(KEYINPUT60), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1219), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT60), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n702), .B1(new_n1219), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1259), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1242), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(G384), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1261), .B1(new_n1258), .B2(new_n1219), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n857), .B1(new_n1266), .B2(new_n1242), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1257), .B1(new_n1268), .B2(KEYINPUT125), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT125), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1257), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n1270), .B(new_n1271), .C1(new_n1265), .C2(new_n1267), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n1269), .A2(new_n1272), .B1(KEYINPUT125), .B2(new_n1268), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1251), .B1(new_n1256), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT127), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT127), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1276), .B(new_n1251), .C1(new_n1256), .C2(new_n1273), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1268), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1256), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(KEYINPUT62), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT62), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1256), .A2(new_n1281), .A3(new_n1278), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1275), .A2(new_n1277), .A3(new_n1280), .A4(new_n1282), .ZN(new_n1283));
  AND2_X1   g1083(.A1(G393), .A2(G396), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(new_n1247), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT126), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1285), .B1(G387), .B2(new_n1286), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n1247), .B(new_n1284), .C1(new_n985), .C2(new_n1012), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1246), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G387), .A2(new_n1285), .ZN(new_n1290));
  AOI21_X1  g1090(.A(KEYINPUT126), .B1(new_n985), .B2(new_n1012), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1290), .B(G390), .C1(new_n1285), .C2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1289), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1283), .A2(new_n1294), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1293), .B(new_n1251), .C1(new_n1256), .C2(new_n1273), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1256), .A2(KEYINPUT63), .A3(new_n1278), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT63), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1279), .A2(KEYINPUT124), .A3(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT124), .B1(new_n1279), .B2(new_n1299), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1297), .B(new_n1298), .C1(new_n1300), .C2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1295), .A2(new_n1302), .ZN(G405));
  INV_X1    g1103(.A(new_n1253), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1157), .B1(new_n1189), .B2(new_n1217), .ZN(new_n1305));
  OR3_X1    g1105(.A1(new_n1304), .A2(new_n1305), .A3(new_n1278), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1278), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1308), .B(new_n1294), .ZN(G402));
endmodule


