//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1146,
    new_n1147, new_n1148, new_n1150, new_n1151, new_n1152, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT65), .B(KEYINPUT0), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G58), .ZN(new_n212));
  INV_X1    g0012(.A(G232), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n214), .B(new_n218), .C1(G107), .C2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G97), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT66), .B(G68), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n207), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n201), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G50), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n211), .B(new_n230), .C1(new_n233), .C2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  AOI21_X1  g0052(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT67), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT67), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G222), .A2(G1698), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(G223), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n264), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n259), .B(new_n268), .C1(G77), .C2(new_n264), .ZN(new_n269));
  INV_X1    g0069(.A(G226), .ZN(new_n270));
  INV_X1    g0070(.A(G1), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(G41), .B2(G45), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n256), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G274), .ZN(new_n274));
  OAI221_X1 g0074(.A(new_n269), .B1(new_n270), .B2(new_n273), .C1(new_n274), .C2(new_n272), .ZN(new_n275));
  INV_X1    g0075(.A(G190), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT9), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n271), .A2(G13), .A3(G20), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n202), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n231), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n284), .B1(G1), .B2(new_n232), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n232), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(G150), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n232), .A2(new_n261), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n286), .A2(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(G20), .B2(new_n203), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n281), .B1(new_n202), .B2(new_n285), .C1(new_n291), .C2(new_n284), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n277), .B1(new_n278), .B2(new_n292), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n275), .A2(G200), .B1(KEYINPUT68), .B2(KEYINPUT10), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n293), .B(new_n294), .C1(new_n278), .C2(new_n292), .ZN(new_n295));
  NOR2_X1   g0095(.A1(KEYINPUT68), .A2(KEYINPUT10), .ZN(new_n296));
  XOR2_X1   g0096(.A(new_n295), .B(new_n296), .Z(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n275), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n299), .B(new_n292), .C1(G179), .C2(new_n275), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT16), .ZN(new_n302));
  INV_X1    g0102(.A(G159), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT71), .B1(new_n289), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(G20), .A2(G33), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT71), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n305), .A2(new_n306), .A3(G159), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n201), .B1(new_n225), .B2(G58), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n308), .B1(new_n309), .B2(new_n232), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n262), .A2(new_n232), .A3(new_n263), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT7), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n262), .A2(KEYINPUT7), .A3(new_n232), .A4(new_n263), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n226), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n302), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  AND2_X1   g0116(.A1(KEYINPUT3), .A2(G33), .ZN(new_n317));
  NOR2_X1   g0117(.A1(KEYINPUT3), .A2(G33), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(KEYINPUT7), .B1(new_n319), .B2(new_n232), .ZN(new_n320));
  INV_X1    g0120(.A(new_n314), .ZN(new_n321));
  OAI21_X1  g0121(.A(G68), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G68), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT66), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT66), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G68), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n326), .A3(G58), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n234), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n328), .A2(G20), .B1(new_n304), .B2(new_n307), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n322), .A2(new_n329), .A3(KEYINPUT16), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n316), .A2(new_n330), .A3(new_n283), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT72), .ZN(new_n332));
  NAND2_X1  g0132(.A1(G33), .A2(G87), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n270), .A2(G1698), .ZN(new_n334));
  OAI221_X1 g0134(.A(new_n334), .B1(G223), .B2(G1698), .C1(new_n317), .C2(new_n318), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n333), .A2(new_n335), .B1(new_n254), .B2(new_n258), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n273), .A2(new_n213), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n272), .A2(new_n274), .ZN(new_n338));
  NOR4_X1   g0138(.A1(new_n336), .A2(new_n276), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G200), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n335), .A2(new_n333), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n338), .B1(new_n341), .B2(new_n259), .ZN(new_n342));
  INV_X1    g0142(.A(new_n337), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n286), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n285), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n280), .B2(new_n346), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT72), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n316), .A2(new_n330), .A3(new_n349), .A4(new_n283), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n332), .A2(new_n345), .A3(new_n348), .A4(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT74), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(KEYINPUT17), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  XOR2_X1   g0155(.A(KEYINPUT74), .B(KEYINPUT17), .Z(new_n356));
  NOR2_X1   g0156(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT75), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n332), .A2(new_n348), .A3(new_n350), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT18), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n336), .A2(new_n338), .A3(new_n337), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G179), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n298), .B2(new_n361), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n359), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n360), .B1(new_n359), .B2(new_n363), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT73), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n359), .A2(new_n363), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT18), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT73), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n359), .A2(new_n360), .A3(new_n363), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT75), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n354), .B(new_n372), .C1(new_n351), .C2(new_n356), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n358), .A2(new_n366), .A3(new_n371), .A4(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n273), .A2(new_n221), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n319), .A2(new_n213), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n266), .ZN(new_n378));
  INV_X1    g0178(.A(G107), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n264), .A2(G1698), .ZN(new_n380));
  OAI221_X1 g0180(.A(new_n378), .B1(new_n379), .B2(new_n264), .C1(new_n380), .C2(new_n227), .ZN(new_n381));
  AOI211_X1 g0181(.A(new_n338), .B(new_n376), .C1(new_n381), .C2(new_n259), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G190), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n346), .A2(new_n305), .B1(G20), .B2(G77), .ZN(new_n384));
  XOR2_X1   g0184(.A(KEYINPUT15), .B(G87), .Z(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n384), .B1(new_n287), .B2(new_n386), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(new_n283), .B1(new_n220), .B2(new_n280), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n220), .B2(new_n285), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n383), .B(new_n390), .C1(new_n340), .C2(new_n382), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n301), .A2(new_n375), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT13), .ZN(new_n393));
  OAI211_X1 g0193(.A(G226), .B(new_n266), .C1(new_n317), .C2(new_n318), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT69), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n264), .A2(KEYINPUT69), .A3(G226), .A4(new_n266), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G97), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n377), .A2(G1698), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n259), .ZN(new_n402));
  INV_X1    g0202(.A(new_n338), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n273), .A2(new_n227), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  AND4_X1   g0205(.A1(new_n393), .A2(new_n402), .A3(new_n403), .A4(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n338), .B1(new_n401), .B2(new_n259), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n393), .B1(new_n407), .B2(new_n405), .ZN(new_n408));
  OAI21_X1  g0208(.A(G169), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT14), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n410), .A2(KEYINPUT70), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  OAI221_X1 g0212(.A(G169), .B1(KEYINPUT70), .B2(new_n410), .C1(new_n406), .C2(new_n408), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n406), .A2(new_n408), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G179), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n410), .A2(KEYINPUT70), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n412), .A2(new_n413), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT12), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n225), .A2(new_n418), .A3(new_n279), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n323), .B1(new_n285), .B2(KEYINPUT12), .ZN(new_n420));
  AOI211_X1 g0220(.A(new_n419), .B(new_n420), .C1(new_n418), .C2(new_n279), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n225), .A2(new_n232), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n289), .A2(new_n202), .B1(new_n287), .B2(new_n220), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n283), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n424), .B(KEYINPUT11), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n417), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(G179), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n382), .A2(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n389), .C1(G169), .C2(new_n382), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n414), .A2(G190), .ZN(new_n432));
  INV_X1    g0232(.A(new_n426), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n432), .B(new_n433), .C1(new_n340), .C2(new_n414), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n392), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n264), .A2(G244), .A3(new_n266), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT4), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n437), .A2(new_n438), .B1(G33), .B2(G283), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n264), .A2(KEYINPUT4), .A3(G244), .A4(new_n266), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT76), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n380), .B2(new_n217), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n264), .A2(KEYINPUT76), .A3(G250), .A4(G1698), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n439), .A2(new_n440), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n259), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n271), .A2(G45), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  XNOR2_X1  g0247(.A(KEYINPUT5), .B(G41), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n253), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G257), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n448), .A2(G274), .A3(new_n447), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n445), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT77), .ZN(new_n453));
  INV_X1    g0253(.A(new_n451), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n454), .B1(new_n444), .B2(new_n259), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT77), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n456), .A3(new_n450), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G190), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n379), .A2(KEYINPUT6), .A3(G97), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n222), .A2(new_n379), .ZN(new_n461));
  NOR2_X1   g0261(.A1(G97), .A2(G107), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n460), .B1(new_n463), .B2(KEYINPUT6), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n464), .A2(G20), .B1(G77), .B2(new_n305), .ZN(new_n465));
  OAI21_X1  g0265(.A(G107), .B1(new_n320), .B2(new_n321), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n284), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n284), .B(new_n279), .C1(G1), .C2(new_n261), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(new_n222), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n279), .A2(G97), .ZN(new_n470));
  NOR3_X1   g0270(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n472), .B1(G200), .B2(new_n452), .ZN(new_n473));
  INV_X1    g0273(.A(new_n452), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n471), .B1(new_n474), .B2(new_n428), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n453), .A2(new_n298), .A3(new_n457), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n459), .A2(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT22), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT84), .ZN(new_n479));
  AOI21_X1  g0279(.A(G20), .B1(new_n262), .B2(new_n263), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n479), .B1(new_n480), .B2(G87), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n232), .B(G87), .C1(new_n317), .C2(new_n318), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(KEYINPUT84), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n478), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT23), .B1(new_n232), .B2(G107), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT23), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(new_n379), .A3(G20), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n232), .A2(G33), .A3(G116), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  XNOR2_X1  g0289(.A(new_n489), .B(KEYINPUT85), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n480), .A2(new_n479), .A3(G87), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n482), .A2(KEYINPUT84), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT22), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n484), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT86), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT86), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n484), .A2(new_n490), .A3(new_n496), .A4(new_n493), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(KEYINPUT24), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT24), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n494), .A2(KEYINPUT86), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n283), .A3(new_n500), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n468), .A2(new_n379), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n280), .B(new_n379), .C1(KEYINPUT87), .C2(KEYINPUT25), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT87), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT25), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n504), .B(new_n505), .C1(new_n279), .C2(G107), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n503), .B(new_n506), .C1(new_n504), .C2(new_n505), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n501), .A2(new_n502), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G294), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n264), .A2(new_n266), .ZN(new_n510));
  OAI221_X1 g0310(.A(new_n509), .B1(new_n380), .B2(new_n223), .C1(new_n217), .C2(new_n510), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n511), .A2(new_n259), .B1(G264), .B2(new_n449), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n451), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(G179), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(new_n298), .B2(new_n513), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n477), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n271), .A2(G45), .A3(G274), .ZN(new_n518));
  XNOR2_X1  g0318(.A(new_n518), .B(KEYINPUT78), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n256), .A2(G250), .A3(new_n446), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n254), .A2(new_n258), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n262), .A2(new_n263), .B1(new_n227), .B2(new_n266), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n221), .A2(G1698), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n522), .A2(new_n523), .B1(G33), .B2(G116), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n519), .B(new_n520), .C1(new_n521), .C2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT79), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n522), .A2(new_n523), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G116), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n259), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n531), .A2(KEYINPUT79), .A3(new_n519), .A4(new_n520), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n276), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT83), .ZN(new_n534));
  XNOR2_X1  g0334(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n468), .A2(new_n216), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n232), .B(G68), .C1(new_n317), .C2(new_n318), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n232), .A2(G33), .A3(G97), .ZN(new_n538));
  AND2_X1   g0338(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n539));
  NOR2_X1   g0339(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NOR3_X1   g0342(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n539), .A2(new_n540), .A3(new_n399), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n544), .B1(new_n545), .B2(G20), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT81), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n542), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  OR2_X1    g0348(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n549));
  AND2_X1   g0349(.A1(G33), .A2(G97), .ZN(new_n550));
  NAND2_X1  g0350(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n543), .B1(new_n552), .B2(new_n232), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n537), .A2(new_n541), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT81), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n548), .A2(new_n555), .A3(new_n283), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n386), .A2(new_n280), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT82), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT82), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n556), .A2(new_n560), .A3(new_n557), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n536), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n527), .A2(new_n532), .A3(G200), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n535), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n556), .A2(new_n560), .A3(new_n557), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n560), .B1(new_n556), .B2(new_n557), .ZN(new_n566));
  OAI22_X1  g0366(.A1(new_n565), .A2(new_n566), .B1(new_n386), .B2(new_n468), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n527), .A2(new_n532), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n428), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n567), .B(new_n569), .C1(G169), .C2(new_n568), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n513), .A2(G200), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n513), .A2(new_n276), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n508), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n264), .A2(G264), .A3(G1698), .ZN(new_n577));
  INV_X1    g0377(.A(G303), .ZN(new_n578));
  OAI221_X1 g0378(.A(new_n577), .B1(new_n578), .B2(new_n264), .C1(new_n510), .C2(new_n223), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n259), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n449), .A2(G270), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n580), .A2(new_n451), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(G116), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n280), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G33), .A2(G283), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n585), .B(new_n232), .C1(G33), .C2(new_n222), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n586), .B(new_n283), .C1(new_n232), .C2(G116), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT20), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n587), .A2(new_n588), .ZN(new_n590));
  OAI221_X1 g0390(.A(new_n584), .B1(new_n583), .B2(new_n468), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n582), .A2(G169), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT21), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n582), .A2(new_n428), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n591), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n582), .A2(new_n591), .A3(KEYINPUT21), .A4(G169), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n594), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n591), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n582), .A2(new_n276), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(G200), .B2(new_n582), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n599), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n436), .A2(new_n517), .A3(new_n576), .A4(new_n603), .ZN(new_n604));
  XNOR2_X1  g0404(.A(new_n604), .B(KEYINPUT88), .ZN(G372));
  NAND2_X1  g0405(.A1(new_n476), .A2(new_n475), .ZN(new_n606));
  OAI21_X1  g0406(.A(KEYINPUT26), .B1(new_n571), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n516), .A2(new_n598), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n501), .A2(new_n502), .ZN(new_n609));
  INV_X1    g0409(.A(new_n574), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n609), .A2(new_n507), .A3(new_n610), .A4(new_n572), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT89), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n525), .A2(G200), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n612), .B1(new_n562), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n536), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n615), .B(new_n613), .C1(new_n565), .C2(new_n566), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n616), .A2(KEYINPUT89), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n535), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n608), .A2(new_n611), .A3(new_n618), .A4(new_n477), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n525), .A2(new_n298), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n567), .A2(new_n569), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT26), .ZN(new_n622));
  INV_X1    g0422(.A(new_n606), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n618), .A2(new_n622), .A3(new_n623), .A4(new_n621), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n607), .A2(new_n619), .A3(new_n621), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n436), .A2(new_n625), .ZN(new_n626));
  AND4_X1   g0426(.A1(new_n373), .A2(new_n431), .A3(new_n358), .A4(new_n434), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n368), .A2(new_n370), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n297), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n629), .A2(new_n300), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n626), .A2(new_n630), .ZN(G369));
  INV_X1    g0431(.A(G13), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n632), .A2(G20), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n271), .ZN(new_n634));
  OR2_X1    g0434(.A1(new_n634), .A2(KEYINPUT27), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(KEYINPUT27), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(G213), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(G343), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n591), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n603), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n598), .B2(new_n640), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G330), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n508), .A2(new_n639), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n516), .B1(new_n575), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n639), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n508), .A2(new_n515), .A3(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT90), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n598), .A2(new_n639), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n654), .A2(new_n648), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n652), .A2(new_n655), .ZN(G399));
  INV_X1    g0456(.A(new_n208), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(G41), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G1), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n543), .A2(new_n583), .ZN(new_n661));
  OAI22_X1  g0461(.A1(new_n660), .A2(new_n661), .B1(new_n235), .B2(new_n659), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT28), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n625), .A2(new_n647), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT29), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n623), .A2(new_n564), .A3(new_n622), .A4(new_n570), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n533), .B(KEYINPUT83), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n562), .A2(new_n612), .A3(new_n613), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n616), .A2(KEYINPUT89), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n621), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n671), .A2(new_n606), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n667), .B1(new_n673), .B2(new_n622), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n619), .A2(new_n621), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n647), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT91), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT91), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n678), .B(new_n647), .C1(new_n674), .C2(new_n675), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n666), .B1(new_n680), .B2(new_n665), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n458), .A2(new_n512), .A3(new_n568), .A4(new_n595), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT30), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n525), .A2(new_n428), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n452), .A2(new_n513), .A3(new_n582), .A4(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n684), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n639), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT31), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n576), .A2(new_n517), .A3(new_n603), .A4(new_n647), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n691), .A2(KEYINPUT31), .A3(new_n689), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n681), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n663), .B1(new_n695), .B2(G1), .ZN(G364));
  AOI21_X1  g0496(.A(new_n660), .B1(G45), .B2(new_n633), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n644), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(G330), .B2(new_n642), .ZN(new_n699));
  INV_X1    g0499(.A(new_n697), .ZN(new_n700));
  INV_X1    g0500(.A(G45), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n236), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n657), .A2(new_n264), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n702), .B(new_n703), .C1(new_n251), .C2(new_n701), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n264), .A2(G355), .A3(new_n208), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n704), .B(new_n705), .C1(G116), .C2(new_n208), .ZN(new_n706));
  NOR2_X1   g0506(.A1(G13), .A2(G33), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G20), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n231), .B1(G20), .B2(new_n298), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n700), .B1(new_n706), .B2(new_n711), .ZN(new_n712));
  XOR2_X1   g0512(.A(new_n712), .B(KEYINPUT92), .Z(new_n713));
  NOR2_X1   g0513(.A1(G179), .A2(G200), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n232), .B1(new_n714), .B2(G190), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n222), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n428), .A2(new_n340), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n232), .A2(G190), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n232), .A2(new_n276), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n340), .A2(G179), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI22_X1  g0524(.A1(G68), .A2(new_n720), .B1(new_n724), .B2(G87), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n718), .A2(new_n722), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n379), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n428), .A2(G200), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n718), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n725), .B(new_n728), .C1(new_n220), .C2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n718), .A2(new_n714), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  XNOR2_X1  g0533(.A(KEYINPUT93), .B(G159), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT32), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n721), .A2(new_n729), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n721), .A2(new_n717), .ZN(new_n738));
  OAI221_X1 g0538(.A(new_n264), .B1(new_n737), .B2(new_n212), .C1(new_n202), .C2(new_n738), .ZN(new_n739));
  OR4_X1    g0539(.A1(new_n716), .A2(new_n731), .A3(new_n736), .A4(new_n739), .ZN(new_n740));
  XOR2_X1   g0540(.A(new_n732), .B(KEYINPUT95), .Z(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n726), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n742), .A2(G329), .B1(G283), .B2(new_n743), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT96), .Z(new_n745));
  INV_X1    g0545(.A(new_n738), .ZN(new_n746));
  INV_X1    g0546(.A(new_n715), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n746), .A2(G326), .B1(new_n747), .B2(G294), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT94), .Z(new_n749));
  NOR2_X1   g0549(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n730), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G311), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n264), .B1(new_n724), .B2(G303), .ZN(new_n753));
  INV_X1    g0553(.A(G317), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(KEYINPUT33), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n754), .A2(KEYINPUT33), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n720), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n750), .A2(new_n752), .A3(new_n753), .A4(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G322), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n737), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n740), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n713), .B1(new_n761), .B2(new_n710), .ZN(new_n762));
  INV_X1    g0562(.A(new_n709), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n762), .B1(new_n642), .B2(new_n763), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n699), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(G396));
  OAI21_X1  g0566(.A(new_n391), .B1(new_n390), .B2(new_n647), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n767), .A2(new_n430), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n430), .A2(new_n639), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n625), .A2(new_n647), .A3(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT99), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n694), .B(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n770), .B1(new_n625), .B2(new_n647), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n700), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n726), .A2(new_n216), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n716), .B(new_n778), .C1(new_n742), .C2(G311), .ZN(new_n779));
  INV_X1    g0579(.A(G283), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n379), .A2(new_n723), .B1(new_n719), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G294), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n737), .A2(new_n782), .B1(new_n730), .B2(new_n583), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n781), .A2(new_n783), .A3(new_n264), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n779), .B(new_n784), .C1(new_n578), .C2(new_n738), .ZN(new_n785));
  INV_X1    g0585(.A(new_n737), .ZN(new_n786));
  XNOR2_X1  g0586(.A(KEYINPUT97), .B(G143), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n786), .A2(new_n787), .B1(new_n751), .B2(new_n734), .ZN(new_n788));
  INV_X1    g0588(.A(G137), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n788), .B1(new_n789), .B2(new_n738), .C1(new_n288), .C2(new_n719), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT34), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n319), .B1(new_n724), .B2(G50), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n790), .A2(new_n791), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n742), .A2(G132), .B1(G58), .B2(new_n747), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n792), .A2(new_n793), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n726), .A2(new_n323), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n785), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n710), .A2(new_n707), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n798), .A2(new_n710), .B1(new_n220), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n697), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT98), .Z(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n708), .B2(new_n770), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n777), .A2(new_n803), .ZN(G384));
  INV_X1    g0604(.A(KEYINPUT104), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n417), .A2(new_n426), .A3(new_n639), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT100), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n426), .A2(new_n639), .ZN(new_n808));
  AND4_X1   g0608(.A1(new_n807), .A2(new_n427), .A3(new_n434), .A4(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n426), .B1(new_n417), .B2(new_n639), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n807), .B1(new_n810), .B2(new_n434), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n806), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(KEYINPUT101), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT101), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n814), .B(new_n806), .C1(new_n809), .C2(new_n811), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  AND3_X1   g0616(.A1(new_n690), .A2(new_n692), .A3(new_n770), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n816), .A2(new_n817), .A3(KEYINPUT40), .ZN(new_n818));
  INV_X1    g0618(.A(new_n637), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n359), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n821), .A2(new_n351), .A3(new_n367), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT103), .ZN(new_n823));
  OAI21_X1  g0623(.A(KEYINPUT37), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR3_X1   g0625(.A1(new_n628), .A2(new_n355), .A3(new_n357), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n822), .B(new_n825), .C1(new_n826), .C2(new_n821), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT38), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n827), .B(new_n828), .C1(new_n822), .C2(new_n825), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n330), .A2(new_n283), .ZN(new_n830));
  AOI21_X1  g0630(.A(KEYINPUT16), .B1(new_n322), .B2(new_n329), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n348), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n832), .A2(new_n819), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n374), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT37), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n822), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n832), .B1(new_n363), .B2(new_n819), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n837), .A2(KEYINPUT37), .A3(new_n351), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n834), .A2(KEYINPUT38), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n829), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n805), .B1(new_n818), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n690), .A2(new_n692), .A3(new_n770), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n815), .B2(new_n813), .ZN(new_n843));
  INV_X1    g0643(.A(new_n840), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n843), .A2(KEYINPUT104), .A3(KEYINPUT40), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n834), .A2(new_n836), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT102), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n847), .A2(new_n848), .A3(KEYINPUT38), .A4(new_n838), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n834), .A2(new_n836), .A3(new_n838), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n828), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n851), .A2(KEYINPUT102), .A3(new_n839), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n843), .A2(new_n849), .A3(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT40), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n846), .A2(new_n855), .A3(G330), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n436), .A2(G330), .A3(new_n693), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT105), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n841), .A2(new_n845), .B1(new_n853), .B2(new_n854), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n860), .A2(new_n436), .A3(new_n693), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT106), .Z(new_n863));
  OAI211_X1 g0663(.A(new_n436), .B(new_n666), .C1(new_n680), .C2(new_n665), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n630), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n863), .B(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n852), .A2(KEYINPUT39), .A3(new_n849), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT39), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n840), .A2(new_n868), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n427), .B(new_n639), .C1(new_n867), .C2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n769), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n813), .A2(new_n815), .B1(new_n871), .B2(new_n771), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(new_n849), .A3(new_n852), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n628), .A2(new_n637), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n866), .B(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n271), .B2(new_n633), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n583), .B1(new_n464), .B2(KEYINPUT35), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n879), .B(new_n233), .C1(KEYINPUT35), .C2(new_n464), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n880), .B(KEYINPUT36), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n236), .A2(G77), .A3(new_n327), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(G50), .B2(new_n323), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(G1), .A3(new_n632), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n878), .A2(new_n881), .A3(new_n884), .ZN(G367));
  NAND2_X1  g0685(.A1(new_n618), .A2(new_n621), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n562), .A2(new_n647), .ZN(new_n887));
  MUX2_X1   g0687(.A(new_n886), .B(new_n621), .S(new_n887), .Z(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n709), .ZN(new_n889));
  OAI22_X1  g0689(.A1(new_n737), .A2(new_n578), .B1(new_n730), .B2(new_n780), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n724), .A2(G116), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT46), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(KEYINPUT110), .ZN(new_n894));
  OAI22_X1  g0694(.A1(new_n754), .A2(new_n732), .B1(new_n715), .B2(new_n379), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n892), .B2(new_n891), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n264), .B1(new_n720), .B2(G294), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n743), .A2(G97), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n894), .A2(new_n896), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  AOI211_X1 g0699(.A(new_n890), .B(new_n899), .C1(G311), .C2(new_n746), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n732), .A2(new_n789), .ZN(new_n901));
  INV_X1    g0701(.A(new_n734), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n902), .A2(new_n719), .B1(new_n730), .B2(new_n202), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n903), .B(KEYINPUT111), .Z(new_n904));
  NOR2_X1   g0704(.A1(new_n726), .A2(new_n220), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n264), .B1(new_n723), .B2(new_n212), .ZN(new_n906));
  AOI211_X1 g0706(.A(new_n905), .B(new_n906), .C1(new_n746), .C2(new_n787), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n904), .B(new_n907), .C1(new_n323), .C2(new_n715), .ZN(new_n908));
  AOI211_X1 g0708(.A(new_n901), .B(new_n908), .C1(G150), .C2(new_n786), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n900), .A2(new_n909), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n910), .B(KEYINPUT47), .Z(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n710), .ZN(new_n912));
  INV_X1    g0712(.A(new_n703), .ZN(new_n913));
  OAI221_X1 g0713(.A(new_n711), .B1(new_n208), .B2(new_n386), .C1(new_n244), .C2(new_n913), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n889), .A2(new_n912), .A3(new_n697), .A4(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n633), .A2(G45), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(G1), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT109), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n477), .B1(new_n471), .B2(new_n647), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n606), .B2(new_n647), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT44), .ZN(new_n921));
  AOI211_X1 g0721(.A(new_n920), .B(new_n655), .C1(KEYINPUT107), .C2(new_n921), .ZN(new_n922));
  OR3_X1    g0722(.A1(new_n922), .A2(KEYINPUT107), .A3(new_n921), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n655), .A2(new_n920), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT45), .Z(new_n925));
  OAI21_X1  g0725(.A(new_n922), .B1(KEYINPUT107), .B2(new_n921), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(new_n651), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT108), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n654), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n649), .A2(KEYINPUT108), .A3(new_n653), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n930), .B(new_n931), .C1(new_n649), .C2(new_n653), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(new_n644), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n695), .A2(new_n933), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n928), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n695), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n658), .B(KEYINPUT41), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n918), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT43), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n888), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n649), .A2(new_n477), .A3(new_n608), .A4(new_n653), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT42), .Z(new_n942));
  AOI21_X1  g0742(.A(new_n516), .B1(new_n459), .B2(new_n473), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n647), .B1(new_n943), .B2(new_n623), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n940), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n888), .A2(new_n939), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n651), .A2(new_n920), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n947), .B(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n915), .B1(new_n938), .B2(new_n949), .ZN(G387));
  NAND2_X1  g0750(.A1(new_n933), .A2(new_n918), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n649), .A2(new_n763), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n703), .B1(new_n241), .B2(new_n701), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n661), .A2(new_n208), .A3(new_n264), .ZN(new_n954));
  AOI211_X1 g0754(.A(G45), .B(new_n661), .C1(G68), .C2(G77), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n286), .A2(G50), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT50), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n953), .A2(new_n954), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n208), .A2(G107), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n711), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(KEYINPUT112), .B(G150), .Z(new_n961));
  AOI22_X1  g0761(.A1(G77), .A2(new_n724), .B1(new_n733), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT113), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n747), .A2(new_n385), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n746), .A2(G159), .B1(new_n751), .B2(G68), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n966), .B(new_n264), .C1(new_n286), .C2(new_n719), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n898), .B1(new_n962), .B2(KEYINPUT113), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n737), .A2(new_n202), .ZN(new_n969));
  NOR4_X1   g0769(.A1(new_n965), .A2(new_n967), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n724), .A2(G294), .B1(new_n747), .B2(G283), .ZN(new_n971));
  AOI22_X1  g0771(.A1(G322), .A2(new_n746), .B1(new_n720), .B2(G311), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n578), .B2(new_n730), .C1(new_n754), .C2(new_n737), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT48), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT114), .Z(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(new_n974), .B2(new_n973), .ZN(new_n977));
  XOR2_X1   g0777(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n978));
  OAI22_X1  g0778(.A1(new_n977), .A2(new_n978), .B1(new_n583), .B2(new_n726), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n264), .B(new_n979), .C1(new_n977), .C2(new_n978), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n733), .A2(G326), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n970), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n710), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n697), .B(new_n960), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n934), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n658), .B1(new_n695), .B2(new_n933), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n951), .B1(new_n952), .B2(new_n984), .C1(new_n985), .C2(new_n986), .ZN(G393));
  AOI21_X1  g0787(.A(new_n659), .B1(new_n928), .B2(new_n934), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n935), .A2(new_n988), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n920), .A2(new_n763), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n711), .B1(new_n222), .B2(new_n208), .C1(new_n248), .C2(new_n913), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n738), .A2(new_n288), .B1(new_n737), .B2(new_n303), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT51), .Z(new_n993));
  AOI22_X1  g0793(.A1(new_n346), .A2(new_n751), .B1(new_n733), .B2(new_n787), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n220), .B2(new_n715), .ZN(new_n995));
  NOR4_X1   g0795(.A1(new_n993), .A2(new_n995), .A3(new_n319), .A4(new_n778), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n202), .B2(new_n719), .C1(new_n226), .C2(new_n723), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT116), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G317), .A2(new_n746), .B1(new_n786), .B2(G311), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT52), .Z(new_n1000));
  AOI21_X1  g0800(.A(new_n264), .B1(new_n751), .B2(G294), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n720), .A2(G303), .B1(new_n747), .B2(G116), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n759), .B2(new_n732), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G283), .B2(new_n724), .ZN(new_n1004));
  AND4_X1   g0804(.A1(new_n728), .A2(new_n1000), .A3(new_n1001), .A4(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n710), .B1(new_n998), .B2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n990), .A2(new_n697), .A3(new_n991), .A4(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n918), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n989), .B(new_n1007), .C1(new_n928), .C2(new_n1008), .ZN(G390));
  NAND3_X1  g0809(.A1(new_n816), .A2(new_n817), .A3(G330), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n677), .A2(new_n679), .A3(new_n871), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n768), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n690), .A2(new_n692), .A3(G330), .A4(new_n770), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1014), .A2(new_n815), .A3(new_n813), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1010), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1010), .A2(new_n1015), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n771), .A2(new_n871), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AND3_X1   g0819(.A1(new_n864), .A2(new_n630), .A3(new_n857), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n427), .A2(new_n639), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n867), .B(new_n869), .C1(new_n1023), .C2(new_n872), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1011), .A2(new_n1012), .A3(new_n816), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n840), .A2(new_n1023), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT117), .ZN(new_n1028));
  AND3_X1   g0828(.A1(new_n1024), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1028), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1029), .A2(new_n1030), .A3(new_n1010), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1010), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1022), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(KEYINPUT117), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1010), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1024), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1039), .A2(new_n1032), .A3(new_n1021), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1034), .A2(new_n658), .A3(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n918), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n867), .A2(new_n869), .A3(new_n707), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n264), .B1(new_n742), .B2(G294), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n220), .B2(new_n715), .C1(new_n780), .C2(new_n738), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n737), .A2(new_n583), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n723), .A2(new_n216), .B1(new_n726), .B2(new_n323), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n719), .A2(new_n379), .B1(new_n730), .B2(new_n222), .ZN(new_n1048));
  NOR4_X1   g0848(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  XOR2_X1   g0849(.A(KEYINPUT54), .B(G143), .Z(new_n1050));
  AOI22_X1  g0850(.A1(new_n742), .A2(G125), .B1(new_n751), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n319), .B1(new_n743), .B2(G50), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT118), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n724), .A2(new_n961), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT53), .Z(new_n1056));
  NAND3_X1  g0856(.A1(new_n1051), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G128), .A2(new_n746), .B1(new_n786), .B2(G132), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT119), .Z(new_n1059));
  NOR2_X1   g0859(.A1(new_n715), .A2(new_n303), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n1052), .A2(new_n1053), .B1(new_n789), .B2(new_n719), .ZN(new_n1061));
  NOR4_X1   g0861(.A1(new_n1057), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n710), .B1(new_n1049), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n799), .A2(new_n286), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1043), .A2(new_n697), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1041), .A2(new_n1042), .A3(new_n1065), .ZN(G378));
  NAND3_X1  g0866(.A1(new_n1034), .A2(KEYINPUT120), .A3(new_n1020), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT120), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1021), .B1(new_n1039), .B2(new_n1032), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1020), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n876), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n292), .A2(new_n819), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n301), .B(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1074), .B(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n856), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1076), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n860), .B2(G330), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1072), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n856), .A2(new_n1076), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n860), .A2(G330), .A3(new_n1078), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1081), .A2(new_n876), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1067), .A2(new_n1071), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT57), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT121), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1067), .A2(new_n1071), .A3(new_n1084), .A4(KEYINPUT57), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1090), .A2(new_n658), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1085), .A2(KEYINPUT121), .A3(new_n1086), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1089), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1076), .A2(new_n707), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n719), .A2(new_n222), .ZN(new_n1095));
  AOI211_X1 g0895(.A(G41), .B(new_n264), .C1(new_n742), .C2(G283), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1096), .B1(new_n212), .B2(new_n726), .C1(new_n386), .C2(new_n730), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1095), .B(new_n1097), .C1(G107), .C2(new_n786), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n724), .A2(G77), .B1(new_n747), .B2(G68), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1098), .B(new_n1099), .C1(new_n583), .C2(new_n738), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT58), .Z(new_n1101));
  AOI22_X1  g0901(.A1(G132), .A2(new_n720), .B1(new_n751), .B2(G137), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n746), .A2(G125), .B1(new_n747), .B2(G150), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n786), .A2(G128), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n724), .B2(new_n1050), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT59), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n261), .ZN(new_n1109));
  AOI211_X1 g0909(.A(G41), .B(new_n1109), .C1(G124), .C2(new_n733), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1110), .B1(new_n1107), .B2(new_n1106), .C1(new_n902), .C2(new_n726), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n202), .B1(new_n317), .B2(G41), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n710), .B1(new_n1101), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n799), .A2(new_n202), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1094), .A2(new_n697), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n1084), .B2(new_n918), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1093), .A2(new_n1118), .ZN(G375));
  OR2_X1    g0919(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1120), .A2(new_n1021), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n937), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT122), .Z(new_n1123));
  NAND2_X1  g0923(.A1(new_n799), .A2(new_n323), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n816), .B2(new_n708), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n726), .A2(new_n212), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1050), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n264), .B1(new_n202), .B2(new_n715), .C1(new_n1127), .C2(new_n719), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1126), .B(new_n1128), .C1(G132), .C2(new_n746), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n786), .A2(G137), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n742), .A2(G128), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G159), .A2(new_n724), .B1(new_n751), .B2(G150), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n741), .A2(new_n578), .B1(new_n583), .B2(new_n719), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G107), .B2(new_n751), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n905), .A2(new_n264), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT123), .Z(new_n1137));
  OAI221_X1 g0937(.A(new_n964), .B1(new_n222), .B2(new_n723), .C1(new_n782), .C2(new_n738), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1135), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n737), .A2(new_n780), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1133), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1125), .B1(new_n710), .B2(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1019), .A2(new_n918), .B1(new_n697), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1123), .A2(new_n1144), .ZN(G381));
  NOR2_X1   g0945(.A1(G375), .A2(G378), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(G387), .A2(G390), .ZN(new_n1147));
  NOR4_X1   g0947(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(G407));
  INV_X1    g0949(.A(new_n1146), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n638), .A2(G213), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT124), .ZN(new_n1152));
  OAI211_X1 g0952(.A(G407), .B(G213), .C1(new_n1150), .C2(new_n1152), .ZN(G409));
  INV_X1    g0953(.A(G378), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1067), .A2(new_n1071), .A3(new_n1084), .A4(new_n937), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(new_n1118), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G375), .B2(G378), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT125), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT60), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1120), .A2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n658), .B(new_n1161), .C1(new_n1121), .C2(new_n1160), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1162), .A2(G384), .A3(new_n1144), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(G384), .B1(new_n1162), .B2(new_n1144), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1159), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1165), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1167), .A2(KEYINPUT125), .A3(new_n1163), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1158), .A2(new_n1151), .A3(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1171), .A2(new_n1152), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(G2897), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1169), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n638), .A2(G213), .A3(G2897), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1173), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n1151), .B2(new_n1158), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT63), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1170), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT61), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(G393), .B(new_n765), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(G387), .A2(G390), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1182), .B1(new_n1184), .B2(new_n1147), .ZN(new_n1185));
  OR2_X1    g0985(.A1(G387), .A2(G390), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1182), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1186), .A2(new_n1187), .A3(new_n1183), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n1085), .A2(KEYINPUT121), .A3(new_n1086), .ZN(new_n1191));
  AOI21_X1  g0991(.A(KEYINPUT121), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1090), .A2(new_n658), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1118), .ZN(new_n1195));
  OAI21_X1  g0995(.A(G378), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1196), .A2(new_n1152), .A3(new_n1156), .A4(new_n1169), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1197), .A2(new_n1179), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1180), .A2(new_n1181), .A3(new_n1190), .A4(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT126), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1196), .A2(new_n1152), .A3(new_n1156), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1175), .A2(new_n1169), .B1(new_n1172), .B2(G2897), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1200), .B1(new_n1203), .B2(new_n1181), .ZN(new_n1204));
  AOI211_X1 g1004(.A(KEYINPUT126), .B(KEYINPUT61), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1197), .A2(KEYINPUT62), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT62), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1158), .A2(new_n1207), .A3(new_n1151), .A4(new_n1169), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1204), .A2(new_n1205), .A3(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1199), .B1(new_n1210), .B2(new_n1190), .ZN(G405));
  NAND2_X1  g1011(.A1(new_n1150), .A2(new_n1196), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1212), .A2(new_n1174), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1171), .B1(new_n1150), .B2(new_n1196), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1189), .A2(KEYINPUT127), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1189), .A2(KEYINPUT127), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  OAI211_X1 g1018(.A(KEYINPUT127), .B(new_n1189), .C1(new_n1213), .C2(new_n1214), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(G402));
endmodule


