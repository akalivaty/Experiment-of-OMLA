//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n832, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1057, new_n1058;
  INV_X1    g000(.A(KEYINPUT103), .ZN(new_n202));
  NAND2_X1  g001(.A1(G229gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT97), .ZN(new_n204));
  INV_X1    g003(.A(G50gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n204), .B1(new_n205), .B2(G43gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(G43gat), .ZN(new_n207));
  INV_X1    g006(.A(G43gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n208), .A2(KEYINPUT97), .A3(G50gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT15), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT98), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(KEYINPUT98), .A3(new_n211), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n208), .A2(G50gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n207), .A2(new_n217), .A3(KEYINPUT15), .ZN(new_n218));
  NAND2_X1  g017(.A1(G29gat), .A2(G36gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NOR3_X1   g020(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n218), .B(new_n219), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n216), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n222), .B1(KEYINPUT96), .B2(new_n220), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(KEYINPUT96), .B2(new_n220), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(new_n219), .ZN(new_n228));
  INV_X1    g027(.A(new_n218), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n225), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT17), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n223), .B1(new_n214), .B2(new_n215), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n218), .B1(new_n227), .B2(new_n219), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n232), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G8gat), .ZN(new_n237));
  INV_X1    g036(.A(G15gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(G22gat), .ZN(new_n239));
  INV_X1    g038(.A(G22gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n240), .A2(G15gat), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT99), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(G15gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n238), .A2(G22gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT99), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G1gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT16), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n242), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(G1gat), .B1(new_n242), .B2(new_n246), .ZN(new_n250));
  OAI211_X1 g049(.A(KEYINPUT100), .B(new_n237), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n245), .B1(new_n243), .B2(new_n244), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n247), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n242), .A2(new_n246), .A3(new_n248), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n237), .A2(KEYINPUT100), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT100), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G8gat), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n254), .A2(new_n255), .A3(new_n256), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n251), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n236), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n233), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT101), .ZN(new_n264));
  AOI211_X1 g063(.A(new_n257), .B(G8gat), .C1(new_n254), .C2(new_n255), .ZN(new_n265));
  AND4_X1   g064(.A1(new_n256), .A2(new_n254), .A3(new_n255), .A4(new_n258), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n251), .A2(KEYINPUT101), .A3(new_n259), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT102), .B1(new_n269), .B2(new_n231), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT102), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n234), .A2(new_n235), .ZN(new_n272));
  AOI211_X1 g071(.A(new_n271), .B(new_n272), .C1(new_n267), .C2(new_n268), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n203), .B(new_n263), .C1(new_n270), .C2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT18), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n202), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n251), .A2(KEYINPUT101), .A3(new_n259), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT101), .B1(new_n251), .B2(new_n259), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n231), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(new_n271), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n269), .A2(KEYINPUT102), .A3(new_n231), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n262), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n282), .A2(KEYINPUT103), .A3(KEYINPUT18), .A4(new_n203), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n276), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n280), .A2(new_n281), .ZN(new_n285));
  INV_X1    g084(.A(new_n269), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n272), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n203), .B(KEYINPUT13), .Z(new_n289));
  AOI22_X1  g088(.A1(new_n288), .A2(new_n289), .B1(new_n274), .B2(new_n275), .ZN(new_n290));
  XNOR2_X1  g089(.A(G113gat), .B(G141gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT94), .B(G197gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(KEYINPUT11), .B(G169gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(KEYINPUT12), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n284), .A2(new_n290), .A3(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(KEYINPUT95), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n299), .B1(new_n284), .B2(new_n290), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(KEYINPUT84), .B(KEYINPUT6), .Z(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G225gat), .A2(G233gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT66), .ZN(new_n306));
  INV_X1    g105(.A(G113gat), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n306), .B1(new_n307), .B2(G120gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT67), .ZN(new_n309));
  INV_X1    g108(.A(G120gat), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n309), .B1(new_n310), .B2(G113gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(KEYINPUT66), .A3(G113gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n307), .A2(KEYINPUT67), .A3(G120gat), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n308), .A2(new_n311), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G134gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G127gat), .ZN(new_n316));
  INV_X1    g115(.A(G127gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G134gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT1), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n314), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT77), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n307), .A2(G120gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n310), .A2(G113gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n319), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n316), .A2(new_n318), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n321), .A2(new_n322), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n322), .B1(new_n321), .B2(new_n327), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT2), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n333), .A2(KEYINPUT76), .B1(G155gat), .B2(G162gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(G141gat), .B(G148gat), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n333), .B1(G155gat), .B2(G162gat), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n332), .B(new_n334), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  AND2_X1   g136(.A1(G141gat), .A2(G148gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(G141gat), .A2(G148gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G155gat), .ZN(new_n341));
  INV_X1    g140(.A(G162gat), .ZN(new_n342));
  OAI21_X1  g141(.A(KEYINPUT2), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(new_n341), .B2(new_n342), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n340), .B(new_n343), .C1(new_n331), .C2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n337), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n337), .A2(new_n346), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT3), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n330), .A2(KEYINPUT79), .A3(new_n348), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n321), .A2(new_n327), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT77), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n321), .A2(new_n327), .A3(new_n322), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n353), .A2(new_n350), .A3(new_n348), .A4(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n305), .B1(new_n351), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT5), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n352), .A2(new_n349), .ZN(new_n360));
  XNOR2_X1  g159(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n363), .B1(KEYINPUT4), .B2(new_n360), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n358), .A2(new_n359), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AND2_X1   g166(.A1(new_n337), .A2(new_n346), .ZN(new_n368));
  NOR3_X1   g167(.A1(new_n328), .A2(new_n329), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n360), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n353), .A2(new_n349), .A3(new_n354), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT82), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n304), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT83), .B1(new_n374), .B2(new_n359), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n369), .A2(new_n370), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n353), .A2(new_n370), .A3(new_n349), .A4(new_n354), .ZN(new_n377));
  INV_X1    g176(.A(new_n360), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n305), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT83), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT5), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n375), .A2(new_n382), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n360), .A2(KEYINPUT81), .A3(new_n361), .ZN(new_n384));
  OR2_X1    g183(.A1(new_n378), .A2(KEYINPUT4), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n386), .B1(new_n378), .B2(new_n362), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n384), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n358), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n367), .B1(new_n383), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G1gat), .B(G29gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(KEYINPUT0), .ZN(new_n392));
  XNOR2_X1  g191(.A(G57gat), .B(G85gat), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n392), .B(new_n393), .Z(new_n394));
  AOI21_X1  g193(.A(new_n303), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n394), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n375), .A2(new_n382), .B1(new_n358), .B2(new_n388), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n396), .B1(new_n397), .B2(new_n367), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT5), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n381), .B1(new_n380), .B2(KEYINPUT5), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n389), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n366), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT85), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n403), .A2(new_n404), .A3(new_n396), .A4(new_n303), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT85), .B1(new_n398), .B2(new_n302), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n399), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT74), .ZN(new_n408));
  AND2_X1   g207(.A1(G226gat), .A2(G233gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT29), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT25), .ZN(new_n413));
  NOR2_X1   g212(.A1(G169gat), .A2(G176gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT23), .ZN(new_n415));
  NAND2_X1  g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT23), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n417), .B1(G169gat), .B2(G176gat), .ZN(new_n418));
  AND4_X1   g217(.A1(new_n413), .A2(new_n415), .A3(new_n416), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G183gat), .A2(G190gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT24), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT24), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n422), .A2(G183gat), .A3(G190gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n424), .B1(G183gat), .B2(G190gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n427));
  INV_X1    g226(.A(G190gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT64), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT64), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(G190gat), .ZN(new_n431));
  INV_X1    g230(.A(G183gat), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n427), .B1(new_n433), .B2(new_n424), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n426), .B1(new_n434), .B2(new_n413), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n414), .A2(KEYINPUT26), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT26), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n416), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n436), .B(new_n420), .C1(new_n438), .C2(new_n414), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT28), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT64), .B(G190gat), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT27), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT65), .B1(new_n442), .B2(G183gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n432), .A2(KEYINPUT27), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n442), .A2(G183gat), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT65), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n440), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n441), .A2(KEYINPUT28), .A3(new_n445), .A4(new_n446), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n439), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n412), .B1(new_n435), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n439), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n443), .A2(new_n429), .A3(new_n431), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n445), .A2(new_n446), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT65), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT28), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n449), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n452), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n433), .A2(new_n424), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n462), .A2(KEYINPUT25), .B1(new_n425), .B2(new_n419), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(new_n463), .A3(new_n410), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT22), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT72), .B(G211gat), .ZN(new_n466));
  INV_X1    g265(.A(G218gat), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G197gat), .B(G204gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G211gat), .B(G218gat), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(KEYINPUT73), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n472), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n474), .A2(new_n468), .A3(new_n469), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n451), .A2(new_n464), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n476), .B1(new_n451), .B2(new_n464), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n408), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n451), .A2(new_n464), .ZN(new_n480));
  INV_X1    g279(.A(new_n476), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n451), .A2(new_n464), .A3(new_n476), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(KEYINPUT74), .A3(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G8gat), .B(G36gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(KEYINPUT75), .ZN(new_n486));
  XNOR2_X1  g285(.A(G64gat), .B(G92gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n479), .A2(new_n484), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT30), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n482), .A2(new_n483), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(new_n489), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT30), .A4(new_n488), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n490), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n407), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT86), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT86), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n407), .A2(new_n499), .A3(new_n496), .ZN(new_n500));
  INV_X1    g299(.A(new_n352), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n459), .A2(new_n463), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT68), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n459), .A2(new_n463), .A3(KEYINPUT68), .A4(new_n501), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n352), .B1(new_n435), .B2(new_n450), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(G227gat), .A2(G233gat), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT71), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT32), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n511), .B1(new_n507), .B2(new_n508), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT33), .B1(new_n507), .B2(new_n508), .ZN(new_n513));
  XOR2_X1   g312(.A(G15gat), .B(G43gat), .Z(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT69), .ZN(new_n515));
  XNOR2_X1  g314(.A(G71gat), .B(G99gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n512), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT33), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT70), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n520), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(new_n521), .B2(new_n517), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n512), .A2(new_n523), .ZN(new_n524));
  NOR3_X1   g323(.A1(new_n519), .A2(new_n524), .A3(KEYINPUT34), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT34), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n507), .A2(new_n508), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT32), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n520), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n529), .A3(new_n517), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n523), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n526), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n510), .B1(new_n525), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT34), .B1(new_n519), .B2(new_n524), .ZN(new_n534));
  INV_X1    g333(.A(new_n510), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n530), .A2(new_n526), .A3(new_n531), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G78gat), .B(G106gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT31), .B(G50gat), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n539), .B(new_n540), .Z(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n348), .A2(new_n411), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n481), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(G228gat), .ZN(new_n545));
  INV_X1    g344(.A(G233gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n347), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT29), .B1(new_n470), .B2(new_n471), .ZN(new_n551));
  INV_X1    g350(.A(new_n471), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n468), .A2(new_n552), .A3(new_n469), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n550), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n554), .A2(new_n368), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT29), .B1(new_n473), .B2(new_n475), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n349), .B1(new_n557), .B2(KEYINPUT3), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n548), .B1(new_n558), .B2(new_n544), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n556), .A2(new_n559), .A3(G22gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n544), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n547), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n544), .B(new_n548), .C1(new_n368), .C2(new_n554), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n240), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n542), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT88), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g366(.A(KEYINPUT88), .B(new_n542), .C1(new_n560), .C2(new_n564), .ZN(new_n568));
  OAI21_X1  g367(.A(G22gat), .B1(new_n556), .B2(new_n559), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n562), .A2(new_n240), .A3(new_n563), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n570), .A3(new_n541), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT87), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT87), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n569), .A2(new_n570), .A3(new_n573), .A4(new_n541), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n567), .A2(new_n568), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n538), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT90), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n398), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n403), .A2(KEYINPUT90), .A3(new_n396), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n395), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n581), .A2(new_n405), .A3(new_n406), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n577), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT36), .ZN(new_n585));
  AND3_X1   g384(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n535), .B1(new_n534), .B2(new_n536), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n533), .A2(KEYINPUT36), .A3(new_n537), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n588), .A2(new_n575), .A3(new_n589), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n498), .B(new_n500), .C1(new_n584), .C2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT37), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT92), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n478), .B1(new_n483), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n477), .A2(KEYINPUT92), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n482), .A2(new_n592), .A3(new_n483), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT38), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(new_n598), .A3(new_n489), .ZN(new_n599));
  OAI22_X1  g398(.A1(new_n596), .A2(new_n599), .B1(new_n489), .B2(new_n492), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n479), .A2(new_n484), .A3(KEYINPUT37), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n489), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT93), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT93), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n601), .A2(new_n604), .A3(new_n489), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n603), .A2(new_n605), .A3(new_n597), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n600), .B1(new_n606), .B2(KEYINPUT38), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n581), .A2(new_n405), .A3(new_n406), .A4(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n364), .B1(new_n351), .B2(new_n357), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n609), .A2(new_n304), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n371), .A2(new_n304), .A3(new_n373), .ZN(new_n613));
  OAI211_X1 g412(.A(KEYINPUT39), .B(new_n613), .C1(new_n609), .C2(new_n304), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT40), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT89), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n612), .A2(new_n614), .A3(new_n394), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(new_n495), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n396), .B1(new_n610), .B2(new_n611), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n616), .B1(new_n619), .B2(new_n614), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n621), .A2(new_n579), .A3(new_n580), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT91), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n621), .A2(new_n579), .A3(KEYINPUT91), .A4(new_n580), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n608), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n588), .A2(new_n576), .A3(new_n589), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n575), .B1(new_n533), .B2(new_n537), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n579), .A2(new_n395), .A3(new_n580), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n406), .A2(new_n405), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n628), .B(new_n583), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT35), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n626), .A2(new_n627), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n301), .B1(new_n591), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n407), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n272), .A2(KEYINPUT17), .ZN(new_n636));
  XNOR2_X1  g435(.A(G99gat), .B(G106gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(KEYINPUT107), .ZN(new_n638));
  INV_X1    g437(.A(G99gat), .ZN(new_n639));
  INV_X1    g438(.A(G106gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT107), .ZN(new_n642));
  NAND2_X1  g441(.A1(G99gat), .A2(G106gat), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n638), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(KEYINPUT106), .A2(G85gat), .A3(G92gat), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT7), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g447(.A1(KEYINPUT106), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n643), .A2(KEYINPUT8), .ZN(new_n650));
  INV_X1    g449(.A(G85gat), .ZN(new_n651));
  INV_X1    g450(.A(G92gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n648), .A2(new_n649), .A3(new_n650), .A4(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n645), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n645), .A2(new_n654), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n636), .B(new_n236), .C1(new_n655), .C2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n655), .ZN(new_n659));
  AND2_X1   g458(.A1(G232gat), .A2(G233gat), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n231), .A2(new_n659), .B1(KEYINPUT41), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(G190gat), .B(G218gat), .Z(new_n663));
  AND2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  XOR2_X1   g464(.A(G134gat), .B(G162gat), .Z(new_n666));
  NOR2_X1   g465(.A1(new_n660), .A2(KEYINPUT41), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  OR4_X1    g467(.A1(KEYINPUT108), .A2(new_n664), .A3(new_n665), .A4(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n668), .B(KEYINPUT108), .Z(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(new_n664), .B2(new_n665), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(G71gat), .A2(G78gat), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT9), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n673), .B1(new_n674), .B2(KEYINPUT104), .ZN(new_n675));
  NOR2_X1   g474(.A1(G71gat), .A2(G78gat), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(G57gat), .A2(G64gat), .ZN(new_n678));
  NOR2_X1   g477(.A1(G57gat), .A2(G64gat), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n677), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n681), .A2(new_n678), .A3(new_n679), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n683), .B1(new_n676), .B2(new_n675), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT21), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(G231gat), .A2(G233gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(G127gat), .B(G155gat), .Z(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n689), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(G183gat), .B(G211gat), .Z(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n692), .B(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n685), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT21), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n286), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT105), .B(KEYINPUT19), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n695), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(G230gat), .A2(G233gat), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n685), .B1(new_n657), .B2(new_n655), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n638), .A2(new_n644), .ZN(new_n705));
  INV_X1    g504(.A(new_n654), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n707), .A2(new_n684), .A3(new_n682), .A4(new_n656), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT10), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n704), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n659), .A2(KEYINPUT10), .A3(new_n696), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n703), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n702), .B1(new_n704), .B2(new_n708), .ZN(new_n713));
  XNOR2_X1  g512(.A(G120gat), .B(G148gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT109), .ZN(new_n715));
  XNOR2_X1  g514(.A(G176gat), .B(G204gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n712), .A2(new_n713), .A3(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n702), .B(KEYINPUT110), .Z(new_n720));
  AOI21_X1  g519(.A(new_n720), .B1(new_n710), .B2(new_n711), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n717), .B1(new_n721), .B2(new_n713), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n672), .A2(new_n701), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n634), .A2(new_n635), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g526(.A1(new_n634), .A2(new_n725), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(KEYINPUT16), .B(G8gat), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n729), .A2(new_n496), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n237), .B1(new_n728), .B2(new_n495), .ZN(new_n732));
  OAI21_X1  g531(.A(KEYINPUT42), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(KEYINPUT42), .B2(new_n731), .ZN(G1325gat));
  AND2_X1   g533(.A1(new_n588), .A2(new_n589), .ZN(new_n735));
  OAI21_X1  g534(.A(G15gat), .B1(new_n729), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n728), .A2(new_n238), .A3(new_n538), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(G1326gat));
  NAND2_X1  g537(.A1(new_n728), .A2(new_n575), .ZN(new_n739));
  XNOR2_X1  g538(.A(KEYINPUT43), .B(G22gat), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1327gat));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n591), .A2(new_n633), .ZN(new_n743));
  INV_X1    g542(.A(new_n672), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n701), .A2(new_n723), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(new_n301), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n407), .A2(G29gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT111), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n752), .A2(KEYINPUT111), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n742), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n752), .A2(KEYINPUT111), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n757), .A2(KEYINPUT45), .A3(new_n753), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n743), .A2(KEYINPUT44), .A3(new_n744), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT44), .B1(new_n743), .B2(new_n744), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n759), .A2(new_n760), .A3(new_n749), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(G29gat), .B1(new_n762), .B2(new_n407), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n756), .A2(new_n758), .A3(new_n763), .ZN(G1328gat));
  OAI21_X1  g563(.A(G36gat), .B1(new_n762), .B2(new_n496), .ZN(new_n765));
  NOR4_X1   g564(.A1(new_n745), .A2(G36gat), .A3(new_n496), .A4(new_n749), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT46), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1329gat));
  AND3_X1   g567(.A1(new_n750), .A2(new_n208), .A3(new_n538), .ZN(new_n769));
  INV_X1    g568(.A(new_n760), .ZN(new_n770));
  INV_X1    g569(.A(new_n735), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n672), .B1(new_n591), .B2(new_n633), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT44), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n770), .A2(new_n771), .A3(new_n748), .A4(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n769), .B1(G43gat), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT47), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT47), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n208), .B1(new_n761), .B2(new_n771), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n769), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n779), .ZN(G1330gat));
  NAND2_X1  g579(.A1(new_n575), .A2(new_n205), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n781), .A2(KEYINPUT112), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(KEYINPUT112), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n747), .A2(new_n672), .ZN(new_n784));
  AND4_X1   g583(.A1(new_n634), .A2(new_n782), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n759), .A2(new_n760), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n786), .A2(new_n575), .A3(new_n748), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n785), .B1(new_n787), .B2(G50gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT48), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT48), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n205), .B1(new_n761), .B2(new_n575), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n791), .B2(new_n785), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(G1331gat));
  INV_X1    g592(.A(new_n203), .ZN(new_n794));
  AOI211_X1 g593(.A(new_n794), .B(new_n262), .C1(new_n280), .C2(new_n281), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT103), .B1(new_n795), .B2(KEYINPUT18), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n274), .A2(new_n202), .A3(new_n275), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n290), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n298), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n284), .A2(new_n290), .A3(new_n296), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n701), .ZN(new_n802));
  NOR4_X1   g601(.A1(new_n801), .A2(new_n744), .A3(new_n802), .A4(new_n724), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT113), .B1(new_n743), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n805));
  INV_X1    g604(.A(new_n803), .ZN(new_n806));
  AOI211_X1 g605(.A(new_n805), .B(new_n806), .C1(new_n591), .C2(new_n633), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n635), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g609(.A(new_n496), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(KEYINPUT114), .Z(new_n812));
  NOR3_X1   g611(.A1(new_n804), .A2(new_n807), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n813), .B(new_n814), .ZN(G1333gat));
  NAND2_X1  g614(.A1(new_n743), .A2(new_n803), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n805), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n743), .A2(KEYINPUT113), .A3(new_n803), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(new_n538), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(G71gat), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n735), .A2(new_n820), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n808), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n823), .ZN(new_n825));
  NOR4_X1   g624(.A1(new_n804), .A2(new_n807), .A3(KEYINPUT115), .A4(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n821), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT50), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n829), .B(new_n821), .C1(new_n824), .C2(new_n826), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(G1334gat));
  NAND2_X1  g630(.A1(new_n808), .A2(new_n575), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g632(.A1(new_n301), .A2(new_n802), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT116), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n723), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n759), .A2(new_n760), .A3(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(G85gat), .B1(new_n838), .B2(new_n407), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n772), .A2(new_n835), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n772), .A2(KEYINPUT51), .A3(new_n835), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n844), .A2(new_n651), .A3(new_n635), .A4(new_n723), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n839), .A2(new_n845), .ZN(G1336gat));
  NOR2_X1   g645(.A1(new_n724), .A2(G92gat), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n844), .A2(new_n495), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n652), .B1(new_n837), .B2(new_n495), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT52), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n844), .A2(new_n495), .A3(new_n847), .ZN(new_n851));
  INV_X1    g650(.A(new_n836), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n770), .A2(new_n495), .A3(new_n773), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(G92gat), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n851), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n850), .A2(new_n856), .ZN(G1337gat));
  OAI21_X1  g656(.A(G99gat), .B1(new_n838), .B2(new_n735), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n844), .A2(new_n639), .A3(new_n538), .A4(new_n723), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1338gat));
  NOR2_X1   g659(.A1(new_n724), .A2(G106gat), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n844), .A2(new_n575), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n640), .B1(new_n837), .B2(new_n575), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT53), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n844), .A2(new_n575), .A3(new_n861), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n770), .A2(new_n575), .A3(new_n773), .A4(new_n852), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(G106gat), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n865), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n864), .A2(new_n869), .ZN(G1339gat));
  NAND2_X1  g669(.A1(new_n725), .A2(new_n301), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT55), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n710), .A2(new_n711), .A3(new_n720), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n875), .A2(new_n712), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n710), .A2(new_n711), .ZN(new_n878));
  INV_X1    g677(.A(new_n720), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n717), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n874), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n878), .A2(new_n702), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n710), .A2(new_n711), .A3(new_n720), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(KEYINPUT54), .A3(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n717), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n886), .B1(new_n721), .B2(new_n876), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n885), .A2(KEYINPUT55), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n882), .A2(new_n719), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT117), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n885), .A2(new_n887), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n718), .B1(new_n891), .B2(new_n874), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n893), .A3(new_n888), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n895), .B1(new_n799), .B2(new_n800), .ZN(new_n896));
  INV_X1    g695(.A(new_n289), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n287), .B(new_n897), .C1(new_n270), .C2(new_n273), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT118), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT118), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n285), .A2(new_n900), .A3(new_n287), .A4(new_n897), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n899), .B(new_n901), .C1(new_n203), .C2(new_n282), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n295), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n800), .A2(new_n903), .A3(new_n723), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n873), .B1(new_n896), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n889), .A2(KEYINPUT117), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n893), .B1(new_n892), .B2(new_n888), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n908), .B1(new_n297), .B2(new_n300), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n800), .A2(new_n903), .A3(new_n723), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(KEYINPUT119), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n905), .A2(new_n672), .A3(new_n911), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n744), .A2(new_n800), .A3(new_n908), .A4(new_n903), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n872), .B1(new_n914), .B2(new_n802), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n915), .A2(new_n577), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n407), .A2(new_n495), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n918), .A2(new_n301), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(new_n307), .ZN(G1340gat));
  NOR2_X1   g719(.A1(new_n918), .A2(new_n724), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(new_n310), .ZN(G1341gat));
  INV_X1    g721(.A(new_n918), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n701), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n317), .A2(KEYINPUT120), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n924), .B(new_n925), .ZN(G1342gat));
  AOI21_X1  g725(.A(new_n672), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  OR2_X1    g727(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n928), .B(new_n929), .ZN(G1343gat));
  INV_X1    g729(.A(G141gat), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n735), .A2(new_n917), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n701), .B1(new_n912), .B2(new_n913), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n575), .B1(new_n933), .B2(new_n872), .ZN(new_n934));
  XOR2_X1   g733(.A(KEYINPUT121), .B(KEYINPUT57), .Z(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n889), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n801), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n744), .B1(new_n938), .B2(new_n910), .ZN(new_n939));
  INV_X1    g738(.A(new_n913), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n802), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n871), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT57), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n576), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n932), .B1(new_n936), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n931), .B1(new_n946), .B2(new_n801), .ZN(new_n947));
  INV_X1    g746(.A(new_n934), .ZN(new_n948));
  INV_X1    g747(.A(new_n932), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n801), .A2(new_n931), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(KEYINPUT58), .B1(new_n947), .B2(new_n952), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n950), .A2(new_n951), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT58), .ZN(new_n955));
  AOI211_X1 g754(.A(new_n301), .B(new_n932), .C1(new_n936), .C2(new_n945), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n954), .B(new_n955), .C1(new_n956), .C2(new_n931), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n953), .A2(new_n957), .ZN(G1344gat));
  INV_X1    g757(.A(new_n950), .ZN(new_n959));
  INV_X1    g758(.A(G148gat), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(new_n960), .A3(new_n723), .ZN(new_n961));
  AOI211_X1 g760(.A(KEYINPUT59), .B(new_n960), .C1(new_n946), .C2(new_n723), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT59), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n909), .A2(new_n910), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n744), .B1(new_n964), .B2(new_n873), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n940), .B1(new_n965), .B2(new_n911), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n871), .B1(new_n966), .B2(new_n701), .ZN(new_n967));
  INV_X1    g766(.A(new_n935), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n967), .A2(new_n575), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n938), .A2(new_n910), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(new_n672), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n744), .A2(new_n800), .A3(new_n903), .A4(new_n937), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n701), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT122), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n871), .B(new_n974), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n575), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(new_n943), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n969), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n978), .A2(new_n723), .A3(new_n949), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n963), .B1(new_n979), .B2(G148gat), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n961), .B1(new_n962), .B2(new_n980), .ZN(G1345gat));
  INV_X1    g780(.A(new_n946), .ZN(new_n982));
  OAI21_X1  g781(.A(G155gat), .B1(new_n982), .B2(new_n802), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n959), .A2(new_n341), .A3(new_n701), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(G1346gat));
  OAI21_X1  g784(.A(G162gat), .B1(new_n982), .B2(new_n672), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n672), .A2(G162gat), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT123), .B1(new_n959), .B2(new_n987), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n959), .A2(KEYINPUT123), .A3(new_n987), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(G1347gat));
  NOR2_X1   g789(.A1(new_n635), .A2(new_n496), .ZN(new_n991));
  OAI211_X1 g790(.A(new_n991), .B(new_n628), .C1(new_n933), .C2(new_n872), .ZN(new_n992));
  INV_X1    g791(.A(G169gat), .ZN(new_n993));
  NOR3_X1   g792(.A1(new_n992), .A2(new_n993), .A3(new_n301), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT124), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n995), .B1(new_n915), .B2(new_n635), .ZN(new_n996));
  OAI211_X1 g795(.A(KEYINPUT124), .B(new_n407), .C1(new_n933), .C2(new_n872), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n577), .A2(new_n496), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n998), .A2(new_n801), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g799(.A(new_n994), .B1(new_n1000), .B2(new_n993), .ZN(G1348gat));
  OAI21_X1  g800(.A(G176gat), .B1(new_n992), .B2(new_n724), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n998), .A2(new_n999), .ZN(new_n1003));
  OR2_X1    g802(.A1(new_n724), .A2(G176gat), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(G1349gat));
  NAND4_X1  g804(.A1(new_n916), .A2(KEYINPUT125), .A3(new_n701), .A4(new_n991), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT125), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1007), .B1(new_n992), .B2(new_n802), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1006), .A2(G183gat), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g808(.A1(new_n802), .A2(new_n454), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n998), .A2(new_n999), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1012), .A2(KEYINPUT60), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT60), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n1009), .A2(new_n1011), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1013), .A2(new_n1015), .ZN(G1350gat));
  OAI21_X1  g815(.A(G190gat), .B1(new_n992), .B2(new_n672), .ZN(new_n1017));
  XNOR2_X1  g816(.A(new_n1017), .B(KEYINPUT61), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n744), .A2(new_n441), .ZN(new_n1019));
  OAI21_X1  g818(.A(new_n1018), .B1(new_n1003), .B2(new_n1019), .ZN(G1351gat));
  NAND2_X1  g819(.A1(new_n991), .A2(new_n735), .ZN(new_n1021));
  AOI21_X1  g820(.A(new_n1021), .B1(new_n969), .B2(new_n977), .ZN(new_n1022));
  INV_X1    g821(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g822(.A(G197gat), .B1(new_n1023), .B2(new_n301), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n590), .A2(new_n495), .ZN(new_n1025));
  AOI21_X1  g824(.A(new_n1025), .B1(new_n996), .B2(new_n997), .ZN(new_n1026));
  INV_X1    g825(.A(KEYINPUT126), .ZN(new_n1027));
  NOR2_X1   g826(.A1(new_n301), .A2(G197gat), .ZN(new_n1028));
  AND3_X1   g827(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g828(.A(new_n1027), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1030));
  OAI21_X1  g829(.A(new_n1024), .B1(new_n1029), .B2(new_n1030), .ZN(G1352gat));
  INV_X1    g830(.A(KEYINPUT62), .ZN(new_n1032));
  INV_X1    g831(.A(KEYINPUT127), .ZN(new_n1033));
  INV_X1    g832(.A(new_n1025), .ZN(new_n1034));
  NOR2_X1   g833(.A1(new_n724), .A2(G204gat), .ZN(new_n1035));
  NAND2_X1  g834(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g835(.A(new_n1036), .ZN(new_n1037));
  AOI21_X1  g836(.A(new_n1033), .B1(new_n998), .B2(new_n1037), .ZN(new_n1038));
  AOI211_X1 g837(.A(KEYINPUT127), .B(new_n1036), .C1(new_n996), .C2(new_n997), .ZN(new_n1039));
  OAI21_X1  g838(.A(new_n1032), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g839(.A(KEYINPUT124), .B1(new_n967), .B2(new_n407), .ZN(new_n1041));
  INV_X1    g840(.A(new_n997), .ZN(new_n1042));
  OAI21_X1  g841(.A(new_n1037), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g842(.A1(new_n1043), .A2(KEYINPUT127), .ZN(new_n1044));
  NAND3_X1  g843(.A1(new_n998), .A2(new_n1033), .A3(new_n1037), .ZN(new_n1045));
  NAND3_X1  g844(.A1(new_n1044), .A2(KEYINPUT62), .A3(new_n1045), .ZN(new_n1046));
  OAI21_X1  g845(.A(G204gat), .B1(new_n1023), .B2(new_n724), .ZN(new_n1047));
  NAND3_X1  g846(.A1(new_n1040), .A2(new_n1046), .A3(new_n1047), .ZN(G1353gat));
  NAND3_X1  g847(.A1(new_n1026), .A2(new_n466), .A3(new_n701), .ZN(new_n1049));
  INV_X1    g848(.A(KEYINPUT63), .ZN(new_n1050));
  INV_X1    g849(.A(G211gat), .ZN(new_n1051));
  AOI211_X1 g850(.A(new_n1050), .B(new_n1051), .C1(new_n1022), .C2(new_n701), .ZN(new_n1052));
  INV_X1    g851(.A(new_n1021), .ZN(new_n1053));
  NAND3_X1  g852(.A1(new_n978), .A2(new_n701), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g853(.A(KEYINPUT63), .B1(new_n1054), .B2(G211gat), .ZN(new_n1055));
  OAI21_X1  g854(.A(new_n1049), .B1(new_n1052), .B2(new_n1055), .ZN(G1354gat));
  OAI21_X1  g855(.A(G218gat), .B1(new_n1023), .B2(new_n672), .ZN(new_n1057));
  NAND3_X1  g856(.A1(new_n1026), .A2(new_n467), .A3(new_n744), .ZN(new_n1058));
  NAND2_X1  g857(.A1(new_n1057), .A2(new_n1058), .ZN(G1355gat));
endmodule


