

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769;

  NOR2_X2 U373 ( .A1(n400), .A2(n396), .ZN(n419) );
  OR2_X2 U374 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X2 U375 ( .A(n509), .B(n355), .ZN(n612) );
  NOR2_X2 U376 ( .A1(n658), .A2(G902), .ZN(n549) );
  NOR2_X2 U377 ( .A1(n717), .A2(n716), .ZN(n630) );
  NAND2_X1 U378 ( .A1(n691), .A2(n483), .ZN(n466) );
  XNOR2_X1 U379 ( .A(n438), .B(KEYINPUT73), .ZN(n634) );
  AND2_X1 U380 ( .A1(n466), .A2(G472), .ZN(n394) );
  OR2_X1 U381 ( .A1(n418), .A2(n642), .ZN(n643) );
  NAND2_X1 U382 ( .A1(n429), .A2(n634), .ZN(n437) );
  XNOR2_X1 U383 ( .A(n700), .B(n550), .ZN(n615) );
  NOR2_X1 U384 ( .A1(n600), .A2(n640), .ZN(n601) );
  XNOR2_X1 U385 ( .A(G478), .B(n527), .ZN(n586) );
  XNOR2_X1 U386 ( .A(G131), .B(KEYINPUT69), .ZN(n488) );
  XNOR2_X1 U387 ( .A(n556), .B(n557), .ZN(n736) );
  XNOR2_X2 U388 ( .A(n549), .B(G472), .ZN(n600) );
  INV_X1 U389 ( .A(n615), .ZN(n637) );
  INV_X1 U390 ( .A(n589), .ZN(n389) );
  NOR2_X1 U391 ( .A1(n617), .A2(n403), .ZN(n402) );
  XNOR2_X1 U392 ( .A(n685), .B(KEYINPUT81), .ZN(n617) );
  NAND2_X1 U393 ( .A1(n619), .A2(n404), .ZN(n403) );
  INV_X1 U394 ( .A(KEYINPUT79), .ZN(n373) );
  NOR2_X1 U395 ( .A1(n613), .A2(n697), .ZN(n423) );
  NOR2_X1 U396 ( .A1(n581), .A2(n637), .ZN(n582) );
  XNOR2_X1 U397 ( .A(KEYINPUT71), .B(G469), .ZN(n481) );
  XNOR2_X1 U398 ( .A(n421), .B(n420), .ZN(n562) );
  INV_X1 U399 ( .A(KEYINPUT8), .ZN(n420) );
  NOR2_X1 U400 ( .A1(n465), .A2(n648), .ZN(n464) );
  INV_X1 U401 ( .A(KEYINPUT22), .ZN(n405) );
  AND2_X2 U402 ( .A1(n386), .A2(n466), .ZN(n395) );
  XOR2_X1 U403 ( .A(KEYINPUT101), .B(KEYINPUT7), .Z(n521) );
  XNOR2_X1 U404 ( .A(G107), .B(KEYINPUT9), .ZN(n520) );
  NOR2_X1 U405 ( .A1(n671), .A2(n766), .ZN(n595) );
  OR2_X1 U406 ( .A1(G902), .A2(G237), .ZN(n507) );
  XNOR2_X1 U407 ( .A(n457), .B(G146), .ZN(n500) );
  INV_X1 U408 ( .A(G125), .ZN(n457) );
  NOR2_X1 U409 ( .A1(G953), .A2(G237), .ZN(n547) );
  XNOR2_X1 U410 ( .A(n445), .B(n444), .ZN(n487) );
  XNOR2_X1 U411 ( .A(n486), .B(n484), .ZN(n444) );
  XNOR2_X1 U412 ( .A(n485), .B(n446), .ZN(n445) );
  XNOR2_X1 U413 ( .A(KEYINPUT15), .B(G902), .ZN(n649) );
  XNOR2_X1 U414 ( .A(n419), .B(n636), .ZN(n376) );
  NAND2_X1 U415 ( .A1(n374), .A2(n373), .ZN(n368) );
  XOR2_X1 U416 ( .A(KEYINPUT75), .B(n607), .Z(n613) );
  XNOR2_X1 U417 ( .A(n449), .B(n447), .ZN(n585) );
  XNOR2_X1 U418 ( .A(n529), .B(n448), .ZN(n447) );
  OR2_X1 U419 ( .A1(n528), .A2(G902), .ZN(n449) );
  INV_X1 U420 ( .A(G475), .ZN(n448) );
  XNOR2_X1 U421 ( .A(n500), .B(n367), .ZN(n751) );
  XNOR2_X1 U422 ( .A(G140), .B(KEYINPUT10), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n560), .B(n366), .ZN(n365) );
  XNOR2_X1 U424 ( .A(G128), .B(G110), .ZN(n560) );
  XNOR2_X1 U425 ( .A(G119), .B(G137), .ZN(n366) );
  XNOR2_X1 U426 ( .A(n422), .B(n561), .ZN(n364) );
  INV_X1 U427 ( .A(KEYINPUT24), .ZN(n561) );
  XNOR2_X1 U428 ( .A(KEYINPUT23), .B(KEYINPUT92), .ZN(n422) );
  XNOR2_X1 U429 ( .A(n408), .B(n525), .ZN(n653) );
  XNOR2_X1 U430 ( .A(n526), .B(n426), .ZN(n408) );
  INV_X1 U431 ( .A(n542), .ZN(n426) );
  XNOR2_X1 U432 ( .A(n496), .B(n495), .ZN(n554) );
  INV_X1 U433 ( .A(G110), .ZN(n495) );
  XNOR2_X1 U434 ( .A(G107), .B(G104), .ZN(n496) );
  INV_X1 U435 ( .A(G146), .ZN(n546) );
  AND2_X1 U436 ( .A1(n455), .A2(n678), .ZN(n614) );
  NAND2_X1 U437 ( .A1(n612), .A2(n415), .ZN(n393) );
  XNOR2_X1 U438 ( .A(n624), .B(n625), .ZN(n631) );
  BUF_X1 U439 ( .A(n702), .Z(n418) );
  INV_X1 U440 ( .A(KEYINPUT84), .ZN(n559) );
  AND2_X1 U441 ( .A1(n392), .A2(n391), .ZN(n390) );
  NOR2_X1 U442 ( .A1(n551), .A2(KEYINPUT83), .ZN(n388) );
  NOR2_X1 U443 ( .A1(n473), .A2(n559), .ZN(n470) );
  INV_X1 U444 ( .A(KEYINPUT120), .ZN(n380) );
  NOR2_X1 U445 ( .A1(n729), .A2(n730), .ZN(n381) );
  NOR2_X1 U446 ( .A1(n695), .A2(G953), .ZN(n378) );
  AND2_X2 U447 ( .A1(n745), .A2(n463), .ZN(n456) );
  INV_X1 U448 ( .A(KEYINPUT2), .ZN(n467) );
  XNOR2_X1 U449 ( .A(n417), .B(n416), .ZN(n767) );
  INV_X1 U450 ( .A(KEYINPUT40), .ZN(n416) );
  XOR2_X1 U451 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n485) );
  XNOR2_X1 U452 ( .A(G143), .B(G104), .ZN(n446) );
  XNOR2_X1 U453 ( .A(G122), .B(G113), .ZN(n486) );
  XNOR2_X1 U454 ( .A(n479), .B(G137), .ZN(n478) );
  INV_X1 U455 ( .A(KEYINPUT70), .ZN(n479) );
  XNOR2_X1 U456 ( .A(n498), .B(n499), .ZN(n502) );
  XOR2_X1 U457 ( .A(KEYINPUT18), .B(KEYINPUT87), .Z(n499) );
  XNOR2_X1 U458 ( .A(n397), .B(KEYINPUT46), .ZN(n396) );
  XOR2_X1 U459 ( .A(KEYINPUT93), .B(KEYINPUT20), .Z(n531) );
  XNOR2_X1 U460 ( .A(n548), .B(n538), .ZN(n443) );
  XNOR2_X1 U461 ( .A(n414), .B(n497), .ZN(n537) );
  XNOR2_X1 U462 ( .A(n412), .B(G119), .ZN(n414) );
  XNOR2_X1 U463 ( .A(KEYINPUT3), .B(G101), .ZN(n412) );
  XNOR2_X1 U464 ( .A(G134), .B(n518), .ZN(n542) );
  XNOR2_X1 U465 ( .A(G116), .B(G122), .ZN(n519) );
  XNOR2_X1 U466 ( .A(n595), .B(n361), .ZN(n360) );
  INV_X1 U467 ( .A(KEYINPUT44), .ZN(n361) );
  XNOR2_X1 U468 ( .A(KEYINPUT38), .B(n644), .ZN(n714) );
  AND2_X1 U469 ( .A1(n702), .A2(n409), .ZN(n571) );
  NAND2_X1 U470 ( .A1(n732), .A2(n649), .ZN(n509) );
  NAND2_X1 U471 ( .A1(n551), .A2(KEYINPUT83), .ZN(n391) );
  XNOR2_X1 U472 ( .A(n556), .B(n441), .ZN(n658) );
  XNOR2_X1 U473 ( .A(n537), .B(n442), .ZN(n441) );
  XNOR2_X1 U474 ( .A(n443), .B(n536), .ZN(n442) );
  XOR2_X1 U475 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n536) );
  XNOR2_X1 U476 ( .A(n458), .B(G953), .ZN(n524) );
  INV_X1 U477 ( .A(KEYINPUT64), .ZN(n458) );
  XNOR2_X1 U478 ( .A(n537), .B(n459), .ZN(n504) );
  XNOR2_X1 U479 ( .A(n554), .B(n460), .ZN(n459) );
  XNOR2_X1 U480 ( .A(KEYINPUT16), .B(G122), .ZN(n460) );
  XNOR2_X1 U481 ( .A(n491), .B(n490), .ZN(n528) );
  NAND2_X1 U482 ( .A1(n371), .A2(n373), .ZN(n370) );
  AND2_X1 U483 ( .A1(n369), .A2(n353), .ZN(n372) );
  NOR2_X1 U484 ( .A1(n639), .A2(n640), .ZN(n641) );
  XNOR2_X1 U485 ( .A(n475), .B(KEYINPUT35), .ZN(n765) );
  INV_X1 U486 ( .A(n613), .ZN(n439) );
  BUF_X1 U487 ( .A(n700), .Z(n410) );
  BUF_X1 U488 ( .A(n572), .Z(n583) );
  XNOR2_X1 U489 ( .A(n751), .B(n363), .ZN(n564) );
  XNOR2_X1 U490 ( .A(n365), .B(n364), .ZN(n363) );
  XOR2_X1 U491 ( .A(G101), .B(G140), .Z(n553) );
  OR2_X1 U492 ( .A1(n424), .A2(n473), .ZN(n685) );
  INV_X1 U493 ( .A(KEYINPUT36), .ZN(n425) );
  AND2_X1 U494 ( .A1(n615), .A2(n614), .ZN(n616) );
  BUF_X1 U495 ( .A(n765), .Z(n407) );
  NAND2_X1 U496 ( .A1(n351), .A2(n593), .ZN(n594) );
  XNOR2_X1 U497 ( .A(n384), .B(KEYINPUT74), .ZN(n676) );
  NOR2_X1 U498 ( .A1(n631), .A2(n626), .ZN(n384) );
  INV_X1 U499 ( .A(KEYINPUT102), .ZN(n453) );
  NOR2_X1 U500 ( .A1(n470), .A2(n696), .ZN(n469) );
  INV_X1 U501 ( .A(KEYINPUT122), .ZN(n427) );
  INV_X1 U502 ( .A(KEYINPUT60), .ZN(n433) );
  NAND2_X1 U503 ( .A1(n435), .A2(n656), .ZN(n434) );
  XNOR2_X1 U504 ( .A(n436), .B(n358), .ZN(n435) );
  INV_X1 U505 ( .A(KEYINPUT56), .ZN(n431) );
  OR2_X1 U506 ( .A1(n693), .A2(n456), .ZN(n382) );
  AND2_X1 U507 ( .A1(n379), .A2(n378), .ZN(n377) );
  XOR2_X1 U508 ( .A(KEYINPUT90), .B(n494), .Z(n640) );
  INV_X1 U509 ( .A(n640), .ZN(n415) );
  AND2_X1 U510 ( .A1(n389), .A2(n637), .ZN(n351) );
  XNOR2_X1 U511 ( .A(n539), .B(n503), .ZN(n352) );
  AND2_X1 U512 ( .A1(n368), .A2(n689), .ZN(n353) );
  AND2_X1 U513 ( .A1(n466), .A2(G475), .ZN(n354) );
  XOR2_X1 U514 ( .A(n508), .B(n510), .Z(n355) );
  AND2_X1 U515 ( .A1(n473), .A2(n559), .ZN(n356) );
  AND2_X1 U516 ( .A1(n382), .A2(n377), .ZN(n357) );
  XOR2_X1 U517 ( .A(n493), .B(n492), .Z(n358) );
  NOR2_X1 U518 ( .A1(n755), .A2(G952), .ZN(n740) );
  XNOR2_X1 U519 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n359) );
  INV_X1 U520 ( .A(n690), .ZN(n374) );
  NOR2_X2 U521 ( .A1(n572), .A2(n535), .ZN(n406) );
  NAND2_X1 U522 ( .A1(n360), .A2(n596), .ZN(n597) );
  AND2_X1 U523 ( .A1(n633), .A2(n714), .ZN(n429) );
  XNOR2_X1 U524 ( .A(n601), .B(KEYINPUT30), .ZN(n633) );
  XNOR2_X2 U525 ( .A(n599), .B(KEYINPUT45), .ZN(n745) );
  NAND2_X1 U526 ( .A1(n362), .A2(n588), .ZN(n430) );
  XNOR2_X1 U527 ( .A(n587), .B(KEYINPUT86), .ZN(n362) );
  NAND2_X1 U528 ( .A1(n376), .A2(n375), .ZN(n369) );
  NAND2_X2 U529 ( .A1(n372), .A2(n370), .ZN(n652) );
  INV_X1 U530 ( .A(n376), .ZN(n371) );
  AND2_X1 U531 ( .A1(n690), .A2(KEYINPUT79), .ZN(n375) );
  XNOR2_X1 U532 ( .A(n381), .B(n380), .ZN(n379) );
  NAND2_X1 U533 ( .A1(n383), .A2(n628), .ZN(n401) );
  XNOR2_X1 U534 ( .A(n676), .B(n627), .ZN(n383) );
  NAND2_X1 U535 ( .A1(n385), .A2(n742), .ZN(n506) );
  INV_X1 U536 ( .A(n461), .ZN(n385) );
  XNOR2_X1 U537 ( .A(n462), .B(n352), .ZN(n461) );
  NAND2_X1 U538 ( .A1(n394), .A2(n386), .ZN(n660) );
  NAND2_X1 U539 ( .A1(n354), .A2(n386), .ZN(n436) );
  NOR2_X4 U540 ( .A1(n456), .A2(n464), .ZN(n386) );
  NAND2_X1 U541 ( .A1(n390), .A2(n387), .ZN(n474) );
  NAND2_X1 U542 ( .A1(n389), .A2(n388), .ZN(n387) );
  NAND2_X1 U543 ( .A1(n589), .A2(KEYINPUT83), .ZN(n392) );
  INV_X1 U544 ( .A(n517), .ZN(n626) );
  XNOR2_X2 U545 ( .A(n393), .B(KEYINPUT19), .ZN(n517) );
  NAND2_X1 U546 ( .A1(n395), .A2(G210), .ZN(n734) );
  NAND2_X1 U547 ( .A1(n395), .A2(G478), .ZN(n655) );
  NAND2_X1 U548 ( .A1(n395), .A2(G469), .ZN(n452) );
  NAND2_X1 U549 ( .A1(n395), .A2(G217), .ZN(n737) );
  NAND2_X1 U550 ( .A1(n399), .A2(n398), .ZN(n397) );
  INV_X1 U551 ( .A(n769), .ZN(n398) );
  INV_X1 U552 ( .A(n767), .ZN(n399) );
  NAND2_X1 U553 ( .A1(n401), .A2(n402), .ZN(n400) );
  INV_X1 U554 ( .A(n675), .ZN(n404) );
  XNOR2_X2 U555 ( .A(n406), .B(n405), .ZN(n589) );
  INV_X1 U556 ( .A(n600), .ZN(n700) );
  NAND2_X1 U557 ( .A1(n423), .A2(n696), .ZN(n638) );
  INV_X2 U558 ( .A(KEYINPUT4), .ZN(n480) );
  NAND2_X1 U559 ( .A1(n517), .A2(n516), .ZN(n413) );
  XNOR2_X1 U560 ( .A(n413), .B(KEYINPUT0), .ZN(n572) );
  NAND2_X1 U561 ( .A1(n440), .A2(n439), .ZN(n438) );
  NAND2_X1 U562 ( .A1(n755), .A2(G234), .ZN(n421) );
  XNOR2_X1 U563 ( .A(n616), .B(n425), .ZN(n424) );
  INV_X1 U564 ( .A(n696), .ZN(n409) );
  XNOR2_X1 U565 ( .A(n622), .B(KEYINPUT1), .ZN(n702) );
  XNOR2_X1 U566 ( .A(n502), .B(n411), .ZN(n462) );
  XNOR2_X1 U567 ( .A(n500), .B(n501), .ZN(n411) );
  INV_X1 U568 ( .A(n612), .ZN(n644) );
  NOR2_X1 U569 ( .A1(n600), .A2(n638), .ZN(n621) );
  NAND2_X1 U570 ( .A1(n646), .A2(n678), .ZN(n417) );
  XNOR2_X2 U571 ( .A(n477), .B(n546), .ZN(n556) );
  NOR2_X1 U572 ( .A1(n697), .A2(n696), .ZN(n703) );
  NOR2_X2 U573 ( .A1(n736), .A2(G902), .ZN(n558) );
  INV_X1 U574 ( .A(n418), .ZN(n473) );
  XNOR2_X1 U575 ( .A(n428), .B(n427), .ZN(G63) );
  NAND2_X1 U576 ( .A1(n657), .A2(n656), .ZN(n428) );
  XNOR2_X1 U577 ( .A(n539), .B(n478), .ZN(n541) );
  XNOR2_X1 U578 ( .A(n430), .B(KEYINPUT85), .ZN(n598) );
  XNOR2_X1 U579 ( .A(n432), .B(n431), .ZN(G51) );
  NAND2_X1 U580 ( .A1(n735), .A2(n656), .ZN(n432) );
  NAND2_X2 U581 ( .A1(n544), .A2(n545), .ZN(n477) );
  XNOR2_X1 U582 ( .A(n434), .B(n433), .ZN(G60) );
  XNOR2_X2 U583 ( .A(n437), .B(n635), .ZN(n646) );
  INV_X1 U584 ( .A(n608), .ZN(n440) );
  NAND2_X1 U585 ( .A1(n754), .A2(n745), .ZN(n691) );
  XNOR2_X2 U586 ( .A(n652), .B(n647), .ZN(n754) );
  AND2_X1 U587 ( .A1(n450), .A2(n656), .ZN(G54) );
  XNOR2_X1 U588 ( .A(n452), .B(n451), .ZN(n450) );
  XNOR2_X1 U589 ( .A(n736), .B(n359), .ZN(n451) );
  XNOR2_X2 U590 ( .A(n454), .B(n453), .ZN(n678) );
  NAND2_X1 U591 ( .A1(n570), .A2(n586), .ZN(n454) );
  AND2_X1 U592 ( .A1(n612), .A2(n482), .ZN(n455) );
  NAND2_X1 U593 ( .A1(n524), .A2(G224), .ZN(n498) );
  NAND2_X1 U594 ( .A1(n461), .A2(n504), .ZN(n505) );
  NOR2_X1 U595 ( .A1(n652), .A2(n467), .ZN(n463) );
  INV_X1 U596 ( .A(n483), .ZN(n465) );
  NOR2_X1 U597 ( .A1(n472), .A2(n468), .ZN(n664) );
  NAND2_X1 U598 ( .A1(n471), .A2(n469), .ZN(n468) );
  NAND2_X1 U599 ( .A1(n474), .A2(n356), .ZN(n471) );
  NOR2_X1 U600 ( .A1(n474), .A2(n559), .ZN(n472) );
  NAND2_X1 U601 ( .A1(n765), .A2(KEYINPUT44), .ZN(n587) );
  NAND2_X1 U602 ( .A1(n476), .A2(n609), .ZN(n475) );
  XNOR2_X1 U603 ( .A(n584), .B(KEYINPUT34), .ZN(n476) );
  XNOR2_X1 U604 ( .A(n477), .B(n752), .ZN(n757) );
  XNOR2_X2 U605 ( .A(n480), .B(KEYINPUT65), .ZN(n539) );
  XNOR2_X2 U606 ( .A(n558), .B(n481), .ZN(n622) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n543) );
  NOR2_X1 U608 ( .A1(n638), .A2(n640), .ZN(n482) );
  XOR2_X1 U609 ( .A(n651), .B(KEYINPUT67), .Z(n483) );
  INV_X1 U610 ( .A(KEYINPUT72), .ZN(n538) );
  XNOR2_X1 U611 ( .A(KEYINPUT103), .B(KEYINPUT6), .ZN(n550) );
  INV_X1 U612 ( .A(n697), .ZN(n533) );
  INV_X1 U613 ( .A(n649), .ZN(n648) );
  XNOR2_X1 U614 ( .A(n540), .B(n489), .ZN(n490) );
  INV_X1 U615 ( .A(KEYINPUT78), .ZN(n647) );
  INV_X1 U616 ( .A(n740), .ZN(n656) );
  INV_X1 U617 ( .A(n685), .ZN(n686) );
  INV_X1 U618 ( .A(KEYINPUT63), .ZN(n662) );
  XNOR2_X1 U619 ( .A(KEYINPUT121), .B(KEYINPUT66), .ZN(n493) );
  INV_X1 U620 ( .A(KEYINPUT11), .ZN(n484) );
  XNOR2_X1 U621 ( .A(n751), .B(n487), .ZN(n491) );
  XNOR2_X1 U622 ( .A(n488), .B(KEYINPUT68), .ZN(n540) );
  AND2_X1 U623 ( .A1(n547), .A2(G214), .ZN(n489) );
  XNOR2_X1 U624 ( .A(n528), .B(KEYINPUT59), .ZN(n492) );
  NAND2_X1 U625 ( .A1(G214), .A2(n507), .ZN(n494) );
  INV_X1 U626 ( .A(KEYINPUT89), .ZN(n510) );
  XNOR2_X1 U627 ( .A(G116), .B(G113), .ZN(n497) );
  INV_X1 U628 ( .A(n504), .ZN(n742) );
  XNOR2_X1 U629 ( .A(KEYINPUT88), .B(KEYINPUT17), .ZN(n501) );
  XNOR2_X1 U630 ( .A(G143), .B(G128), .ZN(n518) );
  INV_X1 U631 ( .A(n518), .ZN(n503) );
  NAND2_X1 U632 ( .A1(n506), .A2(n505), .ZN(n732) );
  NAND2_X1 U633 ( .A1(G210), .A2(n507), .ZN(n508) );
  INV_X1 U634 ( .A(G953), .ZN(n746) );
  NOR2_X1 U635 ( .A1(G898), .A2(n746), .ZN(n741) );
  NAND2_X1 U636 ( .A1(G237), .A2(G234), .ZN(n511) );
  XNOR2_X1 U637 ( .A(n511), .B(KEYINPUT14), .ZN(n513) );
  NAND2_X1 U638 ( .A1(n513), .A2(G902), .ZN(n512) );
  XNOR2_X1 U639 ( .A(n512), .B(KEYINPUT91), .ZN(n602) );
  NAND2_X1 U640 ( .A1(n741), .A2(n602), .ZN(n515) );
  NAND2_X1 U641 ( .A1(G952), .A2(n513), .ZN(n730) );
  NOR2_X1 U642 ( .A1(G953), .A2(n730), .ZN(n606) );
  INV_X1 U643 ( .A(n606), .ZN(n514) );
  NAND2_X1 U644 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U645 ( .A(n519), .B(KEYINPUT100), .ZN(n523) );
  XNOR2_X1 U646 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U647 ( .A(n523), .B(n522), .Z(n526) );
  BUF_X2 U648 ( .A(n524), .Z(n755) );
  NAND2_X1 U649 ( .A1(G217), .A2(n562), .ZN(n525) );
  NOR2_X1 U650 ( .A1(n653), .A2(G902), .ZN(n527) );
  XNOR2_X1 U651 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n529) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n716) );
  INV_X1 U653 ( .A(n716), .ZN(n534) );
  NAND2_X1 U654 ( .A1(G234), .A2(n649), .ZN(n530) );
  XNOR2_X1 U655 ( .A(n531), .B(n530), .ZN(n565) );
  NAND2_X1 U656 ( .A1(n565), .A2(G221), .ZN(n532) );
  XNOR2_X1 U657 ( .A(n532), .B(KEYINPUT21), .ZN(n697) );
  NAND2_X1 U658 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U659 ( .A1(n543), .A2(n542), .ZN(n545) );
  AND2_X1 U660 ( .A1(n547), .A2(G210), .ZN(n548) );
  INV_X1 U661 ( .A(n637), .ZN(n551) );
  NAND2_X1 U662 ( .A1(G227), .A2(n755), .ZN(n552) );
  XNOR2_X1 U663 ( .A(n553), .B(n552), .ZN(n555) );
  XNOR2_X1 U664 ( .A(n555), .B(n554), .ZN(n557) );
  NAND2_X1 U665 ( .A1(G221), .A2(n562), .ZN(n563) );
  XNOR2_X1 U666 ( .A(n564), .B(n563), .ZN(n738) );
  NOR2_X1 U667 ( .A1(n738), .A2(G902), .ZN(n569) );
  XOR2_X1 U668 ( .A(KEYINPUT94), .B(KEYINPUT25), .Z(n567) );
  NAND2_X1 U669 ( .A1(n565), .A2(G217), .ZN(n566) );
  XNOR2_X1 U670 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X2 U671 ( .A(n569), .B(n568), .ZN(n696) );
  INV_X1 U672 ( .A(n585), .ZN(n570) );
  NOR2_X1 U673 ( .A1(n570), .A2(n586), .ZN(n681) );
  NOR2_X1 U674 ( .A1(n681), .A2(n678), .ZN(n718) );
  XOR2_X1 U675 ( .A(KEYINPUT31), .B(KEYINPUT97), .Z(n575) );
  NAND2_X1 U676 ( .A1(n571), .A2(n533), .ZN(n581) );
  NOR2_X1 U677 ( .A1(n600), .A2(n581), .ZN(n709) );
  INV_X1 U678 ( .A(n583), .ZN(n573) );
  NAND2_X1 U679 ( .A1(n709), .A2(n573), .ZN(n574) );
  XNOR2_X1 U680 ( .A(n575), .B(n574), .ZN(n682) );
  NAND2_X1 U681 ( .A1(n622), .A2(n703), .ZN(n608) );
  NOR2_X1 U682 ( .A1(n583), .A2(n608), .ZN(n576) );
  XNOR2_X1 U683 ( .A(n576), .B(KEYINPUT95), .ZN(n577) );
  NOR2_X1 U684 ( .A1(n410), .A2(n577), .ZN(n666) );
  NOR2_X1 U685 ( .A1(n682), .A2(n666), .ZN(n578) );
  NOR2_X1 U686 ( .A1(n718), .A2(n578), .ZN(n579) );
  NOR2_X1 U687 ( .A1(n664), .A2(n579), .ZN(n580) );
  XNOR2_X1 U688 ( .A(n580), .B(KEYINPUT104), .ZN(n588) );
  XNOR2_X1 U689 ( .A(n582), .B(KEYINPUT33), .ZN(n694) );
  NOR2_X1 U690 ( .A1(n583), .A2(n694), .ZN(n584) );
  NOR2_X1 U691 ( .A1(n586), .A2(n585), .ZN(n609) );
  NOR2_X1 U692 ( .A1(n589), .A2(n418), .ZN(n590) );
  NAND2_X1 U693 ( .A1(n590), .A2(n696), .ZN(n591) );
  NOR2_X1 U694 ( .A1(n410), .A2(n591), .ZN(n671) );
  NAND2_X1 U695 ( .A1(n696), .A2(n418), .ZN(n592) );
  XNOR2_X1 U696 ( .A(KEYINPUT105), .B(n592), .ZN(n593) );
  XOR2_X1 U697 ( .A(KEYINPUT32), .B(n594), .Z(n766) );
  NAND2_X1 U698 ( .A1(n595), .A2(n407), .ZN(n596) );
  NAND2_X1 U699 ( .A1(n598), .A2(n597), .ZN(n599) );
  INV_X1 U700 ( .A(n755), .ZN(n603) );
  NAND2_X1 U701 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U702 ( .A1(G900), .A2(n604), .ZN(n605) );
  NOR2_X1 U703 ( .A1(n606), .A2(n605), .ZN(n607) );
  AND2_X1 U704 ( .A1(n633), .A2(n634), .ZN(n610) );
  NAND2_X1 U705 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U706 ( .A1(n644), .A2(n611), .ZN(n675) );
  NAND2_X1 U707 ( .A1(n718), .A2(KEYINPUT47), .ZN(n618) );
  XNOR2_X1 U708 ( .A(n618), .B(KEYINPUT76), .ZN(n619) );
  INV_X1 U709 ( .A(KEYINPUT47), .ZN(n627) );
  INV_X1 U710 ( .A(KEYINPUT107), .ZN(n625) );
  XNOR2_X1 U711 ( .A(KEYINPUT28), .B(KEYINPUT106), .ZN(n620) );
  XNOR2_X1 U712 ( .A(n621), .B(n620), .ZN(n623) );
  NAND2_X1 U713 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U714 ( .A1(n627), .A2(n718), .ZN(n628) );
  NAND2_X1 U715 ( .A1(n714), .A2(n415), .ZN(n717) );
  XNOR2_X1 U716 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n629) );
  XNOR2_X1 U717 ( .A(n630), .B(n629), .ZN(n712) );
  NOR2_X1 U718 ( .A1(n631), .A2(n712), .ZN(n632) );
  XNOR2_X1 U719 ( .A(KEYINPUT42), .B(n632), .ZN(n769) );
  XNOR2_X1 U720 ( .A(KEYINPUT82), .B(KEYINPUT39), .ZN(n635) );
  XNOR2_X1 U721 ( .A(KEYINPUT80), .B(KEYINPUT48), .ZN(n636) );
  OR2_X1 U722 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U723 ( .A1(n641), .A2(n678), .ZN(n642) );
  XNOR2_X1 U724 ( .A(n643), .B(KEYINPUT43), .ZN(n645) );
  NAND2_X1 U725 ( .A1(n645), .A2(n644), .ZN(n690) );
  NAND2_X1 U726 ( .A1(n681), .A2(n646), .ZN(n689) );
  XNOR2_X1 U727 ( .A(KEYINPUT77), .B(n649), .ZN(n650) );
  NAND2_X1 U728 ( .A1(n650), .A2(KEYINPUT2), .ZN(n651) );
  INV_X1 U729 ( .A(n653), .ZN(n654) );
  XNOR2_X1 U730 ( .A(n655), .B(n654), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n658), .B(KEYINPUT62), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n660), .B(n659), .ZN(n661) );
  NOR2_X2 U733 ( .A1(n661), .A2(n740), .ZN(n663) );
  XNOR2_X1 U734 ( .A(n663), .B(n662), .ZN(G57) );
  XOR2_X1 U735 ( .A(n664), .B(G101), .Z(G3) );
  NAND2_X1 U736 ( .A1(n678), .A2(n666), .ZN(n665) );
  XNOR2_X1 U737 ( .A(n665), .B(G104), .ZN(G6) );
  XOR2_X1 U738 ( .A(KEYINPUT109), .B(KEYINPUT27), .Z(n668) );
  NAND2_X1 U739 ( .A1(n666), .A2(n681), .ZN(n667) );
  XNOR2_X1 U740 ( .A(n668), .B(n667), .ZN(n670) );
  XOR2_X1 U741 ( .A(G107), .B(KEYINPUT26), .Z(n669) );
  XNOR2_X1 U742 ( .A(n670), .B(n669), .ZN(G9) );
  XOR2_X1 U743 ( .A(G110), .B(n671), .Z(G12) );
  XOR2_X1 U744 ( .A(KEYINPUT110), .B(KEYINPUT29), .Z(n673) );
  NAND2_X1 U745 ( .A1(n681), .A2(n676), .ZN(n672) );
  XNOR2_X1 U746 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U747 ( .A(G128), .B(n674), .ZN(G30) );
  XOR2_X1 U748 ( .A(G143), .B(n675), .Z(G45) );
  NAND2_X1 U749 ( .A1(n676), .A2(n678), .ZN(n677) );
  XNOR2_X1 U750 ( .A(n677), .B(G146), .ZN(G48) );
  XOR2_X1 U751 ( .A(G113), .B(KEYINPUT111), .Z(n680) );
  NAND2_X1 U752 ( .A1(n682), .A2(n678), .ZN(n679) );
  XNOR2_X1 U753 ( .A(n680), .B(n679), .ZN(G15) );
  NAND2_X1 U754 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U755 ( .A(n683), .B(KEYINPUT112), .ZN(n684) );
  XNOR2_X1 U756 ( .A(G116), .B(n684), .ZN(G18) );
  XOR2_X1 U757 ( .A(KEYINPUT113), .B(KEYINPUT37), .Z(n688) );
  XNOR2_X1 U758 ( .A(G125), .B(n686), .ZN(n687) );
  XNOR2_X1 U759 ( .A(n688), .B(n687), .ZN(G27) );
  XNOR2_X1 U760 ( .A(G134), .B(n689), .ZN(G36) );
  XNOR2_X1 U761 ( .A(G140), .B(n690), .ZN(G42) );
  INV_X1 U762 ( .A(n691), .ZN(n692) );
  NOR2_X1 U763 ( .A1(KEYINPUT2), .A2(n692), .ZN(n693) );
  BUF_X1 U764 ( .A(n694), .Z(n722) );
  NOR2_X1 U765 ( .A1(n712), .A2(n722), .ZN(n695) );
  NAND2_X1 U766 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U767 ( .A(KEYINPUT49), .B(n698), .ZN(n699) );
  NOR2_X1 U768 ( .A1(n410), .A2(n699), .ZN(n701) );
  XOR2_X1 U769 ( .A(KEYINPUT114), .B(n701), .Z(n707) );
  NOR2_X1 U770 ( .A1(n703), .A2(n418), .ZN(n704) );
  XOR2_X1 U771 ( .A(KEYINPUT50), .B(n704), .Z(n705) );
  XNOR2_X1 U772 ( .A(KEYINPUT115), .B(n705), .ZN(n706) );
  NOR2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U774 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U775 ( .A(KEYINPUT51), .B(n710), .Z(n711) );
  NOR2_X1 U776 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U777 ( .A(KEYINPUT116), .B(n713), .ZN(n726) );
  NOR2_X1 U778 ( .A1(n714), .A2(n415), .ZN(n715) );
  NOR2_X1 U779 ( .A1(n716), .A2(n715), .ZN(n721) );
  NOR2_X1 U780 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U781 ( .A(KEYINPUT117), .B(n719), .Z(n720) );
  NOR2_X1 U782 ( .A1(n721), .A2(n720), .ZN(n723) );
  NOR2_X1 U783 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U784 ( .A(KEYINPUT118), .B(n724), .ZN(n725) );
  NOR2_X1 U785 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U786 ( .A(n727), .B(KEYINPUT119), .Z(n728) );
  XNOR2_X1 U787 ( .A(KEYINPUT52), .B(n728), .ZN(n729) );
  XNOR2_X1 U788 ( .A(n357), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U789 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n731) );
  XNOR2_X1 U790 ( .A(n732), .B(n731), .ZN(n733) );
  XNOR2_X1 U791 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U792 ( .A(n738), .B(n737), .ZN(n739) );
  NOR2_X1 U793 ( .A1(n740), .A2(n739), .ZN(G66) );
  NOR2_X1 U794 ( .A1(n742), .A2(n741), .ZN(n750) );
  NAND2_X1 U795 ( .A1(G953), .A2(G224), .ZN(n743) );
  XNOR2_X1 U796 ( .A(KEYINPUT61), .B(n743), .ZN(n744) );
  NAND2_X1 U797 ( .A1(n744), .A2(G898), .ZN(n748) );
  NAND2_X1 U798 ( .A1(n745), .A2(n746), .ZN(n747) );
  NAND2_X1 U799 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U800 ( .A(n750), .B(n749), .ZN(G69) );
  XOR2_X1 U801 ( .A(n751), .B(KEYINPUT123), .Z(n752) );
  INV_X1 U802 ( .A(n757), .ZN(n753) );
  XNOR2_X1 U803 ( .A(n754), .B(n753), .ZN(n756) );
  NAND2_X1 U804 ( .A1(n756), .A2(n755), .ZN(n764) );
  XNOR2_X1 U805 ( .A(n757), .B(KEYINPUT124), .ZN(n758) );
  XNOR2_X1 U806 ( .A(G227), .B(n758), .ZN(n759) );
  NAND2_X1 U807 ( .A1(G900), .A2(n759), .ZN(n760) );
  XOR2_X1 U808 ( .A(KEYINPUT125), .B(n760), .Z(n761) );
  NAND2_X1 U809 ( .A1(G953), .A2(n761), .ZN(n762) );
  XNOR2_X1 U810 ( .A(KEYINPUT126), .B(n762), .ZN(n763) );
  NAND2_X1 U811 ( .A1(n764), .A2(n763), .ZN(G72) );
  XOR2_X1 U812 ( .A(n407), .B(G122), .Z(G24) );
  XOR2_X1 U813 ( .A(G119), .B(n766), .Z(G21) );
  XNOR2_X1 U814 ( .A(G131), .B(KEYINPUT127), .ZN(n768) );
  XNOR2_X1 U815 ( .A(n768), .B(n767), .ZN(G33) );
  XOR2_X1 U816 ( .A(G137), .B(n769), .Z(G39) );
endmodule

