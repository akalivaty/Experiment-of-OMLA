//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n448, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n540, new_n541, new_n542, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n560, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n591, new_n592, new_n594, new_n595, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT64), .Z(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT65), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(new_n455), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2106), .ZN(new_n461));
  INV_X1    g036(.A(new_n457), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G567), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(new_n467), .A3(G2104), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n476), .A2(new_n470), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT66), .B1(new_n469), .B2(KEYINPUT3), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n477), .A2(G137), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n478), .A2(G101), .A3(G2104), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT67), .ZN(new_n482));
  AND3_X1   g057(.A1(new_n474), .A2(new_n480), .A3(new_n482), .ZN(G160));
  NAND4_X1  g058(.A1(new_n479), .A2(new_n476), .A3(G2105), .A4(new_n470), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n478), .A2(G112), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n487));
  OAI22_X1  g062(.A1(new_n484), .A2(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n488), .B1(new_n490), .B2(G136), .ZN(G162));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n479), .A2(new_n476), .A3(new_n470), .A4(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n468), .A2(new_n470), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n492), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n494), .A2(KEYINPUT4), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G114), .C2(new_n478), .ZN(new_n499));
  INV_X1    g074(.A(G126), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n484), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n497), .A2(new_n501), .ZN(G164));
  XNOR2_X1  g077(.A(KEYINPUT6), .B(G651), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT5), .B(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT68), .B(G88), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n503), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n509), .A2(new_n512), .ZN(G166));
  NAND3_X1  g088(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT7), .ZN(new_n515));
  INV_X1    g090(.A(new_n505), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G89), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n518));
  INV_X1    g093(.A(G51), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n507), .B2(new_n519), .ZN(new_n520));
  OAI211_X1 g095(.A(new_n515), .B(new_n517), .C1(new_n520), .C2(KEYINPUT69), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n520), .A2(KEYINPUT69), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(G168));
  NAND2_X1  g098(.A1(new_n516), .A2(G90), .ZN(new_n524));
  INV_X1    g099(.A(new_n507), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G52), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n524), .B(new_n526), .C1(new_n511), .C2(new_n527), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(KEYINPUT70), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(KEYINPUT70), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(G171));
  INV_X1    g106(.A(G81), .ZN(new_n532));
  INV_X1    g107(.A(G43), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n505), .A2(new_n532), .B1(new_n507), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n511), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G860), .ZN(G153));
  NAND4_X1  g113(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g114(.A1(G1), .A2(G3), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT71), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT8), .ZN(new_n542));
  NAND4_X1  g117(.A1(G319), .A2(G483), .A3(G661), .A4(new_n542), .ZN(G188));
  INV_X1    g118(.A(G53), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n544), .B1(new_n545), .B2(KEYINPUT9), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n525), .B(new_n546), .C1(new_n545), .C2(KEYINPUT9), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT9), .ZN(new_n548));
  OAI211_X1 g123(.A(KEYINPUT72), .B(new_n548), .C1(new_n507), .C2(new_n544), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n516), .A2(G91), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  XOR2_X1   g126(.A(KEYINPUT73), .B(G65), .Z(new_n552));
  AOI22_X1  g127(.A1(new_n552), .A2(new_n504), .B1(G78), .B2(G543), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n511), .B1(new_n553), .B2(KEYINPUT74), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n554), .B1(KEYINPUT74), .B2(new_n553), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(G299));
  INV_X1    g131(.A(G171), .ZN(G301));
  INV_X1    g132(.A(G168), .ZN(G286));
  INV_X1    g133(.A(G166), .ZN(G303));
  NAND2_X1  g134(.A1(new_n516), .A2(G87), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n525), .A2(G49), .ZN(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(G288));
  AOI22_X1  g138(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(new_n511), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n516), .A2(G86), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n525), .A2(G48), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G305));
  AOI22_X1  g144(.A1(G85), .A2(new_n516), .B1(new_n525), .B2(G47), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n570), .B(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n573), .A2(new_n511), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(G290));
  AND3_X1   g150(.A1(new_n504), .A2(new_n503), .A3(G92), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT10), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n579), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n504), .A2(G66), .ZN(new_n582));
  NAND2_X1  g157(.A1(G79), .A2(G543), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n511), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(G54), .B2(new_n525), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n580), .A2(new_n581), .A3(new_n585), .ZN(new_n586));
  MUX2_X1   g161(.A(new_n586), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g162(.A(new_n586), .B(G301), .S(G868), .Z(G321));
  MUX2_X1   g163(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g164(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g165(.A(new_n586), .ZN(new_n591));
  INV_X1    g166(.A(G559), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(G860), .ZN(G148));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G868), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(G868), .B2(new_n537), .ZN(G323));
  XNOR2_X1  g171(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g172(.A1(new_n469), .A2(G2105), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n495), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT12), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT13), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(G2100), .ZN(new_n602));
  OR2_X1    g177(.A1(G99), .A2(G2105), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n603), .B(G2104), .C1(G111), .C2(new_n478), .ZN(new_n604));
  INV_X1    g179(.A(G123), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n484), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(new_n490), .B2(G135), .ZN(new_n607));
  INV_X1    g182(.A(G2096), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n602), .A2(new_n609), .A3(new_n610), .ZN(G156));
  INV_X1    g186(.A(G14), .ZN(new_n612));
  XNOR2_X1  g187(.A(G2427), .B(G2438), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2430), .ZN(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT15), .B(G2435), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n616), .A2(KEYINPUT14), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(G2443), .B(G2446), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(G2451), .B(G2454), .Z(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n620), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(G1341), .B(G1348), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n612), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  AND2_X1   g202(.A1(new_n627), .A2(KEYINPUT78), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n627), .A2(KEYINPUT78), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(G401));
  NOR2_X1   g206(.A1(G2072), .A2(G2078), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n444), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT17), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2067), .B(G2678), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT79), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n633), .A2(KEYINPUT80), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n633), .A2(KEYINPUT80), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2084), .B(G2090), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n638), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT81), .ZN(new_n644));
  INV_X1    g219(.A(new_n633), .ZN(new_n645));
  NOR3_X1   g220(.A1(new_n636), .A2(new_n645), .A3(new_n642), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT18), .ZN(new_n647));
  OR3_X1    g222(.A1(new_n634), .A2(new_n637), .A3(new_n642), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n644), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2096), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT82), .B(G2100), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n652), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(G227));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT84), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT83), .B(KEYINPUT19), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1956), .B(G2474), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n659), .B2(new_n663), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n659), .A2(new_n664), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1991), .B(G1996), .Z(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n676), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  AND3_X1   g254(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n679), .B1(new_n677), .B2(new_n678), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(G229));
  MUX2_X1   g257(.A(G6), .B(G305), .S(G16), .Z(new_n683));
  XOR2_X1   g258(.A(KEYINPUT32), .B(G1981), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G22), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G166), .B2(new_n686), .ZN(new_n688));
  INV_X1    g263(.A(G1971), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n686), .A2(G23), .ZN(new_n691));
  INV_X1    g266(.A(G288), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(new_n686), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT33), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n685), .A2(new_n690), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT34), .Z(new_n697));
  NOR2_X1   g272(.A1(G25), .A2(G29), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n490), .A2(G131), .ZN(new_n699));
  INV_X1    g274(.A(G119), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n478), .A2(G107), .ZN(new_n701));
  OAI21_X1  g276(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n702));
  OAI22_X1  g277(.A1(new_n484), .A2(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n698), .B1(new_n704), .B2(G29), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT86), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT35), .B(G1991), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n708), .A2(KEYINPUT87), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(KEYINPUT87), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT88), .ZN(new_n711));
  OR2_X1    g286(.A1(G16), .A2(G24), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G290), .B2(new_n686), .ZN(new_n713));
  INV_X1    g288(.A(G1986), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n711), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n714), .B2(new_n713), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n697), .A2(new_n709), .A3(new_n710), .A4(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT36), .Z(new_n718));
  NAND3_X1  g293(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT25), .Z(new_n720));
  INV_X1    g295(.A(G139), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n495), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n722));
  OAI221_X1 g297(.A(new_n720), .B1(new_n489), .B2(new_n721), .C1(new_n478), .C2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT92), .Z(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n725), .B2(G33), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(new_n442), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT93), .Z(new_n729));
  NAND2_X1  g304(.A1(G164), .A2(G29), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G27), .B2(G29), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n731), .A2(new_n443), .ZN(new_n732));
  NAND3_X1  g307(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT26), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n735), .A2(new_n736), .B1(G105), .B2(new_n598), .ZN(new_n737));
  INV_X1    g312(.A(G129), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n484), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n490), .B2(G141), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(new_n725), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n725), .B2(G32), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT27), .B(G1996), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT94), .ZN(new_n744));
  OAI22_X1  g319(.A1(new_n742), .A2(new_n744), .B1(new_n443), .B2(new_n731), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n686), .A2(G5), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G171), .B2(new_n686), .ZN(new_n747));
  AOI211_X1 g322(.A(new_n732), .B(new_n745), .C1(G1961), .C2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(G160), .A2(G29), .ZN(new_n749));
  INV_X1    g324(.A(G34), .ZN(new_n750));
  AOI21_X1  g325(.A(G29), .B1(new_n750), .B2(KEYINPUT24), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(KEYINPUT24), .B2(new_n750), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(G2084), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(G2084), .ZN(new_n755));
  INV_X1    g330(.A(G11), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(KEYINPUT31), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(KEYINPUT31), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT30), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n759), .A2(G28), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n725), .B1(new_n759), .B2(G28), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n757), .B(new_n758), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n607), .B2(G29), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n754), .A2(new_n755), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n727), .B2(new_n442), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n748), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n725), .A2(G35), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G162), .B2(new_n725), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT29), .Z(new_n769));
  INV_X1    g344(.A(G2090), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n686), .A2(G21), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G168), .B2(new_n686), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT95), .B(G1966), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n742), .A2(new_n744), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n775), .B(new_n776), .C1(G1961), .C2(new_n747), .ZN(new_n777));
  NOR4_X1   g352(.A1(new_n729), .A2(new_n766), .A3(new_n771), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n686), .A2(G20), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT23), .Z(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G299), .B2(G16), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G1956), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n770), .B2(new_n769), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT96), .Z(new_n784));
  NOR2_X1   g359(.A1(G4), .A2(G16), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n591), .B2(G16), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT89), .B(G1348), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n725), .A2(G26), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT28), .ZN(new_n790));
  OAI21_X1  g365(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n791));
  INV_X1    g366(.A(G116), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(G2105), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT90), .ZN(new_n794));
  INV_X1    g369(.A(G128), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n484), .ZN(new_n796));
  INV_X1    g371(.A(G140), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n489), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n790), .B1(new_n799), .B2(new_n725), .ZN(new_n800));
  INV_X1    g375(.A(G2067), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n686), .A2(G19), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n537), .B2(new_n686), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(G1341), .Z(new_n805));
  NAND3_X1  g380(.A1(new_n788), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT91), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n778), .A2(new_n784), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(KEYINPUT97), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT97), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n778), .A2(new_n810), .A3(new_n784), .A4(new_n807), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n718), .B1(new_n809), .B2(new_n811), .ZN(G311));
  INV_X1    g387(.A(G311), .ZN(G150));
  INV_X1    g388(.A(G93), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT98), .B(G55), .Z(new_n815));
  OAI22_X1  g390(.A1(new_n505), .A2(new_n814), .B1(new_n507), .B2(new_n815), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(new_n511), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(G860), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT37), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n586), .A2(new_n592), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT38), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n537), .A2(new_n819), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n537), .A2(new_n819), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n824), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT99), .Z(new_n830));
  OAI21_X1  g405(.A(new_n820), .B1(new_n828), .B2(KEYINPUT39), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n822), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT100), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(G145));
  OAI21_X1  g409(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT102), .ZN(new_n836));
  INV_X1    g411(.A(G118), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n835), .A2(new_n836), .B1(new_n837), .B2(G2105), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(new_n836), .B2(new_n835), .ZN(new_n839));
  INV_X1    g414(.A(G130), .ZN(new_n840));
  INV_X1    g415(.A(G142), .ZN(new_n841));
  OAI221_X1 g416(.A(new_n839), .B1(new_n840), .B2(new_n484), .C1(new_n489), .C2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n600), .ZN(new_n843));
  OR3_X1    g418(.A1(new_n796), .A2(G164), .A3(new_n798), .ZN(new_n844));
  OAI21_X1  g419(.A(G164), .B1(new_n796), .B2(new_n798), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n740), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n844), .A2(new_n740), .A3(new_n845), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n848), .A2(new_n723), .A3(new_n849), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n850), .A2(KEYINPUT101), .ZN(new_n851));
  INV_X1    g426(.A(new_n849), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n740), .B1(new_n844), .B2(new_n845), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n724), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT101), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n848), .A2(new_n855), .A3(new_n723), .A4(new_n849), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n704), .B1(new_n851), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n850), .A2(KEYINPUT101), .ZN(new_n859));
  INV_X1    g434(.A(new_n704), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n859), .A2(new_n860), .A3(new_n854), .A4(new_n856), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n843), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n858), .A2(new_n843), .A3(new_n861), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(G162), .B(new_n607), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(G160), .Z(new_n867));
  AOI21_X1  g442(.A(G37), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT103), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n858), .A2(new_n843), .A3(new_n861), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n870), .A2(new_n862), .ZN(new_n871));
  INV_X1    g446(.A(new_n867), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NOR4_X1   g448(.A1(new_n870), .A2(new_n862), .A3(KEYINPUT103), .A4(new_n867), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n868), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g451(.A(new_n827), .B(KEYINPUT104), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n594), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n586), .A2(G299), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n551), .A2(new_n555), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n880), .A2(new_n580), .A3(new_n581), .A4(new_n585), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT41), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT41), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n879), .A2(new_n884), .A3(new_n881), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n878), .A2(new_n886), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n887), .A2(KEYINPUT105), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(KEYINPUT105), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n878), .A2(new_n882), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(G290), .A2(G288), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n572), .A2(new_n692), .A3(new_n574), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n894), .A2(new_n895), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT106), .ZN(new_n900));
  XNOR2_X1  g475(.A(G303), .B(G305), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n900), .A2(new_n901), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n905), .B1(KEYINPUT107), .B2(KEYINPUT42), .ZN(new_n906));
  INV_X1    g481(.A(new_n892), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n888), .A2(new_n907), .A3(new_n889), .A4(new_n890), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n893), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n906), .B1(new_n893), .B2(new_n908), .ZN(new_n910));
  OAI21_X1  g485(.A(G868), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(G868), .B2(new_n819), .ZN(G295));
  OAI21_X1  g487(.A(new_n911), .B1(G868), .B2(new_n819), .ZN(G331));
  NAND2_X1  g488(.A1(G171), .A2(G168), .ZN(new_n914));
  NAND3_X1  g489(.A1(G286), .A2(new_n529), .A3(new_n530), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n827), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n914), .A2(new_n825), .A3(new_n826), .A4(new_n915), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(new_n882), .ZN(new_n920));
  AOI22_X1  g495(.A1(new_n883), .A2(new_n885), .B1(new_n917), .B2(new_n918), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(G37), .B1(new_n905), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n904), .B1(new_n920), .B2(new_n921), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n885), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n879), .A2(new_n881), .A3(KEYINPUT109), .A4(new_n884), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n883), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT110), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(new_n933), .A3(new_n919), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n932), .A2(new_n919), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT110), .B1(new_n919), .B2(new_n882), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n904), .B(new_n934), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n923), .A2(new_n937), .A3(new_n926), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n928), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n925), .A2(new_n927), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n923), .A2(new_n937), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n940), .B1(KEYINPUT43), .B2(new_n941), .ZN(new_n942));
  MUX2_X1   g517(.A(new_n939), .B(new_n942), .S(KEYINPUT44), .Z(G397));
  INV_X1    g518(.A(KEYINPUT126), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n474), .A2(new_n480), .A3(G40), .A4(new_n482), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n947));
  INV_X1    g522(.A(G1384), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n497), .B2(new_n501), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n799), .B(new_n801), .ZN(new_n952));
  INV_X1    g527(.A(G1996), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n740), .B(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n704), .B(new_n707), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(G290), .B(new_n714), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n951), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n949), .A2(KEYINPUT50), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT50), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n962), .B(new_n948), .C1(new_n497), .C2(new_n501), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n946), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT118), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1348), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n945), .B1(new_n949), .B2(KEYINPUT50), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(KEYINPUT118), .A3(new_n963), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT119), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n949), .A2(new_n945), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n801), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n971), .B1(new_n970), .B2(new_n973), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G1956), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n961), .A2(new_n946), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT115), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n963), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n968), .A2(KEYINPUT115), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n977), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(G299), .A2(KEYINPUT57), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT57), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(new_n551), .B2(new_n555), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n949), .A2(new_n947), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n945), .B1(new_n949), .B2(new_n947), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT56), .B(G2072), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n982), .A2(new_n986), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n976), .A2(new_n591), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n963), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n993), .B1(new_n968), .B2(KEYINPUT115), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n978), .A2(new_n979), .ZN(new_n995));
  AOI21_X1  g570(.A(G1956), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n990), .ZN(new_n997));
  OAI22_X1  g572(.A1(new_n996), .A2(new_n997), .B1(new_n985), .B2(new_n983), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n992), .A2(new_n998), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n974), .A2(new_n975), .A3(KEYINPUT60), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT60), .B1(new_n974), .B2(new_n975), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n591), .ZN(new_n1002));
  OAI211_X1 g577(.A(KEYINPUT60), .B(new_n586), .C1(new_n974), .C2(new_n975), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1000), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n987), .A2(new_n988), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT58), .B(G1341), .ZN(new_n1006));
  OAI22_X1  g581(.A1(new_n1005), .A2(G1996), .B1(new_n972), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n537), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1008), .B(KEYINPUT59), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n998), .A2(new_n991), .A3(KEYINPUT61), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT120), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n998), .A2(new_n991), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT61), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n998), .B2(new_n1011), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1009), .B(new_n1010), .C1(new_n1012), .C2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n999), .B1(new_n1004), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT121), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT121), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n999), .B(new_n1018), .C1(new_n1004), .C2(new_n1015), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT116), .B(G2084), .Z(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT117), .B1(new_n964), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1005), .A2(new_n774), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1020), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n968), .A2(new_n1023), .A3(new_n963), .A4(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1021), .A2(new_n1022), .A3(G168), .A4(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT51), .B1(new_n1026), .B2(G8), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1026), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(KEYINPUT122), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT122), .ZN(new_n1031));
  INV_X1    g606(.A(G8), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n1033), .B2(new_n1021), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1027), .A2(new_n1031), .B1(new_n1034), .B2(G286), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1030), .A2(new_n1035), .ZN(new_n1036));
  XOR2_X1   g611(.A(KEYINPUT111), .B(G2090), .Z(new_n1037));
  NAND3_X1  g612(.A1(new_n994), .A2(new_n995), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1971), .B1(new_n987), .B2(new_n988), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1032), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(G166), .A2(new_n1032), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(G166), .B2(new_n1032), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n1041), .A2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n972), .A2(new_n1032), .ZN(new_n1049));
  INV_X1    g624(.A(G1976), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT52), .B1(G288), .B2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1049), .B(new_n1051), .C1(new_n1050), .C2(G288), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1049), .ZN(new_n1053));
  NOR2_X1   g628(.A1(G288), .A2(new_n1050), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT52), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n567), .A2(new_n568), .ZN(new_n1056));
  OAI21_X1  g631(.A(G1981), .B1(new_n1056), .B2(new_n565), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n1058));
  INV_X1    g633(.A(G1981), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n566), .A2(new_n1059), .A3(new_n567), .A4(new_n568), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1057), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(G305), .A2(KEYINPUT114), .A3(G1981), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1063), .A2(KEYINPUT49), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1049), .B1(new_n1063), .B2(KEYINPUT49), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1052), .B(new_n1055), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1037), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1040), .B(KEYINPUT112), .C1(new_n964), .C2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT112), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n964), .A2(new_n1068), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1070), .B1(new_n1071), .B2(new_n1039), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1069), .A2(new_n1072), .A3(new_n1047), .A4(G8), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1048), .A2(new_n1067), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n987), .A2(new_n988), .A3(new_n443), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1076), .B(KEYINPUT53), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n966), .A2(new_n969), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1077), .B1(new_n1078), .B2(G1961), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(G171), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1077), .B(G301), .C1(G1961), .C2(new_n1078), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1081), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1036), .B(new_n1075), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1017), .A2(new_n1019), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1036), .A2(KEYINPUT62), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1030), .A2(new_n1035), .A3(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1074), .A2(new_n1080), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1060), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1094));
  NOR2_X1   g669(.A1(G288), .A2(G1976), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI22_X1  g671(.A1(new_n1096), .A2(new_n1053), .B1(new_n1073), .B2(new_n1066), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT63), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1034), .A2(G168), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1098), .B1(new_n1074), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1098), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1069), .A2(G8), .A3(new_n1072), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1102), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1101), .A2(new_n1073), .A3(new_n1067), .A4(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1097), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1092), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n960), .B1(new_n1087), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n950), .A2(new_n953), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(KEYINPUT46), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n950), .B1(new_n952), .B2(new_n847), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT123), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n1112), .A2(KEYINPUT47), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(KEYINPUT47), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n860), .A2(new_n707), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n955), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n799), .A2(new_n801), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n951), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT48), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n950), .A2(new_n714), .A3(new_n572), .A4(new_n574), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1120), .B(KEYINPUT124), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1119), .A2(new_n1121), .B1(new_n957), .B2(new_n950), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1121), .A2(new_n1119), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1118), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1113), .A2(new_n1114), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1125), .B(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n944), .B1(new_n1107), .B2(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1125), .B(KEYINPUT125), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1092), .A2(new_n1105), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1085), .B1(new_n1016), .B2(KEYINPUT121), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1130), .B1(new_n1131), .B2(new_n1019), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1129), .B(KEYINPUT126), .C1(new_n1132), .C2(new_n960), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1128), .A2(new_n1133), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g709(.A(new_n464), .B1(new_n653), .B2(new_n654), .ZN(new_n1136));
  OAI211_X1 g710(.A(new_n1136), .B(new_n630), .C1(new_n680), .C2(new_n681), .ZN(new_n1137));
  AOI21_X1  g711(.A(new_n1137), .B1(new_n928), .B2(new_n938), .ZN(new_n1138));
  AND3_X1   g712(.A1(new_n875), .A2(new_n1138), .A3(KEYINPUT127), .ZN(new_n1139));
  AOI21_X1  g713(.A(KEYINPUT127), .B1(new_n875), .B2(new_n1138), .ZN(new_n1140));
  NOR2_X1   g714(.A1(new_n1139), .A2(new_n1140), .ZN(G308));
  NAND2_X1  g715(.A1(new_n875), .A2(new_n1138), .ZN(G225));
endmodule


