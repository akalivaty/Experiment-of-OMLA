

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599;

  AND2_X2 U323 ( .A1(n474), .A2(n473), .ZN(n292) );
  XNOR2_X1 U324 ( .A(n303), .B(n302), .ZN(n325) );
  NOR2_X1 U325 ( .A1(n374), .A2(n373), .ZN(n492) );
  AND2_X1 U326 ( .A1(n580), .A2(n579), .ZN(n585) );
  XNOR2_X1 U327 ( .A(n308), .B(n291), .ZN(n309) );
  XOR2_X1 U328 ( .A(KEYINPUT106), .B(n458), .Z(n531) );
  XOR2_X1 U329 ( .A(n359), .B(n358), .Z(n580) );
  XOR2_X1 U330 ( .A(G148GAT), .B(G85GAT), .Z(n291) );
  INV_X1 U331 ( .A(n594), .ZN(n473) );
  INV_X1 U332 ( .A(KEYINPUT3), .ZN(n300) );
  XNOR2_X1 U333 ( .A(G155GAT), .B(KEYINPUT86), .ZN(n299) );
  XNOR2_X1 U334 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U335 ( .A(G99GAT), .B(G85GAT), .Z(n452) );
  NOR2_X1 U336 ( .A1(n550), .A2(n522), .ZN(n533) );
  XNOR2_X1 U337 ( .A(n425), .B(n330), .ZN(n331) );
  XNOR2_X1 U338 ( .A(n332), .B(n331), .ZN(n334) );
  XNOR2_X1 U339 ( .A(n310), .B(n309), .ZN(n368) );
  XOR2_X1 U340 ( .A(n415), .B(n414), .Z(n586) );
  INV_X1 U341 ( .A(G106GAT), .ZN(n459) );
  XOR2_X1 U342 ( .A(KEYINPUT38), .B(n506), .Z(n513) );
  XNOR2_X1 U343 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U344 ( .A(n462), .B(n461), .ZN(G1339GAT) );
  XOR2_X1 U345 ( .A(G29GAT), .B(G134GAT), .Z(n396) );
  XOR2_X1 U346 ( .A(n396), .B(KEYINPUT89), .Z(n294) );
  NAND2_X1 U347 ( .A1(G225GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U348 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U349 ( .A(KEYINPUT5), .B(KEYINPUT91), .Z(n296) );
  XNOR2_X1 U350 ( .A(KEYINPUT90), .B(KEYINPUT1), .ZN(n295) );
  XNOR2_X1 U351 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U352 ( .A(n298), .B(n297), .Z(n305) );
  XOR2_X1 U353 ( .A(G113GAT), .B(KEYINPUT0), .Z(n353) );
  XNOR2_X1 U354 ( .A(n299), .B(KEYINPUT2), .ZN(n303) );
  XNOR2_X1 U355 ( .A(G141GAT), .B(G162GAT), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n353), .B(n325), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n310) );
  XOR2_X1 U358 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n307) );
  XOR2_X1 U359 ( .A(G1GAT), .B(G127GAT), .Z(n379) );
  XOR2_X1 U360 ( .A(G120GAT), .B(G57GAT), .Z(n441) );
  XNOR2_X1 U361 ( .A(n379), .B(n441), .ZN(n306) );
  XNOR2_X1 U362 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U363 ( .A(KEYINPUT87), .B(KEYINPUT24), .Z(n312) );
  XNOR2_X1 U364 ( .A(KEYINPUT88), .B(KEYINPUT22), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U366 ( .A(n313), .B(KEYINPUT23), .Z(n315) );
  XOR2_X1 U367 ( .A(G50GAT), .B(KEYINPUT75), .Z(n404) );
  XNOR2_X1 U368 ( .A(G22GAT), .B(n404), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n315), .B(n314), .ZN(n321) );
  XOR2_X1 U370 ( .A(G78GAT), .B(G148GAT), .Z(n317) );
  XNOR2_X1 U371 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n446) );
  XOR2_X1 U373 ( .A(G204GAT), .B(n446), .Z(n319) );
  NAND2_X1 U374 ( .A1(G228GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U375 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U376 ( .A(n321), .B(n320), .Z(n327) );
  XOR2_X1 U377 ( .A(KEYINPUT21), .B(G218GAT), .Z(n323) );
  XNOR2_X1 U378 ( .A(KEYINPUT85), .B(G211GAT), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U380 ( .A(G197GAT), .B(n324), .Z(n329) );
  XNOR2_X1 U381 ( .A(n325), .B(n329), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n571) );
  XNOR2_X1 U383 ( .A(G36GAT), .B(G190GAT), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n328), .B(KEYINPUT78), .ZN(n395) );
  XNOR2_X1 U385 ( .A(n329), .B(n395), .ZN(n332) );
  XOR2_X1 U386 ( .A(G169GAT), .B(G8GAT), .Z(n425) );
  XOR2_X1 U387 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n330) );
  AND2_X1 U388 ( .A1(G226GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n340) );
  XOR2_X1 U390 ( .A(G183GAT), .B(KEYINPUT17), .Z(n336) );
  XNOR2_X1 U391 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n341) );
  XOR2_X1 U393 ( .A(G64GAT), .B(G92GAT), .Z(n338) );
  XNOR2_X1 U394 ( .A(G176GAT), .B(G204GAT), .ZN(n337) );
  XNOR2_X1 U395 ( .A(n338), .B(n337), .ZN(n440) );
  XOR2_X1 U396 ( .A(n341), .B(n440), .Z(n339) );
  XNOR2_X1 U397 ( .A(n340), .B(n339), .ZN(n528) );
  XOR2_X1 U398 ( .A(n341), .B(G15GAT), .Z(n343) );
  NAND2_X1 U399 ( .A1(G227GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n343), .B(n342), .ZN(n359) );
  XOR2_X1 U401 ( .A(G120GAT), .B(G127GAT), .Z(n345) );
  XNOR2_X1 U402 ( .A(KEYINPUT66), .B(G71GAT), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U404 ( .A(G176GAT), .B(KEYINPUT20), .Z(n347) );
  XNOR2_X1 U405 ( .A(G169GAT), .B(KEYINPUT82), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n357) );
  XOR2_X1 U408 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n351) );
  XNOR2_X1 U409 ( .A(G99GAT), .B(G190GAT), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U411 ( .A(n352), .B(G134GAT), .Z(n355) );
  XNOR2_X1 U412 ( .A(G43GAT), .B(n353), .ZN(n354) );
  XNOR2_X1 U413 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U414 ( .A(n357), .B(n356), .ZN(n358) );
  AND2_X1 U415 ( .A1(n528), .A2(n580), .ZN(n360) );
  NOR2_X1 U416 ( .A1(n571), .A2(n360), .ZN(n361) );
  XOR2_X1 U417 ( .A(KEYINPUT25), .B(n361), .Z(n365) );
  INV_X1 U418 ( .A(n580), .ZN(n535) );
  NAND2_X1 U419 ( .A1(n535), .A2(n571), .ZN(n362) );
  XNOR2_X1 U420 ( .A(n362), .B(KEYINPUT26), .ZN(n551) );
  XNOR2_X1 U421 ( .A(KEYINPUT27), .B(n528), .ZN(n369) );
  INV_X1 U422 ( .A(n369), .ZN(n363) );
  NOR2_X1 U423 ( .A1(n551), .A2(n363), .ZN(n364) );
  NOR2_X1 U424 ( .A1(n365), .A2(n364), .ZN(n366) );
  XOR2_X1 U425 ( .A(KEYINPUT97), .B(n366), .Z(n367) );
  NOR2_X1 U426 ( .A1(n368), .A2(n367), .ZN(n374) );
  INV_X1 U427 ( .A(KEYINPUT96), .ZN(n372) );
  XNOR2_X1 U428 ( .A(KEYINPUT92), .B(n368), .ZN(n526) );
  NAND2_X1 U429 ( .A1(n369), .A2(n526), .ZN(n550) );
  XNOR2_X1 U430 ( .A(n571), .B(KEYINPUT28), .ZN(n522) );
  XOR2_X1 U431 ( .A(n533), .B(KEYINPUT95), .Z(n370) );
  NAND2_X1 U432 ( .A1(n370), .A2(n535), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U434 ( .A(G57GAT), .B(G78GAT), .Z(n376) );
  XNOR2_X1 U435 ( .A(G8GAT), .B(G211GAT), .ZN(n375) );
  XOR2_X1 U436 ( .A(n376), .B(n375), .Z(n391) );
  XOR2_X1 U437 ( .A(KEYINPUT80), .B(KEYINPUT14), .Z(n378) );
  XNOR2_X1 U438 ( .A(G64GAT), .B(KEYINPUT79), .ZN(n377) );
  XNOR2_X1 U439 ( .A(n378), .B(n377), .ZN(n383) );
  XOR2_X1 U440 ( .A(G71GAT), .B(KEYINPUT13), .Z(n445) );
  XOR2_X1 U441 ( .A(n379), .B(n445), .Z(n381) );
  XNOR2_X1 U442 ( .A(G183GAT), .B(G155GAT), .ZN(n380) );
  XNOR2_X1 U443 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U444 ( .A(n383), .B(n382), .Z(n385) );
  NAND2_X1 U445 ( .A1(G231GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U446 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U447 ( .A(n386), .B(KEYINPUT15), .Z(n389) );
  XNOR2_X1 U448 ( .A(G15GAT), .B(G22GAT), .ZN(n387) );
  XNOR2_X1 U449 ( .A(n387), .B(KEYINPUT71), .ZN(n433) );
  XNOR2_X1 U450 ( .A(n433), .B(KEYINPUT12), .ZN(n388) );
  XNOR2_X1 U451 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U452 ( .A(n391), .B(n390), .ZN(n564) );
  INV_X1 U453 ( .A(n564), .ZN(n598) );
  NOR2_X1 U454 ( .A1(n492), .A2(n598), .ZN(n392) );
  XNOR2_X1 U455 ( .A(n392), .B(KEYINPUT103), .ZN(n417) );
  XOR2_X1 U456 ( .A(KEYINPUT36), .B(KEYINPUT102), .Z(n416) );
  XOR2_X1 U457 ( .A(KEYINPUT10), .B(G92GAT), .Z(n394) );
  XNOR2_X1 U458 ( .A(G106GAT), .B(KEYINPUT77), .ZN(n393) );
  XNOR2_X1 U459 ( .A(n394), .B(n393), .ZN(n415) );
  XNOR2_X1 U460 ( .A(n396), .B(n395), .ZN(n397) );
  AND2_X1 U461 ( .A1(G232GAT), .A2(G233GAT), .ZN(n398) );
  NAND2_X1 U462 ( .A1(n397), .A2(n398), .ZN(n402) );
  INV_X1 U463 ( .A(n397), .ZN(n400) );
  INV_X1 U464 ( .A(n398), .ZN(n399) );
  NAND2_X1 U465 ( .A1(n400), .A2(n399), .ZN(n401) );
  NAND2_X1 U466 ( .A1(n402), .A2(n401), .ZN(n403) );
  XNOR2_X1 U467 ( .A(n403), .B(G162GAT), .ZN(n409) );
  XOR2_X1 U468 ( .A(KEYINPUT11), .B(n452), .Z(n406) );
  XNOR2_X1 U469 ( .A(G218GAT), .B(n404), .ZN(n405) );
  XNOR2_X1 U470 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U471 ( .A(n407), .B(KEYINPUT67), .Z(n408) );
  XNOR2_X1 U472 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U473 ( .A(n410), .B(KEYINPUT9), .ZN(n413) );
  XNOR2_X1 U474 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n411), .B(KEYINPUT7), .ZN(n434) );
  XOR2_X1 U476 ( .A(n434), .B(KEYINPUT76), .Z(n412) );
  XNOR2_X1 U477 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U478 ( .A(n416), .B(n586), .ZN(n484) );
  NOR2_X1 U479 ( .A1(n417), .A2(n484), .ZN(n419) );
  XOR2_X1 U480 ( .A(KEYINPUT104), .B(KEYINPUT37), .Z(n418) );
  XNOR2_X1 U481 ( .A(n419), .B(n418), .ZN(n505) );
  XOR2_X1 U482 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n421) );
  XNOR2_X1 U483 ( .A(KEYINPUT29), .B(G1GAT), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n429) );
  XOR2_X1 U485 ( .A(G197GAT), .B(G141GAT), .Z(n423) );
  XNOR2_X1 U486 ( .A(G36GAT), .B(G113GAT), .ZN(n422) );
  XNOR2_X1 U487 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U488 ( .A(n424), .B(G50GAT), .Z(n427) );
  XNOR2_X1 U489 ( .A(n425), .B(G29GAT), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n438) );
  XOR2_X1 U492 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n431) );
  NAND2_X1 U493 ( .A1(G229GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U495 ( .A(n432), .B(KEYINPUT72), .Z(n436) );
  XNOR2_X1 U496 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U497 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U498 ( .A(n438), .B(n437), .Z(n589) );
  INV_X1 U499 ( .A(n589), .ZN(n554) );
  INV_X1 U500 ( .A(n441), .ZN(n439) );
  NAND2_X1 U501 ( .A1(n440), .A2(n439), .ZN(n444) );
  INV_X1 U502 ( .A(n440), .ZN(n442) );
  NAND2_X1 U503 ( .A1(n442), .A2(n441), .ZN(n443) );
  NAND2_X1 U504 ( .A1(n444), .A2(n443), .ZN(n448) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n448), .B(n447), .ZN(n456) );
  XOR2_X1 U507 ( .A(KEYINPUT73), .B(KEYINPUT31), .Z(n450) );
  XNOR2_X1 U508 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n449) );
  XNOR2_X1 U509 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U510 ( .A(n452), .B(n451), .Z(n454) );
  NAND2_X1 U511 ( .A1(G230GAT), .A2(G233GAT), .ZN(n453) );
  XNOR2_X1 U512 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U513 ( .A(n456), .B(n455), .Z(n594) );
  XOR2_X1 U514 ( .A(KEYINPUT41), .B(n594), .Z(n581) );
  NAND2_X1 U515 ( .A1(n554), .A2(n581), .ZN(n515) );
  INV_X1 U516 ( .A(n515), .ZN(n457) );
  NAND2_X1 U517 ( .A1(n505), .A2(n457), .ZN(n458) );
  NAND2_X1 U518 ( .A1(n531), .A2(n522), .ZN(n462) );
  XOR2_X1 U519 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n460) );
  INV_X1 U520 ( .A(G218GAT), .ZN(n488) );
  XNOR2_X1 U521 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n478) );
  INV_X1 U522 ( .A(n581), .ZN(n559) );
  NOR2_X1 U523 ( .A1(n554), .A2(n559), .ZN(n463) );
  XNOR2_X1 U524 ( .A(n463), .B(KEYINPUT46), .ZN(n464) );
  NOR2_X1 U525 ( .A1(n598), .A2(n464), .ZN(n465) );
  INV_X1 U526 ( .A(n586), .ZN(n567) );
  NAND2_X1 U527 ( .A1(n465), .A2(n567), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n466), .B(KEYINPUT109), .ZN(n467) );
  NAND2_X1 U529 ( .A1(n467), .A2(KEYINPUT47), .ZN(n471) );
  INV_X1 U530 ( .A(n467), .ZN(n469) );
  INV_X1 U531 ( .A(KEYINPUT47), .ZN(n468) );
  NAND2_X1 U532 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U533 ( .A1(n471), .A2(n470), .ZN(n476) );
  NOR2_X1 U534 ( .A1(n484), .A2(n564), .ZN(n472) );
  XNOR2_X1 U535 ( .A(n472), .B(KEYINPUT45), .ZN(n474) );
  NAND2_X1 U536 ( .A1(n292), .A2(n554), .ZN(n475) );
  NAND2_X1 U537 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(n552) );
  NAND2_X1 U539 ( .A1(n528), .A2(n552), .ZN(n480) );
  XOR2_X1 U540 ( .A(KEYINPUT54), .B(KEYINPUT121), .Z(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(n481) );
  NOR2_X1 U542 ( .A1(n481), .A2(n526), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n482), .B(KEYINPUT65), .ZN(n570) );
  NOR2_X1 U544 ( .A1(n551), .A2(n570), .ZN(n597) );
  INV_X1 U545 ( .A(n597), .ZN(n483) );
  NOR2_X1 U546 ( .A1(n484), .A2(n483), .ZN(n486) );
  XNOR2_X1 U547 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(G1355GAT) );
  XNOR2_X1 U550 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n496) );
  XOR2_X1 U551 ( .A(KEYINPUT81), .B(KEYINPUT16), .Z(n490) );
  NAND2_X1 U552 ( .A1(n598), .A2(n567), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n490), .B(n489), .ZN(n491) );
  NOR2_X1 U554 ( .A1(n492), .A2(n491), .ZN(n493) );
  XOR2_X1 U555 ( .A(KEYINPUT98), .B(n493), .Z(n516) );
  NOR2_X1 U556 ( .A1(n554), .A2(n594), .ZN(n504) );
  INV_X1 U557 ( .A(n504), .ZN(n494) );
  NOR2_X1 U558 ( .A1(n516), .A2(n494), .ZN(n501) );
  NAND2_X1 U559 ( .A1(n501), .A2(n526), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n496), .B(n495), .ZN(G1324GAT) );
  XOR2_X1 U561 ( .A(G8GAT), .B(KEYINPUT99), .Z(n498) );
  NAND2_X1 U562 ( .A1(n501), .A2(n528), .ZN(n497) );
  XNOR2_X1 U563 ( .A(n498), .B(n497), .ZN(G1325GAT) );
  XOR2_X1 U564 ( .A(G15GAT), .B(KEYINPUT35), .Z(n500) );
  NAND2_X1 U565 ( .A1(n501), .A2(n580), .ZN(n499) );
  XNOR2_X1 U566 ( .A(n500), .B(n499), .ZN(G1326GAT) );
  NAND2_X1 U567 ( .A1(n522), .A2(n501), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n502), .B(KEYINPUT100), .ZN(n503) );
  XNOR2_X1 U569 ( .A(G22GAT), .B(n503), .ZN(G1327GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n508) );
  NAND2_X1 U571 ( .A1(n505), .A2(n504), .ZN(n506) );
  NAND2_X1 U572 ( .A1(n513), .A2(n526), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U574 ( .A(n509), .B(G29GAT), .Z(G1328GAT) );
  NAND2_X1 U575 ( .A1(n513), .A2(n528), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n510), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U577 ( .A1(n513), .A2(n580), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n511), .B(KEYINPUT40), .ZN(n512) );
  XNOR2_X1 U579 ( .A(G43GAT), .B(n512), .ZN(G1330GAT) );
  NAND2_X1 U580 ( .A1(n513), .A2(n522), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n514), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n518) );
  NOR2_X1 U583 ( .A1(n516), .A2(n515), .ZN(n523) );
  NAND2_X1 U584 ( .A1(n523), .A2(n526), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U586 ( .A(G57GAT), .B(n519), .ZN(G1332GAT) );
  NAND2_X1 U587 ( .A1(n528), .A2(n523), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n520), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U589 ( .A1(n523), .A2(n580), .ZN(n521) );
  XNOR2_X1 U590 ( .A(n521), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U591 ( .A(G78GAT), .B(KEYINPUT43), .Z(n525) );
  NAND2_X1 U592 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U593 ( .A(n525), .B(n524), .ZN(G1335GAT) );
  NAND2_X1 U594 ( .A1(n526), .A2(n531), .ZN(n527) );
  XNOR2_X1 U595 ( .A(G85GAT), .B(n527), .ZN(G1336GAT) );
  XOR2_X1 U596 ( .A(G92GAT), .B(KEYINPUT107), .Z(n530) );
  NAND2_X1 U597 ( .A1(n531), .A2(n528), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n530), .B(n529), .ZN(G1337GAT) );
  NAND2_X1 U599 ( .A1(n531), .A2(n580), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n532), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U601 ( .A1(n533), .A2(n552), .ZN(n534) );
  NOR2_X1 U602 ( .A1(n535), .A2(n534), .ZN(n545) );
  NAND2_X1 U603 ( .A1(n589), .A2(n545), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n536), .B(KEYINPUT110), .ZN(n537) );
  XNOR2_X1 U605 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT49), .B(KEYINPUT112), .Z(n539) );
  NAND2_X1 U607 ( .A1(n545), .A2(n581), .ZN(n538) );
  XNOR2_X1 U608 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U609 ( .A(G120GAT), .B(KEYINPUT111), .Z(n540) );
  XNOR2_X1 U610 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n543) );
  NAND2_X1 U612 ( .A1(n545), .A2(n598), .ZN(n542) );
  XNOR2_X1 U613 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U614 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U616 ( .A1(n545), .A2(n586), .ZN(n546) );
  XNOR2_X1 U617 ( .A(n547), .B(n546), .ZN(n549) );
  XOR2_X1 U618 ( .A(G134GAT), .B(KEYINPUT115), .Z(n548) );
  XNOR2_X1 U619 ( .A(n549), .B(n548), .ZN(G1343GAT) );
  NOR2_X1 U620 ( .A1(n551), .A2(n550), .ZN(n553) );
  NAND2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n566) );
  NOR2_X1 U622 ( .A1(n554), .A2(n566), .ZN(n555) );
  XOR2_X1 U623 ( .A(KEYINPUT116), .B(n555), .Z(n556) );
  XNOR2_X1 U624 ( .A(G141GAT), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n558) );
  XNOR2_X1 U626 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n557) );
  XNOR2_X1 U627 ( .A(n558), .B(n557), .ZN(n563) );
  NOR2_X1 U628 ( .A1(n559), .A2(n566), .ZN(n561) );
  XNOR2_X1 U629 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n560) );
  XNOR2_X1 U630 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U631 ( .A(n563), .B(n562), .Z(G1345GAT) );
  NOR2_X1 U632 ( .A1(n564), .A2(n566), .ZN(n565) );
  XOR2_X1 U633 ( .A(G155GAT), .B(n565), .Z(G1346GAT) );
  NOR2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U635 ( .A(KEYINPUT120), .B(n568), .Z(n569) );
  XNOR2_X1 U636 ( .A(G162GAT), .B(n569), .ZN(G1347GAT) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U638 ( .A(n572), .B(KEYINPUT55), .Z(n579) );
  AND2_X1 U639 ( .A1(n580), .A2(n589), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n579), .A2(n573), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n574), .B(KEYINPUT122), .ZN(n575) );
  XNOR2_X1 U642 ( .A(G169GAT), .B(n575), .ZN(G1348GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n577) );
  XNOR2_X1 U644 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n576) );
  XNOR2_X1 U645 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U646 ( .A(KEYINPUT56), .B(n578), .Z(n583) );
  NAND2_X1 U647 ( .A1(n585), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1349GAT) );
  NAND2_X1 U649 ( .A1(n585), .A2(n598), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n584), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U651 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n588) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1351GAT) );
  XOR2_X1 U654 ( .A(G197GAT), .B(KEYINPUT125), .Z(n591) );
  NAND2_X1 U655 ( .A1(n597), .A2(n589), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n591), .B(n590), .ZN(n593) );
  XOR2_X1 U657 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n592) );
  XNOR2_X1 U658 ( .A(n593), .B(n592), .ZN(G1352GAT) );
  XOR2_X1 U659 ( .A(G204GAT), .B(KEYINPUT61), .Z(n596) );
  NAND2_X1 U660 ( .A1(n597), .A2(n594), .ZN(n595) );
  XNOR2_X1 U661 ( .A(n596), .B(n595), .ZN(G1353GAT) );
  NAND2_X1 U662 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U663 ( .A(n599), .B(G211GAT), .ZN(G1354GAT) );
endmodule

