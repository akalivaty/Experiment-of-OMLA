

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(G2104), .A2(G2105), .ZN(n542) );
  AND2_X1 U551 ( .A1(n549), .A2(G2104), .ZN(n886) );
  BUF_X1 U552 ( .A(n885), .Z(n517) );
  XNOR2_X1 U553 ( .A(n542), .B(n541), .ZN(n885) );
  AND2_X1 U554 ( .A1(n786), .A2(n691), .ZN(n716) );
  AND2_X1 U555 ( .A1(n716), .A2(G1996), .ZN(n702) );
  INV_X1 U556 ( .A(KEYINPUT31), .ZN(n699) );
  XOR2_X1 U557 ( .A(n745), .B(KEYINPUT94), .Z(n518) );
  INV_X1 U558 ( .A(n974), .ZN(n703) );
  AND2_X1 U559 ( .A1(n704), .A2(n703), .ZN(n705) );
  AND2_X1 U560 ( .A1(n706), .A2(n705), .ZN(n710) );
  INV_X1 U561 ( .A(KEYINPUT29), .ZN(n727) );
  XNOR2_X1 U562 ( .A(n728), .B(n727), .ZN(n731) );
  INV_X1 U563 ( .A(KEYINPUT95), .ZN(n734) );
  INV_X1 U564 ( .A(n787), .ZN(n691) );
  NOR2_X1 U565 ( .A1(n758), .A2(n757), .ZN(n759) );
  INV_X1 U566 ( .A(n716), .ZN(n736) );
  NOR2_X1 U567 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U568 ( .A1(G8), .A2(n736), .ZN(n778) );
  AND2_X1 U569 ( .A1(n885), .A2(G138), .ZN(n563) );
  NOR2_X2 U570 ( .A1(G651), .A2(n627), .ZN(n647) );
  INV_X1 U571 ( .A(KEYINPUT17), .ZN(n541) );
  XOR2_X1 U572 ( .A(KEYINPUT73), .B(n590), .Z(n970) );
  AND2_X1 U573 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U574 ( .A1(n830), .A2(n829), .ZN(n831) );
  INV_X1 U575 ( .A(G651), .ZN(n523) );
  NOR2_X1 U576 ( .A1(G543), .A2(n523), .ZN(n520) );
  XNOR2_X1 U577 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n519) );
  XNOR2_X1 U578 ( .A(n520), .B(n519), .ZN(n648) );
  NAND2_X1 U579 ( .A1(G64), .A2(n648), .ZN(n522) );
  XOR2_X1 U580 ( .A(KEYINPUT0), .B(G543), .Z(n627) );
  NAND2_X1 U581 ( .A1(G52), .A2(n647), .ZN(n521) );
  NAND2_X1 U582 ( .A1(n522), .A2(n521), .ZN(n528) );
  NOR2_X1 U583 ( .A1(G651), .A2(G543), .ZN(n651) );
  NAND2_X1 U584 ( .A1(G90), .A2(n651), .ZN(n525) );
  NOR2_X1 U585 ( .A1(n627), .A2(n523), .ZN(n655) );
  NAND2_X1 U586 ( .A1(G77), .A2(n655), .ZN(n524) );
  NAND2_X1 U587 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U588 ( .A(KEYINPUT9), .B(n526), .Z(n527) );
  NOR2_X1 U589 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U590 ( .A(KEYINPUT68), .B(n529), .Z(G301) );
  INV_X1 U591 ( .A(G301), .ZN(G171) );
  XOR2_X1 U592 ( .A(G2438), .B(G2454), .Z(n531) );
  XNOR2_X1 U593 ( .A(G2435), .B(G2430), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U595 ( .A(n532), .B(G2427), .Z(n534) );
  XNOR2_X1 U596 ( .A(G1341), .B(G1348), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n534), .B(n533), .ZN(n538) );
  XOR2_X1 U598 ( .A(G2443), .B(G2446), .Z(n536) );
  XNOR2_X1 U599 ( .A(KEYINPUT102), .B(G2451), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U601 ( .A(n538), .B(n537), .Z(n539) );
  AND2_X1 U602 ( .A1(G14), .A2(n539), .ZN(G401) );
  AND2_X1 U603 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U604 ( .A(G2105), .ZN(n549) );
  NOR2_X1 U605 ( .A1(G2104), .A2(n549), .ZN(n881) );
  NAND2_X1 U606 ( .A1(n881), .A2(G123), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n540), .B(KEYINPUT18), .ZN(n544) );
  NAND2_X1 U608 ( .A1(G135), .A2(n517), .ZN(n543) );
  NAND2_X1 U609 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U610 ( .A(KEYINPUT78), .B(n545), .ZN(n548) );
  AND2_X1 U611 ( .A1(G2104), .A2(G2105), .ZN(n882) );
  NAND2_X1 U612 ( .A1(G111), .A2(n882), .ZN(n546) );
  XNOR2_X1 U613 ( .A(KEYINPUT79), .B(n546), .ZN(n547) );
  NOR2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n551) );
  NAND2_X1 U615 ( .A1(n886), .A2(G99), .ZN(n550) );
  NAND2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n923) );
  XNOR2_X1 U617 ( .A(G2096), .B(n923), .ZN(n552) );
  OR2_X1 U618 ( .A1(G2100), .A2(n552), .ZN(G156) );
  NAND2_X1 U619 ( .A1(G65), .A2(n648), .ZN(n554) );
  NAND2_X1 U620 ( .A1(G53), .A2(n647), .ZN(n553) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U622 ( .A1(G91), .A2(n651), .ZN(n556) );
  NAND2_X1 U623 ( .A1(G78), .A2(n655), .ZN(n555) );
  NAND2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n967) );
  INV_X1 U626 ( .A(n967), .ZN(G299) );
  NAND2_X1 U627 ( .A1(G126), .A2(n881), .ZN(n560) );
  NAND2_X1 U628 ( .A1(G114), .A2(n882), .ZN(n559) );
  NAND2_X1 U629 ( .A1(n560), .A2(n559), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n886), .A2(G102), .ZN(n561) );
  XOR2_X1 U631 ( .A(KEYINPUT85), .B(n561), .Z(n565) );
  INV_X1 U632 ( .A(KEYINPUT86), .ZN(n562) );
  XNOR2_X1 U633 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U634 ( .A(n566), .B(KEYINPUT87), .ZN(n567) );
  NOR2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n690) );
  BUF_X1 U636 ( .A(n690), .Z(G164) );
  INV_X1 U637 ( .A(G132), .ZN(G219) );
  INV_X1 U638 ( .A(G82), .ZN(G220) );
  NAND2_X1 U639 ( .A1(G7), .A2(G661), .ZN(n569) );
  XNOR2_X1 U640 ( .A(n569), .B(KEYINPUT10), .ZN(n570) );
  XOR2_X1 U641 ( .A(KEYINPUT70), .B(n570), .Z(n915) );
  NAND2_X1 U642 ( .A1(n915), .A2(G567), .ZN(n571) );
  XOR2_X1 U643 ( .A(KEYINPUT11), .B(n571), .Z(G234) );
  INV_X1 U644 ( .A(G860), .ZN(n616) );
  NAND2_X1 U645 ( .A1(G56), .A2(n648), .ZN(n572) );
  XOR2_X1 U646 ( .A(KEYINPUT14), .B(n572), .Z(n578) );
  NAND2_X1 U647 ( .A1(n651), .A2(G81), .ZN(n573) );
  XNOR2_X1 U648 ( .A(n573), .B(KEYINPUT12), .ZN(n575) );
  NAND2_X1 U649 ( .A1(G68), .A2(n655), .ZN(n574) );
  NAND2_X1 U650 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U651 ( .A(KEYINPUT13), .B(n576), .Z(n577) );
  NOR2_X1 U652 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U653 ( .A1(n647), .A2(G43), .ZN(n579) );
  NAND2_X1 U654 ( .A1(n580), .A2(n579), .ZN(n974) );
  NOR2_X1 U655 ( .A1(n616), .A2(n974), .ZN(n581) );
  XNOR2_X1 U656 ( .A(n581), .B(KEYINPUT71), .ZN(G153) );
  NAND2_X1 U657 ( .A1(G301), .A2(G868), .ZN(n592) );
  NAND2_X1 U658 ( .A1(G79), .A2(n655), .ZN(n588) );
  NAND2_X1 U659 ( .A1(G92), .A2(n651), .ZN(n583) );
  NAND2_X1 U660 ( .A1(G66), .A2(n648), .ZN(n582) );
  NAND2_X1 U661 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U662 ( .A1(n647), .A2(G54), .ZN(n584) );
  XOR2_X1 U663 ( .A(KEYINPUT72), .B(n584), .Z(n585) );
  NAND2_X1 U664 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U665 ( .A(n589), .B(KEYINPUT15), .ZN(n590) );
  INV_X1 U666 ( .A(n970), .ZN(n712) );
  INV_X1 U667 ( .A(G868), .ZN(n609) );
  NAND2_X1 U668 ( .A1(n712), .A2(n609), .ZN(n591) );
  NAND2_X1 U669 ( .A1(n592), .A2(n591), .ZN(G284) );
  NAND2_X1 U670 ( .A1(n651), .A2(G89), .ZN(n593) );
  XNOR2_X1 U671 ( .A(n593), .B(KEYINPUT4), .ZN(n595) );
  NAND2_X1 U672 ( .A1(G76), .A2(n655), .ZN(n594) );
  NAND2_X1 U673 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U674 ( .A(n596), .B(KEYINPUT5), .ZN(n601) );
  NAND2_X1 U675 ( .A1(G63), .A2(n648), .ZN(n598) );
  NAND2_X1 U676 ( .A1(G51), .A2(n647), .ZN(n597) );
  NAND2_X1 U677 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U678 ( .A(KEYINPUT6), .B(n599), .Z(n600) );
  NAND2_X1 U679 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U680 ( .A(n602), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U681 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U682 ( .A1(G286), .A2(n609), .ZN(n603) );
  XNOR2_X1 U683 ( .A(n603), .B(KEYINPUT74), .ZN(n605) );
  NOR2_X1 U684 ( .A1(G299), .A2(G868), .ZN(n604) );
  NOR2_X1 U685 ( .A1(n605), .A2(n604), .ZN(G297) );
  NAND2_X1 U686 ( .A1(n616), .A2(G559), .ZN(n606) );
  NAND2_X1 U687 ( .A1(n606), .A2(n970), .ZN(n607) );
  XNOR2_X1 U688 ( .A(n607), .B(KEYINPUT16), .ZN(n608) );
  XOR2_X1 U689 ( .A(KEYINPUT75), .B(n608), .Z(G148) );
  NOR2_X1 U690 ( .A1(n712), .A2(n609), .ZN(n610) );
  XOR2_X1 U691 ( .A(KEYINPUT76), .B(n610), .Z(n611) );
  NOR2_X1 U692 ( .A1(G559), .A2(n611), .ZN(n612) );
  XOR2_X1 U693 ( .A(KEYINPUT77), .B(n612), .Z(n614) );
  NOR2_X1 U694 ( .A1(G868), .A2(n974), .ZN(n613) );
  NOR2_X1 U695 ( .A1(n614), .A2(n613), .ZN(G282) );
  NAND2_X1 U696 ( .A1(G559), .A2(n970), .ZN(n615) );
  XOR2_X1 U697 ( .A(n974), .B(n615), .Z(n663) );
  NAND2_X1 U698 ( .A1(n616), .A2(n663), .ZN(n623) );
  NAND2_X1 U699 ( .A1(G67), .A2(n648), .ZN(n618) );
  NAND2_X1 U700 ( .A1(G55), .A2(n647), .ZN(n617) );
  NAND2_X1 U701 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U702 ( .A1(G93), .A2(n651), .ZN(n620) );
  NAND2_X1 U703 ( .A1(G80), .A2(n655), .ZN(n619) );
  NAND2_X1 U704 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U705 ( .A1(n622), .A2(n621), .ZN(n665) );
  XOR2_X1 U706 ( .A(n623), .B(n665), .Z(G145) );
  NAND2_X1 U707 ( .A1(G49), .A2(n647), .ZN(n625) );
  NAND2_X1 U708 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U709 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U710 ( .A1(n648), .A2(n626), .ZN(n629) );
  NAND2_X1 U711 ( .A1(n627), .A2(G87), .ZN(n628) );
  NAND2_X1 U712 ( .A1(n629), .A2(n628), .ZN(G288) );
  XOR2_X1 U713 ( .A(KEYINPUT2), .B(KEYINPUT81), .Z(n631) );
  NAND2_X1 U714 ( .A1(G73), .A2(n655), .ZN(n630) );
  XNOR2_X1 U715 ( .A(n631), .B(n630), .ZN(n638) );
  NAND2_X1 U716 ( .A1(G61), .A2(n648), .ZN(n633) );
  NAND2_X1 U717 ( .A1(G48), .A2(n647), .ZN(n632) );
  NAND2_X1 U718 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U719 ( .A1(n651), .A2(G86), .ZN(n634) );
  XOR2_X1 U720 ( .A(KEYINPUT80), .B(n634), .Z(n635) );
  NOR2_X1 U721 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U722 ( .A1(n638), .A2(n637), .ZN(G305) );
  NAND2_X1 U723 ( .A1(G62), .A2(n648), .ZN(n640) );
  NAND2_X1 U724 ( .A1(G50), .A2(n647), .ZN(n639) );
  NAND2_X1 U725 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U726 ( .A(KEYINPUT82), .B(n641), .ZN(n645) );
  NAND2_X1 U727 ( .A1(G88), .A2(n651), .ZN(n643) );
  NAND2_X1 U728 ( .A1(G75), .A2(n655), .ZN(n642) );
  NAND2_X1 U729 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U730 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U731 ( .A(KEYINPUT83), .B(n646), .ZN(G303) );
  INV_X1 U732 ( .A(G303), .ZN(G166) );
  NAND2_X1 U733 ( .A1(n647), .A2(G47), .ZN(n650) );
  NAND2_X1 U734 ( .A1(n648), .A2(G60), .ZN(n649) );
  NAND2_X1 U735 ( .A1(n650), .A2(n649), .ZN(n654) );
  NAND2_X1 U736 ( .A1(G85), .A2(n651), .ZN(n652) );
  XOR2_X1 U737 ( .A(KEYINPUT66), .B(n652), .Z(n653) );
  NOR2_X1 U738 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U739 ( .A1(n655), .A2(G72), .ZN(n656) );
  NAND2_X1 U740 ( .A1(n657), .A2(n656), .ZN(G290) );
  XNOR2_X1 U741 ( .A(KEYINPUT19), .B(G288), .ZN(n662) );
  XNOR2_X1 U742 ( .A(n665), .B(G305), .ZN(n658) );
  XOR2_X1 U743 ( .A(n658), .B(G166), .Z(n659) );
  XOR2_X1 U744 ( .A(G299), .B(n659), .Z(n660) );
  XNOR2_X1 U745 ( .A(n660), .B(G290), .ZN(n661) );
  XNOR2_X1 U746 ( .A(n662), .B(n661), .ZN(n901) );
  XNOR2_X1 U747 ( .A(n663), .B(n901), .ZN(n664) );
  NAND2_X1 U748 ( .A1(n664), .A2(G868), .ZN(n667) );
  OR2_X1 U749 ( .A1(G868), .A2(n665), .ZN(n666) );
  NAND2_X1 U750 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U751 ( .A1(G2084), .A2(G2078), .ZN(n668) );
  XOR2_X1 U752 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U753 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U754 ( .A(KEYINPUT21), .B(n670), .ZN(n671) );
  NAND2_X1 U755 ( .A1(n671), .A2(G2072), .ZN(n672) );
  XNOR2_X1 U756 ( .A(KEYINPUT84), .B(n672), .ZN(G158) );
  XNOR2_X1 U757 ( .A(KEYINPUT69), .B(G57), .ZN(G237) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U759 ( .A1(G108), .A2(G120), .ZN(n673) );
  NOR2_X1 U760 ( .A1(G237), .A2(n673), .ZN(n674) );
  NAND2_X1 U761 ( .A1(G69), .A2(n674), .ZN(n913) );
  NAND2_X1 U762 ( .A1(n913), .A2(G567), .ZN(n679) );
  NOR2_X1 U763 ( .A1(G220), .A2(G219), .ZN(n675) );
  XOR2_X1 U764 ( .A(KEYINPUT22), .B(n675), .Z(n676) );
  NOR2_X1 U765 ( .A1(G218), .A2(n676), .ZN(n677) );
  NAND2_X1 U766 ( .A1(G96), .A2(n677), .ZN(n914) );
  NAND2_X1 U767 ( .A1(n914), .A2(G2106), .ZN(n678) );
  NAND2_X1 U768 ( .A1(n679), .A2(n678), .ZN(n857) );
  NAND2_X1 U769 ( .A1(G661), .A2(G483), .ZN(n680) );
  NOR2_X1 U770 ( .A1(n857), .A2(n680), .ZN(n835) );
  NAND2_X1 U771 ( .A1(n835), .A2(G36), .ZN(G176) );
  XOR2_X1 U772 ( .A(KEYINPUT23), .B(KEYINPUT64), .Z(n682) );
  NAND2_X1 U773 ( .A1(G101), .A2(n886), .ZN(n681) );
  XNOR2_X1 U774 ( .A(n682), .B(n681), .ZN(n685) );
  NAND2_X1 U775 ( .A1(G113), .A2(n882), .ZN(n683) );
  XOR2_X1 U776 ( .A(KEYINPUT65), .B(n683), .Z(n684) );
  NAND2_X1 U777 ( .A1(n685), .A2(n684), .ZN(n689) );
  NAND2_X1 U778 ( .A1(G137), .A2(n517), .ZN(n687) );
  NAND2_X1 U779 ( .A1(G125), .A2(n881), .ZN(n686) );
  NAND2_X1 U780 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U781 ( .A1(n689), .A2(n688), .ZN(G160) );
  NOR2_X1 U782 ( .A1(n690), .A2(G1384), .ZN(n786) );
  NAND2_X1 U783 ( .A1(G160), .A2(G40), .ZN(n787) );
  NOR2_X1 U784 ( .A1(G1966), .A2(n778), .ZN(n746) );
  NOR2_X1 U785 ( .A1(G2084), .A2(n736), .ZN(n744) );
  NOR2_X1 U786 ( .A1(n746), .A2(n744), .ZN(n692) );
  NAND2_X1 U787 ( .A1(G8), .A2(n692), .ZN(n693) );
  XNOR2_X1 U788 ( .A(KEYINPUT30), .B(n693), .ZN(n694) );
  NOR2_X1 U789 ( .A1(n694), .A2(G168), .ZN(n698) );
  OR2_X1 U790 ( .A1(n716), .A2(G1961), .ZN(n696) );
  XNOR2_X1 U791 ( .A(G2078), .B(KEYINPUT25), .ZN(n942) );
  NAND2_X1 U792 ( .A1(n716), .A2(n942), .ZN(n695) );
  NAND2_X1 U793 ( .A1(n696), .A2(n695), .ZN(n729) );
  NOR2_X1 U794 ( .A1(n729), .A2(G171), .ZN(n697) );
  NOR2_X1 U795 ( .A1(n698), .A2(n697), .ZN(n700) );
  XNOR2_X1 U796 ( .A(n700), .B(n699), .ZN(n733) );
  INV_X1 U797 ( .A(KEYINPUT26), .ZN(n701) );
  XNOR2_X1 U798 ( .A(n702), .B(n701), .ZN(n706) );
  NAND2_X1 U799 ( .A1(n736), .A2(G1341), .ZN(n704) );
  NAND2_X1 U800 ( .A1(G1348), .A2(n736), .ZN(n708) );
  NAND2_X1 U801 ( .A1(G2067), .A2(n716), .ZN(n707) );
  NAND2_X1 U802 ( .A1(n708), .A2(n707), .ZN(n711) );
  NOR2_X1 U803 ( .A1(n712), .A2(n711), .ZN(n709) );
  OR2_X1 U804 ( .A1(n710), .A2(n709), .ZN(n714) );
  NAND2_X1 U805 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U806 ( .A1(n714), .A2(n713), .ZN(n721) );
  NAND2_X1 U807 ( .A1(n716), .A2(G2072), .ZN(n715) );
  XNOR2_X1 U808 ( .A(KEYINPUT27), .B(n715), .ZN(n719) );
  XNOR2_X1 U809 ( .A(G1956), .B(KEYINPUT91), .ZN(n1004) );
  NOR2_X1 U810 ( .A1(n716), .A2(n1004), .ZN(n717) );
  XNOR2_X1 U811 ( .A(n717), .B(KEYINPUT92), .ZN(n718) );
  NOR2_X1 U812 ( .A1(n719), .A2(n718), .ZN(n722) );
  NAND2_X1 U813 ( .A1(n967), .A2(n722), .ZN(n720) );
  NAND2_X1 U814 ( .A1(n721), .A2(n720), .ZN(n726) );
  NOR2_X1 U815 ( .A1(n967), .A2(n722), .ZN(n724) );
  XNOR2_X1 U816 ( .A(KEYINPUT93), .B(KEYINPUT28), .ZN(n723) );
  XNOR2_X1 U817 ( .A(n724), .B(n723), .ZN(n725) );
  NAND2_X1 U818 ( .A1(n726), .A2(n725), .ZN(n728) );
  NAND2_X1 U819 ( .A1(n729), .A2(G171), .ZN(n730) );
  NAND2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U821 ( .A1(n733), .A2(n732), .ZN(n745) );
  NAND2_X1 U822 ( .A1(G286), .A2(n745), .ZN(n735) );
  XNOR2_X1 U823 ( .A(n735), .B(n734), .ZN(n741) );
  NOR2_X1 U824 ( .A1(G1971), .A2(n778), .ZN(n738) );
  NOR2_X1 U825 ( .A1(G2090), .A2(n736), .ZN(n737) );
  NOR2_X1 U826 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U827 ( .A1(G303), .A2(n739), .ZN(n740) );
  NAND2_X1 U828 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U829 ( .A1(n742), .A2(G8), .ZN(n743) );
  XNOR2_X1 U830 ( .A(n743), .B(KEYINPUT32), .ZN(n768) );
  NAND2_X1 U831 ( .A1(G8), .A2(n744), .ZN(n748) );
  NOR2_X1 U832 ( .A1(n746), .A2(n518), .ZN(n747) );
  NAND2_X1 U833 ( .A1(n748), .A2(n747), .ZN(n769) );
  NAND2_X1 U834 ( .A1(G288), .A2(G1976), .ZN(n749) );
  XNOR2_X1 U835 ( .A(n749), .B(KEYINPUT96), .ZN(n979) );
  INV_X1 U836 ( .A(n979), .ZN(n750) );
  OR2_X1 U837 ( .A1(n750), .A2(n778), .ZN(n754) );
  INV_X1 U838 ( .A(n754), .ZN(n751) );
  AND2_X1 U839 ( .A1(n769), .A2(n751), .ZN(n752) );
  AND2_X1 U840 ( .A1(n768), .A2(n752), .ZN(n758) );
  NOR2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n761) );
  NOR2_X1 U842 ( .A1(G1971), .A2(G303), .ZN(n753) );
  NOR2_X1 U843 ( .A1(n761), .A2(n753), .ZN(n978) );
  OR2_X1 U844 ( .A1(n754), .A2(n978), .ZN(n756) );
  INV_X1 U845 ( .A(KEYINPUT33), .ZN(n755) );
  NAND2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U847 ( .A(n759), .B(KEYINPUT97), .ZN(n765) );
  XNOR2_X1 U848 ( .A(G1981), .B(KEYINPUT98), .ZN(n760) );
  XNOR2_X1 U849 ( .A(n760), .B(G305), .ZN(n965) );
  NAND2_X1 U850 ( .A1(n761), .A2(KEYINPUT33), .ZN(n762) );
  NOR2_X1 U851 ( .A1(n778), .A2(n762), .ZN(n763) );
  NOR2_X1 U852 ( .A1(n965), .A2(n763), .ZN(n764) );
  NAND2_X1 U853 ( .A1(n765), .A2(n764), .ZN(n774) );
  NOR2_X1 U854 ( .A1(G2090), .A2(G303), .ZN(n766) );
  XOR2_X1 U855 ( .A(KEYINPUT99), .B(n766), .Z(n767) );
  NAND2_X1 U856 ( .A1(G8), .A2(n767), .ZN(n771) );
  NAND2_X1 U857 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U859 ( .A1(n772), .A2(n778), .ZN(n773) );
  NAND2_X1 U860 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U861 ( .A(n775), .B(KEYINPUT100), .ZN(n821) );
  NOR2_X1 U862 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U863 ( .A(n776), .B(KEYINPUT24), .Z(n777) );
  NOR2_X1 U864 ( .A1(n778), .A2(n777), .ZN(n819) );
  XOR2_X1 U865 ( .A(KEYINPUT39), .B(KEYINPUT101), .Z(n805) );
  NAND2_X1 U866 ( .A1(G141), .A2(n517), .ZN(n780) );
  NAND2_X1 U867 ( .A1(G129), .A2(n881), .ZN(n779) );
  NAND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n783) );
  NAND2_X1 U869 ( .A1(n886), .A2(G105), .ZN(n781) );
  XOR2_X1 U870 ( .A(KEYINPUT38), .B(n781), .Z(n782) );
  NOR2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n882), .A2(G117), .ZN(n784) );
  NAND2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n877) );
  NOR2_X1 U874 ( .A1(G1996), .A2(n877), .ZN(n926) );
  NOR2_X1 U875 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U876 ( .A(n788), .B(KEYINPUT88), .ZN(n824) );
  AND2_X1 U877 ( .A1(n877), .A2(G1996), .ZN(n798) );
  NAND2_X1 U878 ( .A1(G107), .A2(n882), .ZN(n789) );
  XNOR2_X1 U879 ( .A(n789), .B(KEYINPUT90), .ZN(n792) );
  NAND2_X1 U880 ( .A1(G119), .A2(n881), .ZN(n790) );
  XOR2_X1 U881 ( .A(KEYINPUT89), .B(n790), .Z(n791) );
  NAND2_X1 U882 ( .A1(n792), .A2(n791), .ZN(n796) );
  NAND2_X1 U883 ( .A1(G131), .A2(n517), .ZN(n794) );
  NAND2_X1 U884 ( .A1(G95), .A2(n886), .ZN(n793) );
  NAND2_X1 U885 ( .A1(n794), .A2(n793), .ZN(n795) );
  OR2_X1 U886 ( .A1(n796), .A2(n795), .ZN(n892) );
  AND2_X1 U887 ( .A1(n892), .A2(G1991), .ZN(n797) );
  NOR2_X1 U888 ( .A1(n798), .A2(n797), .ZN(n924) );
  INV_X1 U889 ( .A(n924), .ZN(n799) );
  NAND2_X1 U890 ( .A1(n824), .A2(n799), .ZN(n823) );
  INV_X1 U891 ( .A(n823), .ZN(n802) );
  NOR2_X1 U892 ( .A1(G1991), .A2(n892), .ZN(n922) );
  NOR2_X1 U893 ( .A1(G1986), .A2(G290), .ZN(n800) );
  NOR2_X1 U894 ( .A1(n922), .A2(n800), .ZN(n801) );
  NOR2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U896 ( .A1(n926), .A2(n803), .ZN(n804) );
  XNOR2_X1 U897 ( .A(n805), .B(n804), .ZN(n815) );
  XNOR2_X1 U898 ( .A(KEYINPUT37), .B(G2067), .ZN(n816) );
  NAND2_X1 U899 ( .A1(G140), .A2(n517), .ZN(n807) );
  NAND2_X1 U900 ( .A1(G104), .A2(n886), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U902 ( .A(KEYINPUT34), .B(n808), .ZN(n813) );
  NAND2_X1 U903 ( .A1(G128), .A2(n881), .ZN(n810) );
  NAND2_X1 U904 ( .A1(G116), .A2(n882), .ZN(n809) );
  NAND2_X1 U905 ( .A1(n810), .A2(n809), .ZN(n811) );
  XOR2_X1 U906 ( .A(KEYINPUT35), .B(n811), .Z(n812) );
  NOR2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U908 ( .A(KEYINPUT36), .B(n814), .ZN(n878) );
  NOR2_X1 U909 ( .A1(n816), .A2(n878), .ZN(n933) );
  NAND2_X1 U910 ( .A1(n933), .A2(n824), .ZN(n822) );
  NAND2_X1 U911 ( .A1(n815), .A2(n822), .ZN(n817) );
  NAND2_X1 U912 ( .A1(n816), .A2(n878), .ZN(n937) );
  NAND2_X1 U913 ( .A1(n817), .A2(n937), .ZN(n818) );
  AND2_X1 U914 ( .A1(n818), .A2(n824), .ZN(n828) );
  OR2_X1 U915 ( .A1(n819), .A2(n828), .ZN(n820) );
  NOR2_X1 U916 ( .A1(n821), .A2(n820), .ZN(n830) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n826) );
  XNOR2_X1 U918 ( .A(G1986), .B(G290), .ZN(n969) );
  AND2_X1 U919 ( .A1(n969), .A2(n824), .ZN(n825) );
  NOR2_X1 U920 ( .A1(n826), .A2(n825), .ZN(n827) );
  NOR2_X1 U921 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U922 ( .A(n831), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n915), .ZN(G217) );
  NAND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n832) );
  XNOR2_X1 U925 ( .A(KEYINPUT103), .B(n832), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n833), .A2(G661), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U928 ( .A1(n835), .A2(n834), .ZN(G188) );
  XOR2_X1 U929 ( .A(G1971), .B(G1956), .Z(n837) );
  XNOR2_X1 U930 ( .A(G1996), .B(G1991), .ZN(n836) );
  XNOR2_X1 U931 ( .A(n837), .B(n836), .ZN(n847) );
  XOR2_X1 U932 ( .A(G2474), .B(KEYINPUT41), .Z(n839) );
  XNOR2_X1 U933 ( .A(G1961), .B(KEYINPUT107), .ZN(n838) );
  XNOR2_X1 U934 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U935 ( .A(G1976), .B(G1966), .Z(n841) );
  XNOR2_X1 U936 ( .A(G1986), .B(G1981), .ZN(n840) );
  XNOR2_X1 U937 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U938 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U939 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n844) );
  XNOR2_X1 U940 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U941 ( .A(n847), .B(n846), .Z(G229) );
  XOR2_X1 U942 ( .A(G2096), .B(KEYINPUT43), .Z(n849) );
  XNOR2_X1 U943 ( .A(G2072), .B(KEYINPUT104), .ZN(n848) );
  XNOR2_X1 U944 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U945 ( .A(n850), .B(G2678), .Z(n852) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2090), .ZN(n851) );
  XNOR2_X1 U947 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U948 ( .A(KEYINPUT42), .B(G2100), .Z(n854) );
  XNOR2_X1 U949 ( .A(G2084), .B(G2078), .ZN(n853) );
  XNOR2_X1 U950 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U951 ( .A(n856), .B(n855), .ZN(G227) );
  INV_X1 U952 ( .A(n857), .ZN(G319) );
  NAND2_X1 U953 ( .A1(G136), .A2(n517), .ZN(n858) );
  XNOR2_X1 U954 ( .A(n858), .B(KEYINPUT108), .ZN(n865) );
  NAND2_X1 U955 ( .A1(G100), .A2(n886), .ZN(n860) );
  NAND2_X1 U956 ( .A1(G112), .A2(n882), .ZN(n859) );
  NAND2_X1 U957 ( .A1(n860), .A2(n859), .ZN(n863) );
  NAND2_X1 U958 ( .A1(n881), .A2(G124), .ZN(n861) );
  XOR2_X1 U959 ( .A(KEYINPUT44), .B(n861), .Z(n862) );
  NOR2_X1 U960 ( .A1(n863), .A2(n862), .ZN(n864) );
  NAND2_X1 U961 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U962 ( .A(KEYINPUT109), .B(n866), .ZN(G162) );
  NAND2_X1 U963 ( .A1(G139), .A2(n517), .ZN(n868) );
  NAND2_X1 U964 ( .A1(G103), .A2(n886), .ZN(n867) );
  NAND2_X1 U965 ( .A1(n868), .A2(n867), .ZN(n873) );
  NAND2_X1 U966 ( .A1(G127), .A2(n881), .ZN(n870) );
  NAND2_X1 U967 ( .A1(G115), .A2(n882), .ZN(n869) );
  NAND2_X1 U968 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U969 ( .A(KEYINPUT47), .B(n871), .Z(n872) );
  NOR2_X1 U970 ( .A1(n873), .A2(n872), .ZN(n916) );
  XOR2_X1 U971 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n875) );
  XNOR2_X1 U972 ( .A(KEYINPUT111), .B(KEYINPUT110), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n916), .B(n876), .ZN(n880) );
  XOR2_X1 U975 ( .A(n878), .B(n877), .Z(n879) );
  XNOR2_X1 U976 ( .A(n880), .B(n879), .ZN(n895) );
  NAND2_X1 U977 ( .A1(G130), .A2(n881), .ZN(n884) );
  NAND2_X1 U978 ( .A1(G118), .A2(n882), .ZN(n883) );
  NAND2_X1 U979 ( .A1(n884), .A2(n883), .ZN(n891) );
  NAND2_X1 U980 ( .A1(G142), .A2(n517), .ZN(n888) );
  NAND2_X1 U981 ( .A1(G106), .A2(n886), .ZN(n887) );
  NAND2_X1 U982 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U983 ( .A(n889), .B(KEYINPUT45), .Z(n890) );
  NOR2_X1 U984 ( .A1(n891), .A2(n890), .ZN(n893) );
  XNOR2_X1 U985 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U986 ( .A(n895), .B(n894), .Z(n897) );
  XNOR2_X1 U987 ( .A(G164), .B(G160), .ZN(n896) );
  XNOR2_X1 U988 ( .A(n897), .B(n896), .ZN(n899) );
  XOR2_X1 U989 ( .A(n923), .B(G162), .Z(n898) );
  XNOR2_X1 U990 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U991 ( .A1(G37), .A2(n900), .ZN(G395) );
  XNOR2_X1 U992 ( .A(n901), .B(n974), .ZN(n902) );
  XOR2_X1 U993 ( .A(n902), .B(n970), .Z(n904) );
  XOR2_X1 U994 ( .A(G286), .B(G171), .Z(n903) );
  XNOR2_X1 U995 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U996 ( .A1(G37), .A2(n905), .ZN(G397) );
  NOR2_X1 U997 ( .A1(G229), .A2(G227), .ZN(n906) );
  XOR2_X1 U998 ( .A(KEYINPUT112), .B(n906), .Z(n907) );
  XNOR2_X1 U999 ( .A(KEYINPUT49), .B(n907), .ZN(n912) );
  NOR2_X1 U1000 ( .A1(G395), .A2(G397), .ZN(n908) );
  XOR2_X1 U1001 ( .A(KEYINPUT113), .B(n908), .Z(n909) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n909), .ZN(n910) );
  NOR2_X1 U1003 ( .A1(G401), .A2(n910), .ZN(n911) );
  NAND2_X1 U1004 ( .A1(n912), .A2(n911), .ZN(G225) );
  XOR2_X1 U1005 ( .A(KEYINPUT114), .B(G225), .Z(G308) );
  INV_X1 U1007 ( .A(G120), .ZN(G236) );
  INV_X1 U1008 ( .A(G108), .ZN(G238) );
  INV_X1 U1009 ( .A(G96), .ZN(G221) );
  INV_X1 U1010 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(G325) );
  INV_X1 U1012 ( .A(G325), .ZN(G261) );
  INV_X1 U1013 ( .A(n915), .ZN(G223) );
  XNOR2_X1 U1014 ( .A(KEYINPUT116), .B(KEYINPUT50), .ZN(n920) );
  XNOR2_X1 U1015 ( .A(G2072), .B(n916), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(G164), .B(G2078), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1018 ( .A(n920), .B(n919), .ZN(n936) );
  XOR2_X1 U1019 ( .A(G160), .B(G2084), .Z(n921) );
  NOR2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n931) );
  NAND2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n929) );
  XOR2_X1 U1022 ( .A(G2090), .B(G162), .Z(n925) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(n927), .B(KEYINPUT51), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1028 ( .A(n934), .B(KEYINPUT115), .ZN(n935) );
  NOR2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n938) );
  NAND2_X1 U1030 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1031 ( .A(KEYINPUT52), .B(n939), .ZN(n940) );
  NAND2_X1 U1032 ( .A1(n940), .A2(G29), .ZN(n1023) );
  XNOR2_X1 U1033 ( .A(G2084), .B(G34), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(n941), .B(KEYINPUT54), .ZN(n959) );
  XOR2_X1 U1035 ( .A(G2090), .B(G35), .Z(n957) );
  XNOR2_X1 U1036 ( .A(G27), .B(n942), .ZN(n946) );
  XNOR2_X1 U1037 ( .A(G2067), .B(G26), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(G32), .B(G1996), .ZN(n943) );
  NOR2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n949) );
  XOR2_X1 U1041 ( .A(KEYINPUT117), .B(G2072), .Z(n947) );
  XNOR2_X1 U1042 ( .A(G33), .B(n947), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1044 ( .A(KEYINPUT118), .B(n950), .Z(n952) );
  XNOR2_X1 U1045 ( .A(G1991), .B(G25), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n953), .A2(G28), .ZN(n954) );
  XOR2_X1 U1048 ( .A(KEYINPUT53), .B(n954), .Z(n955) );
  XNOR2_X1 U1049 ( .A(n955), .B(KEYINPUT119), .ZN(n956) );
  NAND2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(n960), .B(KEYINPUT120), .ZN(n961) );
  NOR2_X1 U1053 ( .A1(G29), .A2(n961), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(KEYINPUT55), .B(n962), .ZN(n963) );
  NAND2_X1 U1055 ( .A1(n963), .A2(G11), .ZN(n1021) );
  INV_X1 U1056 ( .A(G16), .ZN(n1017) );
  XOR2_X1 U1057 ( .A(n1017), .B(KEYINPUT56), .Z(n990) );
  XOR2_X1 U1058 ( .A(G168), .B(G1966), .Z(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1060 ( .A(KEYINPUT57), .B(n966), .Z(n988) );
  XOR2_X1 U1061 ( .A(G1956), .B(n967), .Z(n968) );
  NOR2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n973) );
  XNOR2_X1 U1063 ( .A(G1348), .B(KEYINPUT121), .ZN(n971) );
  XOR2_X1 U1064 ( .A(n971), .B(n970), .Z(n972) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n977) );
  XOR2_X1 U1066 ( .A(G1341), .B(n974), .Z(n975) );
  XNOR2_X1 U1067 ( .A(KEYINPUT123), .B(n975), .ZN(n976) );
  NOR2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n984) );
  AND2_X1 U1069 ( .A1(G303), .A2(G1971), .ZN(n981) );
  NAND2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1072 ( .A(n982), .B(KEYINPUT122), .ZN(n983) );
  NAND2_X1 U1073 ( .A1(n984), .A2(n983), .ZN(n986) );
  XOR2_X1 U1074 ( .A(G1961), .B(G171), .Z(n985) );
  NOR2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1077 ( .A1(n990), .A2(n989), .ZN(n1019) );
  XOR2_X1 U1078 ( .A(G1986), .B(G24), .Z(n994) );
  XNOR2_X1 U1079 ( .A(G1971), .B(G22), .ZN(n992) );
  XNOR2_X1 U1080 ( .A(G23), .B(G1976), .ZN(n991) );
  NOR2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(KEYINPUT58), .B(KEYINPUT127), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(n996), .B(n995), .ZN(n1012) );
  XNOR2_X1 U1085 ( .A(KEYINPUT125), .B(G1341), .ZN(n997) );
  XNOR2_X1 U1086 ( .A(n997), .B(G19), .ZN(n1003) );
  XOR2_X1 U1087 ( .A(G4), .B(KEYINPUT126), .Z(n999) );
  XNOR2_X1 U1088 ( .A(G1348), .B(KEYINPUT59), .ZN(n998) );
  XNOR2_X1 U1089 ( .A(n999), .B(n998), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(G1981), .B(G6), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1007) );
  XOR2_X1 U1093 ( .A(G20), .B(n1004), .Z(n1005) );
  XNOR2_X1 U1094 ( .A(KEYINPUT124), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1096 ( .A(KEYINPUT60), .B(n1008), .Z(n1010) );
  XNOR2_X1 U1097 ( .A(G1966), .B(G21), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(G5), .B(G1961), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1015), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1024), .ZN(G150) );
  INV_X1 U1108 ( .A(G150), .ZN(G311) );
endmodule

