

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755;

  INV_X1 U371 ( .A(KEYINPUT1), .ZN(n351) );
  XNOR2_X1 U372 ( .A(n502), .B(n501), .ZN(n742) );
  XNOR2_X1 U373 ( .A(n500), .B(G134), .ZN(n502) );
  BUF_X1 U374 ( .A(G107), .Z(n349) );
  XNOR2_X1 U375 ( .A(n437), .B(KEYINPUT69), .ZN(n522) );
  XNOR2_X1 U376 ( .A(n444), .B(n443), .ZN(n473) );
  INV_X1 U377 ( .A(G146), .ZN(n503) );
  INV_X2 U378 ( .A(G953), .ZN(n745) );
  NAND2_X1 U379 ( .A1(n350), .A2(n645), .ZN(n571) );
  XNOR2_X1 U380 ( .A(n558), .B(KEYINPUT85), .ZN(n350) );
  XNOR2_X1 U381 ( .A(n568), .B(KEYINPUT35), .ZN(n645) );
  INV_X1 U382 ( .A(n563), .ZN(n535) );
  NAND2_X1 U383 ( .A1(n563), .A2(n685), .ZN(n572) );
  XNOR2_X2 U384 ( .A(n590), .B(n351), .ZN(n563) );
  AND2_X2 U385 ( .A1(n620), .A2(n619), .ZN(n743) );
  NAND2_X1 U386 ( .A1(n352), .A2(n397), .ZN(n404) );
  NAND2_X1 U387 ( .A1(n400), .A2(n401), .ZN(n352) );
  NOR2_X1 U388 ( .A1(n560), .A2(n559), .ZN(n562) );
  XNOR2_X2 U389 ( .A(n520), .B(n521), .ZN(n560) );
  XNOR2_X2 U390 ( .A(G101), .B(KEYINPUT68), .ZN(n437) );
  XNOR2_X2 U391 ( .A(n478), .B(KEYINPUT71), .ZN(n500) );
  XNOR2_X2 U392 ( .A(n499), .B(KEYINPUT22), .ZN(n555) );
  XNOR2_X1 U393 ( .A(n423), .B(n422), .ZN(n755) );
  NAND2_X1 U394 ( .A1(n361), .A2(n395), .ZN(n394) );
  AND2_X1 U395 ( .A1(n743), .A2(n494), .ZN(n413) );
  XNOR2_X1 U396 ( .A(n407), .B(KEYINPUT41), .ZN(n709) );
  XNOR2_X1 U397 ( .A(n591), .B(KEYINPUT30), .ZN(n373) );
  XNOR2_X1 U398 ( .A(n688), .B(n532), .ZN(n564) );
  OR2_X1 U399 ( .A1(n623), .A2(G902), .ZN(n409) );
  OR2_X1 U400 ( .A1(n722), .A2(G902), .ZN(n520) );
  XOR2_X1 U401 ( .A(KEYINPUT62), .B(n623), .Z(n624) );
  XNOR2_X1 U402 ( .A(n436), .B(n726), .ZN(n507) );
  XNOR2_X2 U403 ( .A(G116), .B(G107), .ZN(n444) );
  XNOR2_X2 U404 ( .A(n742), .B(n503), .ZN(n530) );
  NOR2_X1 U405 ( .A1(n605), .A2(n381), .ZN(n380) );
  XNOR2_X1 U406 ( .A(n446), .B(KEYINPUT3), .ZN(n523) );
  XNOR2_X1 U407 ( .A(G119), .B(G113), .ZN(n446) );
  AND2_X1 U408 ( .A1(n368), .A2(n367), .ZN(n366) );
  NAND2_X1 U409 ( .A1(n365), .A2(n622), .ZN(n364) );
  NOR2_X1 U410 ( .A1(n583), .A2(n566), .ZN(n606) );
  INV_X1 U411 ( .A(G237), .ZN(n454) );
  NAND2_X1 U412 ( .A1(n435), .A2(G902), .ZN(n433) );
  NOR2_X1 U413 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U414 ( .A(n406), .B(n615), .ZN(n620) );
  NAND2_X1 U415 ( .A1(n404), .A2(n402), .ZN(n406) );
  NOR2_X1 U416 ( .A1(n379), .A2(n376), .ZN(n402) );
  XNOR2_X1 U417 ( .A(n528), .B(n522), .ZN(n412) );
  XNOR2_X1 U418 ( .A(G116), .B(G137), .ZN(n526) );
  INV_X1 U419 ( .A(n523), .ZN(n411) );
  XNOR2_X1 U420 ( .A(n491), .B(n490), .ZN(n631) );
  XNOR2_X1 U421 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U422 ( .A(n530), .B(n508), .ZN(n715) );
  XNOR2_X1 U423 ( .A(n507), .B(n506), .ZN(n508) );
  NAND2_X1 U424 ( .A1(n386), .A2(KEYINPUT2), .ZN(n420) );
  INV_X1 U425 ( .A(n408), .ZN(n386) );
  XNOR2_X1 U426 ( .A(n360), .B(n419), .ZN(n637) );
  XNOR2_X1 U427 ( .A(n725), .B(n507), .ZN(n360) );
  INV_X1 U428 ( .A(n420), .ZN(n706) );
  INV_X1 U429 ( .A(KEYINPUT108), .ZN(n549) );
  OR2_X1 U430 ( .A1(n674), .A2(n676), .ZN(n407) );
  INV_X1 U431 ( .A(n373), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n426), .B(n424), .ZN(n519) );
  XNOR2_X1 U433 ( .A(n516), .B(n513), .ZN(n426) );
  NAND2_X1 U434 ( .A1(n512), .A2(G221), .ZN(n424) );
  XNOR2_X1 U435 ( .A(n378), .B(n377), .ZN(n376) );
  INV_X1 U436 ( .A(KEYINPUT81), .ZN(n377) );
  NAND2_X1 U437 ( .A1(n456), .A2(n494), .ZN(n367) );
  INV_X1 U438 ( .A(KEYINPUT44), .ZN(n570) );
  XOR2_X1 U439 ( .A(G140), .B(G122), .Z(n477) );
  XNOR2_X1 U440 ( .A(G143), .B(G104), .ZN(n486) );
  AND2_X1 U441 ( .A1(n374), .A2(n494), .ZN(n389) );
  NAND2_X1 U442 ( .A1(n375), .A2(n704), .ZN(n374) );
  XNOR2_X1 U443 ( .A(n522), .B(KEYINPUT74), .ZN(n436) );
  NAND2_X1 U444 ( .A1(G234), .A2(G237), .ZN(n458) );
  AND2_X1 U445 ( .A1(n672), .A2(n592), .ZN(n372) );
  XNOR2_X1 U446 ( .A(n543), .B(KEYINPUT73), .ZN(n589) );
  INV_X1 U447 ( .A(KEYINPUT70), .ZN(n561) );
  OR2_X2 U448 ( .A1(n432), .A2(n429), .ZN(n590) );
  NAND2_X1 U449 ( .A1(n434), .A2(n433), .ZN(n432) );
  NAND2_X1 U450 ( .A1(G469), .A2(n431), .ZN(n430) );
  XNOR2_X1 U451 ( .A(n447), .B(n523), .ZN(n725) );
  INV_X1 U452 ( .A(KEYINPUT16), .ZN(n445) );
  XNOR2_X1 U453 ( .A(n466), .B(n425), .ZN(n512) );
  INV_X1 U454 ( .A(KEYINPUT8), .ZN(n425) );
  XNOR2_X1 U455 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U456 ( .A(G128), .B(G119), .ZN(n515) );
  XOR2_X1 U457 ( .A(G110), .B(KEYINPUT23), .Z(n513) );
  XNOR2_X1 U458 ( .A(G143), .B(G128), .ZN(n470) );
  NAND2_X1 U459 ( .A1(n608), .A2(n671), .ZN(n369) );
  AND2_X1 U460 ( .A1(n383), .A2(n382), .ZN(n609) );
  INV_X1 U461 ( .A(n590), .ZN(n382) );
  XNOR2_X1 U462 ( .A(n385), .B(n384), .ZN(n383) );
  INV_X1 U463 ( .A(KEYINPUT28), .ZN(n384) );
  XNOR2_X1 U464 ( .A(n574), .B(KEYINPUT93), .ZN(n578) );
  XNOR2_X1 U465 ( .A(n410), .B(n525), .ZN(n529) );
  XNOR2_X1 U466 ( .A(n412), .B(n411), .ZN(n410) );
  XNOR2_X1 U467 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U468 ( .A(n637), .B(n638), .ZN(n639) );
  NOR2_X1 U469 ( .A1(n712), .A2(n711), .ZN(n713) );
  AND2_X1 U470 ( .A1(n414), .A2(n599), .ZN(n618) );
  NOR2_X1 U471 ( .A1(n548), .A2(n684), .ZN(n415) );
  INV_X1 U472 ( .A(KEYINPUT40), .ZN(n422) );
  AND2_X1 U473 ( .A1(n462), .A2(n609), .ZN(n658) );
  XNOR2_X1 U474 ( .A(n723), .B(n722), .ZN(n362) );
  XNOR2_X1 U475 ( .A(n720), .B(n719), .ZN(n391) );
  XNOR2_X1 U476 ( .A(n393), .B(n359), .ZN(n392) );
  XNOR2_X1 U477 ( .A(n417), .B(n416), .ZN(G75) );
  XNOR2_X1 U478 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n416) );
  NAND2_X1 U479 ( .A1(n713), .A2(n418), .ZN(n417) );
  AND2_X1 U480 ( .A1(n714), .A2(n745), .ZN(n418) );
  AND2_X1 U481 ( .A1(n619), .A2(KEYINPUT82), .ZN(n353) );
  INV_X1 U482 ( .A(G469), .ZN(n435) );
  AND2_X1 U483 ( .A1(n420), .A2(G210), .ZN(n354) );
  AND2_X1 U484 ( .A1(n595), .A2(n372), .ZN(n355) );
  AND2_X1 U485 ( .A1(n420), .A2(G475), .ZN(n356) );
  INV_X1 U486 ( .A(G902), .ZN(n431) );
  XOR2_X1 U487 ( .A(KEYINPUT87), .B(KEYINPUT33), .Z(n357) );
  NAND2_X2 U488 ( .A1(n366), .A2(n363), .ZN(n608) );
  XOR2_X1 U489 ( .A(n550), .B(n549), .Z(n358) );
  XOR2_X1 U490 ( .A(n717), .B(n716), .Z(n359) );
  XNOR2_X1 U491 ( .A(G902), .B(KEYINPUT15), .ZN(n622) );
  NAND2_X1 U492 ( .A1(n387), .A2(n389), .ZN(n361) );
  NOR2_X1 U493 ( .A1(n362), .A2(n724), .ZN(G66) );
  OR2_X1 U494 ( .A1(n637), .A2(n364), .ZN(n363) );
  INV_X1 U495 ( .A(n456), .ZN(n365) );
  NAND2_X1 U496 ( .A1(n637), .A2(n456), .ZN(n368) );
  XNOR2_X2 U497 ( .A(n369), .B(KEYINPUT19), .ZN(n462) );
  NOR2_X1 U498 ( .A1(n370), .A2(n373), .ZN(n612) );
  NAND2_X1 U499 ( .A1(n595), .A2(n592), .ZN(n370) );
  NAND2_X1 U500 ( .A1(n355), .A2(n371), .ZN(n613) );
  NAND2_X1 U501 ( .A1(n620), .A2(n353), .ZN(n375) );
  NAND2_X1 U502 ( .A1(n598), .A2(n656), .ZN(n378) );
  NAND2_X1 U503 ( .A1(n380), .A2(n403), .ZN(n379) );
  INV_X1 U504 ( .A(n668), .ZN(n381) );
  NAND2_X1 U505 ( .A1(n589), .A2(n688), .ZN(n385) );
  INV_X1 U506 ( .A(n622), .ZN(n494) );
  NAND2_X1 U507 ( .A1(n622), .A2(G234), .ZN(n495) );
  NAND2_X1 U508 ( .A1(n388), .A2(n704), .ZN(n387) );
  INV_X1 U509 ( .A(n730), .ZN(n388) );
  XNOR2_X2 U510 ( .A(n588), .B(KEYINPUT45), .ZN(n730) );
  NAND2_X1 U511 ( .A1(n421), .A2(n354), .ZN(n640) );
  AND2_X2 U512 ( .A1(n421), .A2(n420), .ZN(n721) );
  NAND2_X1 U513 ( .A1(n421), .A2(n356), .ZN(n633) );
  NAND2_X1 U514 ( .A1(n421), .A2(n390), .ZN(n625) );
  AND2_X1 U515 ( .A1(n420), .A2(G472), .ZN(n390) );
  NOR2_X1 U516 ( .A1(n391), .A2(n724), .ZN(G63) );
  NOR2_X1 U517 ( .A1(n392), .A2(n724), .ZN(G54) );
  NAND2_X1 U518 ( .A1(n555), .A2(n440), .ZN(n438) );
  NAND2_X1 U519 ( .A1(n730), .A2(n743), .ZN(n408) );
  NAND2_X1 U520 ( .A1(n721), .A2(G469), .ZN(n393) );
  XNOR2_X2 U521 ( .A(n394), .B(KEYINPUT64), .ZN(n421) );
  NAND2_X1 U522 ( .A1(n396), .A2(n621), .ZN(n395) );
  NAND2_X1 U523 ( .A1(n413), .A2(n730), .ZN(n396) );
  NAND2_X1 U524 ( .A1(n754), .A2(n398), .ZN(n397) );
  INV_X1 U525 ( .A(n614), .ZN(n398) );
  INV_X1 U526 ( .A(n405), .ZN(n400) );
  INV_X1 U527 ( .A(n754), .ZN(n401) );
  NAND2_X1 U528 ( .A1(n755), .A2(n614), .ZN(n403) );
  NOR2_X1 U529 ( .A1(n755), .A2(n614), .ZN(n405) );
  NAND2_X1 U530 ( .A1(n609), .A2(n709), .ZN(n610) );
  NAND2_X1 U531 ( .A1(n672), .A2(n671), .ZN(n676) );
  NAND2_X1 U532 ( .A1(n408), .A2(n704), .ZN(n705) );
  NAND2_X1 U533 ( .A1(n589), .A2(n564), .ZN(n544) );
  XNOR2_X2 U534 ( .A(n409), .B(n531), .ZN(n688) );
  XNOR2_X1 U535 ( .A(n415), .B(n358), .ZN(n414) );
  XNOR2_X1 U536 ( .A(n452), .B(n501), .ZN(n419) );
  NOR2_X2 U537 ( .A1(n574), .A2(n498), .ZN(n499) );
  NAND2_X1 U538 ( .A1(n616), .A2(n657), .ZN(n423) );
  XNOR2_X2 U539 ( .A(n613), .B(KEYINPUT39), .ZN(n616) );
  NAND2_X1 U540 ( .A1(n708), .A2(n578), .ZN(n565) );
  XNOR2_X2 U541 ( .A(n465), .B(n464), .ZN(n574) );
  XNOR2_X2 U542 ( .A(n427), .B(n357), .ZN(n708) );
  NAND2_X1 U543 ( .A1(n428), .A2(n564), .ZN(n427) );
  XNOR2_X1 U544 ( .A(n572), .B(KEYINPUT103), .ZN(n428) );
  NAND2_X1 U545 ( .A1(n715), .A2(n435), .ZN(n434) );
  NOR2_X1 U546 ( .A1(n715), .A2(n430), .ZN(n429) );
  NAND2_X1 U547 ( .A1(n556), .A2(n557), .ZN(n558) );
  XNOR2_X2 U548 ( .A(n438), .B(KEYINPUT102), .ZN(n557) );
  XNOR2_X2 U549 ( .A(n439), .B(KEYINPUT32), .ZN(n556) );
  NAND2_X1 U550 ( .A1(n555), .A2(n554), .ZN(n439) );
  NOR2_X1 U551 ( .A1(n577), .A2(n590), .ZN(n594) );
  AND2_X1 U552 ( .A1(n536), .A2(n580), .ZN(n440) );
  OR2_X1 U553 ( .A1(n540), .A2(n461), .ZN(n441) );
  AND2_X1 U554 ( .A1(n586), .A2(n585), .ZN(n442) );
  XNOR2_X1 U555 ( .A(n477), .B(G113), .ZN(n479) );
  XNOR2_X1 U556 ( .A(KEYINPUT48), .B(KEYINPUT83), .ZN(n615) );
  XNOR2_X1 U557 ( .A(n479), .B(n500), .ZN(n480) );
  INV_X1 U558 ( .A(n671), .ZN(n545) );
  NOR2_X1 U559 ( .A1(n661), .A2(n545), .ZN(n546) );
  NAND2_X1 U560 ( .A1(n547), .A2(n546), .ZN(n600) );
  XNOR2_X1 U561 ( .A(n741), .B(n519), .ZN(n722) );
  AND2_X1 U562 ( .A1(n626), .A2(G953), .ZN(n724) );
  INV_X1 U563 ( .A(G122), .ZN(n443) );
  XNOR2_X1 U564 ( .A(n473), .B(n445), .ZN(n447) );
  NAND2_X1 U565 ( .A1(n745), .A2(G224), .ZN(n448) );
  XNOR2_X1 U566 ( .A(n448), .B(KEYINPUT90), .ZN(n450) );
  XNOR2_X1 U567 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n449) );
  XNOR2_X1 U568 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U569 ( .A(n503), .B(G125), .ZN(n481) );
  XNOR2_X1 U570 ( .A(n481), .B(n451), .ZN(n452) );
  XNOR2_X1 U571 ( .A(n470), .B(KEYINPUT4), .ZN(n501) );
  XOR2_X1 U572 ( .A(G104), .B(KEYINPUT89), .Z(n453) );
  XNOR2_X1 U573 ( .A(n453), .B(G110), .ZN(n726) );
  NAND2_X1 U574 ( .A1(n431), .A2(n454), .ZN(n457) );
  NAND2_X1 U575 ( .A1(n457), .A2(G210), .ZN(n455) );
  XNOR2_X1 U576 ( .A(n455), .B(KEYINPUT91), .ZN(n456) );
  NAND2_X1 U577 ( .A1(n457), .A2(G214), .ZN(n671) );
  XNOR2_X1 U578 ( .A(n458), .B(KEYINPUT14), .ZN(n460) );
  NAND2_X1 U579 ( .A1(G952), .A2(n460), .ZN(n702) );
  NOR2_X1 U580 ( .A1(n702), .A2(G953), .ZN(n540) );
  XNOR2_X1 U581 ( .A(KEYINPUT92), .B(G898), .ZN(n733) );
  AND2_X1 U582 ( .A1(G953), .A2(G902), .ZN(n459) );
  NAND2_X1 U583 ( .A1(n460), .A2(n459), .ZN(n537) );
  NOR2_X1 U584 ( .A1(n733), .A2(n537), .ZN(n461) );
  NAND2_X1 U585 ( .A1(n462), .A2(n441), .ZN(n465) );
  INV_X1 U586 ( .A(KEYINPUT67), .ZN(n463) );
  XNOR2_X1 U587 ( .A(n463), .B(KEYINPUT0), .ZN(n464) );
  XOR2_X1 U588 ( .A(G134), .B(KEYINPUT7), .Z(n468) );
  NAND2_X1 U589 ( .A1(G234), .A2(n745), .ZN(n466) );
  NAND2_X1 U590 ( .A1(G217), .A2(n512), .ZN(n467) );
  XNOR2_X1 U591 ( .A(n468), .B(n467), .ZN(n469) );
  XOR2_X1 U592 ( .A(n469), .B(KEYINPUT100), .Z(n472) );
  XOR2_X1 U593 ( .A(KEYINPUT9), .B(n470), .Z(n471) );
  XNOR2_X1 U594 ( .A(n472), .B(n471), .ZN(n474) );
  XNOR2_X1 U595 ( .A(n474), .B(n473), .ZN(n718) );
  NOR2_X1 U596 ( .A1(n718), .A2(G902), .ZN(n476) );
  INV_X1 U597 ( .A(G478), .ZN(n475) );
  XNOR2_X1 U598 ( .A(n476), .B(n475), .ZN(n583) );
  XNOR2_X1 U599 ( .A(KEYINPUT13), .B(G475), .ZN(n493) );
  XNOR2_X2 U600 ( .A(G131), .B(KEYINPUT72), .ZN(n478) );
  XOR2_X1 U601 ( .A(n480), .B(KEYINPUT11), .Z(n484) );
  XNOR2_X1 U602 ( .A(KEYINPUT10), .B(n481), .ZN(n517) );
  INV_X1 U603 ( .A(n517), .ZN(n482) );
  XNOR2_X1 U604 ( .A(n482), .B(KEYINPUT98), .ZN(n483) );
  XNOR2_X1 U605 ( .A(n484), .B(n483), .ZN(n491) );
  NOR2_X1 U606 ( .A1(G237), .A2(G953), .ZN(n485) );
  XNOR2_X1 U607 ( .A(n485), .B(KEYINPUT76), .ZN(n524) );
  NAND2_X1 U608 ( .A1(n524), .A2(G214), .ZN(n489) );
  XOR2_X1 U609 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n487) );
  XNOR2_X1 U610 ( .A(n487), .B(n486), .ZN(n488) );
  NOR2_X1 U611 ( .A1(G902), .A2(n631), .ZN(n492) );
  XNOR2_X1 U612 ( .A(n493), .B(n492), .ZN(n566) );
  XNOR2_X1 U613 ( .A(n495), .B(KEYINPUT20), .ZN(n496) );
  XNOR2_X1 U614 ( .A(KEYINPUT94), .B(n496), .ZN(n509) );
  AND2_X1 U615 ( .A1(n509), .A2(G221), .ZN(n497) );
  XNOR2_X1 U616 ( .A(n497), .B(KEYINPUT21), .ZN(n689) );
  NAND2_X1 U617 ( .A1(n606), .A2(n689), .ZN(n498) );
  XOR2_X1 U618 ( .A(G137), .B(G140), .Z(n518) );
  XOR2_X1 U619 ( .A(n349), .B(n518), .Z(n505) );
  NAND2_X1 U620 ( .A1(G227), .A2(n745), .ZN(n504) );
  XNOR2_X1 U621 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U622 ( .A(KEYINPUT25), .B(KEYINPUT77), .Z(n511) );
  NAND2_X1 U623 ( .A1(G217), .A2(n509), .ZN(n510) );
  XNOR2_X1 U624 ( .A(n511), .B(n510), .ZN(n521) );
  INV_X1 U625 ( .A(KEYINPUT24), .ZN(n514) );
  XNOR2_X1 U626 ( .A(n518), .B(n517), .ZN(n741) );
  INV_X1 U627 ( .A(n560), .ZN(n690) );
  NAND2_X1 U628 ( .A1(n535), .A2(n690), .ZN(n533) );
  NAND2_X1 U629 ( .A1(G210), .A2(n524), .ZN(n525) );
  XOR2_X1 U630 ( .A(KEYINPUT75), .B(KEYINPUT5), .Z(n527) );
  XNOR2_X1 U631 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U632 ( .A(n530), .B(n529), .ZN(n623) );
  XNOR2_X1 U633 ( .A(G472), .B(KEYINPUT96), .ZN(n531) );
  INV_X1 U634 ( .A(KEYINPUT6), .ZN(n532) );
  NOR2_X1 U635 ( .A1(n533), .A2(n564), .ZN(n534) );
  NAND2_X1 U636 ( .A1(n555), .A2(n534), .ZN(n585) );
  XNOR2_X1 U637 ( .A(n585), .B(G101), .ZN(G3) );
  BUF_X2 U638 ( .A(n563), .Z(n684) );
  NOR2_X1 U639 ( .A1(n684), .A2(n690), .ZN(n536) );
  INV_X1 U640 ( .A(n688), .ZN(n580) );
  XNOR2_X1 U641 ( .A(n557), .B(G110), .ZN(G12) );
  XNOR2_X1 U642 ( .A(n537), .B(KEYINPUT104), .ZN(n538) );
  NOR2_X1 U643 ( .A1(G900), .A2(n538), .ZN(n539) );
  NOR2_X1 U644 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U645 ( .A(KEYINPUT79), .B(n541), .ZN(n592) );
  AND2_X1 U646 ( .A1(n592), .A2(n560), .ZN(n542) );
  NAND2_X1 U647 ( .A1(n542), .A2(n689), .ZN(n543) );
  XNOR2_X1 U648 ( .A(n544), .B(KEYINPUT105), .ZN(n547) );
  INV_X1 U649 ( .A(n566), .ZN(n582) );
  OR2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n661) );
  XNOR2_X1 U651 ( .A(n600), .B(KEYINPUT106), .ZN(n548) );
  XNOR2_X1 U652 ( .A(KEYINPUT43), .B(KEYINPUT107), .ZN(n550) );
  XOR2_X1 U653 ( .A(G140), .B(n618), .Z(G42) );
  NAND2_X1 U654 ( .A1(n684), .A2(n560), .ZN(n551) );
  XOR2_X1 U655 ( .A(KEYINPUT101), .B(n551), .Z(n553) );
  XNOR2_X1 U656 ( .A(n564), .B(KEYINPUT78), .ZN(n552) );
  NOR2_X1 U657 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U658 ( .A(n556), .B(G119), .ZN(G21) );
  INV_X1 U659 ( .A(n689), .ZN(n559) );
  XNOR2_X1 U660 ( .A(n562), .B(n561), .ZN(n577) );
  INV_X1 U661 ( .A(n577), .ZN(n685) );
  XNOR2_X1 U662 ( .A(n565), .B(KEYINPUT34), .ZN(n567) );
  NAND2_X1 U663 ( .A1(n583), .A2(n566), .ZN(n596) );
  NOR2_X2 U664 ( .A1(n567), .A2(n596), .ZN(n568) );
  XNOR2_X1 U665 ( .A(n571), .B(n570), .ZN(n587) );
  NOR2_X1 U666 ( .A1(n580), .A2(n572), .ZN(n573) );
  XNOR2_X1 U667 ( .A(n573), .B(KEYINPUT97), .ZN(n695) );
  BUF_X1 U668 ( .A(n574), .Z(n575) );
  NOR2_X1 U669 ( .A1(n695), .A2(n575), .ZN(n576) );
  XNOR2_X1 U670 ( .A(n576), .B(KEYINPUT31), .ZN(n664) );
  NAND2_X1 U671 ( .A1(n594), .A2(n578), .ZN(n579) );
  XNOR2_X1 U672 ( .A(KEYINPUT95), .B(n579), .ZN(n581) );
  NAND2_X1 U673 ( .A1(n581), .A2(n580), .ZN(n649) );
  NAND2_X1 U674 ( .A1(n664), .A2(n649), .ZN(n584) );
  AND2_X1 U675 ( .A1(n583), .A2(n582), .ZN(n653) );
  INV_X1 U676 ( .A(n653), .ZN(n665) );
  NAND2_X1 U677 ( .A1(n661), .A2(n665), .ZN(n675) );
  NAND2_X1 U678 ( .A1(n584), .A2(n675), .ZN(n586) );
  NAND2_X1 U679 ( .A1(n587), .A2(n442), .ZN(n588) );
  NAND2_X1 U680 ( .A1(n658), .A2(n675), .ZN(n604) );
  NAND2_X1 U681 ( .A1(n604), .A2(KEYINPUT47), .ZN(n598) );
  NAND2_X1 U682 ( .A1(n671), .A2(n688), .ZN(n591) );
  INV_X1 U683 ( .A(KEYINPUT109), .ZN(n593) );
  XNOR2_X1 U684 ( .A(n594), .B(n593), .ZN(n595) );
  INV_X1 U685 ( .A(n608), .ZN(n599) );
  NOR2_X1 U686 ( .A1(n596), .A2(n599), .ZN(n597) );
  NAND2_X1 U687 ( .A1(n612), .A2(n597), .ZN(n656) );
  NOR2_X1 U688 ( .A1(n600), .A2(n599), .ZN(n602) );
  XNOR2_X1 U689 ( .A(KEYINPUT36), .B(KEYINPUT86), .ZN(n601) );
  XNOR2_X1 U690 ( .A(n602), .B(n601), .ZN(n603) );
  NAND2_X1 U691 ( .A1(n684), .A2(n603), .ZN(n668) );
  NOR2_X1 U692 ( .A1(KEYINPUT47), .A2(n604), .ZN(n605) );
  XOR2_X1 U693 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n611) );
  INV_X1 U694 ( .A(n606), .ZN(n674) );
  INV_X1 U695 ( .A(KEYINPUT38), .ZN(n607) );
  XNOR2_X1 U696 ( .A(n608), .B(n607), .ZN(n672) );
  XNOR2_X1 U697 ( .A(n611), .B(n610), .ZN(n754) );
  INV_X1 U698 ( .A(n661), .ZN(n657) );
  XNOR2_X1 U699 ( .A(KEYINPUT46), .B(KEYINPUT84), .ZN(n614) );
  NAND2_X1 U700 ( .A1(n616), .A2(n653), .ZN(n670) );
  INV_X1 U701 ( .A(n670), .ZN(n617) );
  INV_X1 U702 ( .A(KEYINPUT82), .ZN(n621) );
  INV_X1 U703 ( .A(KEYINPUT2), .ZN(n704) );
  XNOR2_X1 U704 ( .A(n625), .B(n624), .ZN(n627) );
  INV_X1 U705 ( .A(G952), .ZN(n626) );
  INV_X1 U706 ( .A(n724), .ZN(n641) );
  NAND2_X1 U707 ( .A1(n627), .A2(n641), .ZN(n628) );
  XNOR2_X1 U708 ( .A(n628), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U709 ( .A(KEYINPUT65), .B(KEYINPUT88), .Z(n629) );
  XNOR2_X1 U710 ( .A(n629), .B(KEYINPUT59), .ZN(n630) );
  XNOR2_X1 U711 ( .A(n633), .B(n632), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n634), .A2(n641), .ZN(n636) );
  XOR2_X1 U713 ( .A(KEYINPUT66), .B(KEYINPUT60), .Z(n635) );
  XNOR2_X1 U714 ( .A(n636), .B(n635), .ZN(G60) );
  XNOR2_X1 U715 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n638) );
  XNOR2_X1 U716 ( .A(n640), .B(n639), .ZN(n642) );
  NAND2_X1 U717 ( .A1(n642), .A2(n641), .ZN(n644) );
  INV_X1 U718 ( .A(KEYINPUT56), .ZN(n643) );
  XNOR2_X1 U719 ( .A(n644), .B(n643), .ZN(G51) );
  BUF_X1 U720 ( .A(n645), .Z(n646) );
  XNOR2_X1 U721 ( .A(n646), .B(G122), .ZN(G24) );
  NOR2_X1 U722 ( .A1(n661), .A2(n649), .ZN(n648) );
  XNOR2_X1 U723 ( .A(G104), .B(KEYINPUT111), .ZN(n647) );
  XNOR2_X1 U724 ( .A(n648), .B(n647), .ZN(G6) );
  NOR2_X1 U725 ( .A1(n665), .A2(n649), .ZN(n651) );
  XNOR2_X1 U726 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n650) );
  XNOR2_X1 U727 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U728 ( .A(n349), .B(n652), .ZN(G9) );
  XOR2_X1 U729 ( .A(G128), .B(KEYINPUT29), .Z(n655) );
  NAND2_X1 U730 ( .A1(n658), .A2(n653), .ZN(n654) );
  XNOR2_X1 U731 ( .A(n655), .B(n654), .ZN(G30) );
  XNOR2_X1 U732 ( .A(G143), .B(n656), .ZN(G45) );
  XNOR2_X1 U733 ( .A(G146), .B(KEYINPUT112), .ZN(n660) );
  NAND2_X1 U734 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U735 ( .A(n660), .B(n659), .ZN(G48) );
  NOR2_X1 U736 ( .A1(n661), .A2(n664), .ZN(n663) );
  XNOR2_X1 U737 ( .A(G113), .B(KEYINPUT113), .ZN(n662) );
  XNOR2_X1 U738 ( .A(n663), .B(n662), .ZN(G15) );
  NOR2_X1 U739 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U740 ( .A(G116), .B(n666), .Z(G18) );
  XOR2_X1 U741 ( .A(KEYINPUT114), .B(KEYINPUT37), .Z(n667) );
  XNOR2_X1 U742 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U743 ( .A(G125), .B(n669), .ZN(G27) );
  XNOR2_X1 U744 ( .A(G134), .B(n670), .ZN(G36) );
  INV_X1 U745 ( .A(n708), .ZN(n682) );
  NOR2_X1 U746 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U747 ( .A1(n674), .A2(n673), .ZN(n679) );
  INV_X1 U748 ( .A(n675), .ZN(n677) );
  NOR2_X1 U749 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U750 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U751 ( .A(KEYINPUT115), .B(n680), .Z(n681) );
  NOR2_X1 U752 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U753 ( .A(KEYINPUT116), .B(n683), .Z(n699) );
  NOR2_X1 U754 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U755 ( .A(n686), .B(KEYINPUT50), .ZN(n687) );
  NOR2_X1 U756 ( .A1(n688), .A2(n687), .ZN(n693) );
  NOR2_X1 U757 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U758 ( .A(n691), .B(KEYINPUT49), .ZN(n692) );
  NAND2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U760 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U761 ( .A(KEYINPUT51), .B(n696), .Z(n697) );
  NAND2_X1 U762 ( .A1(n709), .A2(n697), .ZN(n698) );
  NAND2_X1 U763 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U764 ( .A(KEYINPUT52), .B(n700), .Z(n701) );
  NOR2_X1 U765 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U766 ( .A(KEYINPUT117), .B(n703), .ZN(n714) );
  XOR2_X1 U767 ( .A(KEYINPUT80), .B(n705), .Z(n707) );
  NOR2_X1 U768 ( .A1(n707), .A2(n706), .ZN(n712) );
  NAND2_X1 U769 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U770 ( .A(KEYINPUT118), .B(n710), .Z(n711) );
  XNOR2_X1 U771 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n717) );
  XNOR2_X1 U772 ( .A(n715), .B(KEYINPUT57), .ZN(n716) );
  NAND2_X1 U773 ( .A1(n721), .A2(G478), .ZN(n720) );
  XOR2_X1 U774 ( .A(n718), .B(KEYINPUT121), .Z(n719) );
  NAND2_X1 U775 ( .A1(n721), .A2(G217), .ZN(n723) );
  XNOR2_X1 U776 ( .A(n725), .B(G101), .ZN(n727) );
  XNOR2_X1 U777 ( .A(n727), .B(n726), .ZN(n729) );
  NOR2_X1 U778 ( .A1(n745), .A2(n733), .ZN(n728) );
  NOR2_X1 U779 ( .A1(n729), .A2(n728), .ZN(n739) );
  NAND2_X1 U780 ( .A1(n730), .A2(n745), .ZN(n731) );
  XNOR2_X1 U781 ( .A(n731), .B(KEYINPUT123), .ZN(n737) );
  NAND2_X1 U782 ( .A1(G953), .A2(G224), .ZN(n732) );
  XNOR2_X1 U783 ( .A(n732), .B(KEYINPUT61), .ZN(n734) );
  NAND2_X1 U784 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U785 ( .A(n735), .B(KEYINPUT122), .Z(n736) );
  NOR2_X1 U786 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U787 ( .A(n739), .B(n738), .Z(n740) );
  XNOR2_X1 U788 ( .A(KEYINPUT124), .B(n740), .ZN(G69) );
  XNOR2_X1 U789 ( .A(n742), .B(n741), .ZN(n748) );
  XNOR2_X1 U790 ( .A(n748), .B(n743), .ZN(n744) );
  XNOR2_X1 U791 ( .A(n744), .B(KEYINPUT125), .ZN(n746) );
  NAND2_X1 U792 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U793 ( .A(KEYINPUT126), .B(n747), .ZN(n753) );
  XNOR2_X1 U794 ( .A(G227), .B(n748), .ZN(n749) );
  NAND2_X1 U795 ( .A1(n749), .A2(G900), .ZN(n750) );
  NAND2_X1 U796 ( .A1(G953), .A2(n750), .ZN(n751) );
  XOR2_X1 U797 ( .A(KEYINPUT127), .B(n751), .Z(n752) );
  NAND2_X1 U798 ( .A1(n753), .A2(n752), .ZN(G72) );
  XOR2_X1 U799 ( .A(G137), .B(n754), .Z(G39) );
  XOR2_X1 U800 ( .A(n755), .B(G131), .Z(G33) );
endmodule

