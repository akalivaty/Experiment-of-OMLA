

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U559 ( .A1(G651), .A2(n583), .ZN(n806) );
  INV_X2 U560 ( .A(n636), .ZN(n524) );
  XNOR2_X1 U561 ( .A(n606), .B(n605), .ZN(n607) );
  XOR2_X1 U562 ( .A(KEYINPUT71), .B(n618), .Z(n525) );
  XNOR2_X1 U563 ( .A(KEYINPUT73), .B(n624), .ZN(n526) );
  XNOR2_X1 U564 ( .A(n675), .B(n628), .ZN(n636) );
  NOR2_X1 U565 ( .A1(n988), .A2(n642), .ZN(n643) );
  INV_X1 U566 ( .A(KEYINPUT72), .ZN(n620) );
  AND2_X1 U567 ( .A1(n625), .A2(n526), .ZN(n626) );
  XNOR2_X1 U568 ( .A(KEYINPUT13), .B(KEYINPUT70), .ZN(n605) );
  NOR2_X2 U569 ( .A1(n547), .A2(n583), .ZN(n802) );
  NOR2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  XOR2_X1 U571 ( .A(KEYINPUT17), .B(n527), .Z(n536) );
  NAND2_X1 U572 ( .A1(n536), .A2(G137), .ZN(n530) );
  INV_X1 U573 ( .A(G2104), .ZN(n531) );
  NOR2_X4 U574 ( .A1(G2105), .A2(n531), .ZN(n890) );
  NAND2_X1 U575 ( .A1(G101), .A2(n890), .ZN(n528) );
  XOR2_X1 U576 ( .A(KEYINPUT23), .B(n528), .Z(n529) );
  NAND2_X1 U577 ( .A1(n530), .A2(n529), .ZN(n535) );
  AND2_X1 U578 ( .A1(G2104), .A2(G2105), .ZN(n886) );
  NAND2_X1 U579 ( .A1(G113), .A2(n886), .ZN(n533) );
  AND2_X1 U580 ( .A1(n531), .A2(G2105), .ZN(n887) );
  NAND2_X1 U581 ( .A1(G125), .A2(n887), .ZN(n532) );
  NAND2_X1 U582 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X2 U583 ( .A1(n535), .A2(n534), .ZN(G160) );
  BUF_X1 U584 ( .A(n536), .Z(n891) );
  NAND2_X1 U585 ( .A1(n891), .A2(G138), .ZN(n539) );
  NAND2_X1 U586 ( .A1(G114), .A2(n886), .ZN(n537) );
  XOR2_X1 U587 ( .A(KEYINPUT83), .B(n537), .Z(n538) );
  NAND2_X1 U588 ( .A1(n539), .A2(n538), .ZN(n543) );
  NAND2_X1 U589 ( .A1(G102), .A2(n890), .ZN(n541) );
  NAND2_X1 U590 ( .A1(G126), .A2(n887), .ZN(n540) );
  NAND2_X1 U591 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U592 ( .A1(n543), .A2(n542), .ZN(G164) );
  XOR2_X1 U593 ( .A(G543), .B(KEYINPUT0), .Z(n544) );
  XNOR2_X1 U594 ( .A(KEYINPUT64), .B(n544), .ZN(n583) );
  NAND2_X1 U595 ( .A1(n806), .A2(G53), .ZN(n553) );
  INV_X1 U596 ( .A(G651), .ZN(n547) );
  NAND2_X1 U597 ( .A1(G78), .A2(n802), .ZN(n546) );
  NOR2_X1 U598 ( .A1(G651), .A2(G543), .ZN(n805) );
  NAND2_X1 U599 ( .A1(G91), .A2(n805), .ZN(n545) );
  NAND2_X1 U600 ( .A1(n546), .A2(n545), .ZN(n551) );
  NOR2_X1 U601 ( .A1(G543), .A2(n547), .ZN(n548) );
  XOR2_X2 U602 ( .A(KEYINPUT1), .B(n548), .Z(n801) );
  NAND2_X1 U603 ( .A1(n801), .A2(G65), .ZN(n549) );
  XOR2_X1 U604 ( .A(KEYINPUT66), .B(n549), .Z(n550) );
  NOR2_X1 U605 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U606 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U607 ( .A(KEYINPUT67), .B(n554), .Z(G299) );
  NAND2_X1 U608 ( .A1(G64), .A2(n801), .ZN(n555) );
  XNOR2_X1 U609 ( .A(n555), .B(KEYINPUT65), .ZN(n562) );
  NAND2_X1 U610 ( .A1(G77), .A2(n802), .ZN(n557) );
  NAND2_X1 U611 ( .A1(G90), .A2(n805), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U613 ( .A(n558), .B(KEYINPUT9), .ZN(n560) );
  NAND2_X1 U614 ( .A1(G52), .A2(n806), .ZN(n559) );
  NAND2_X1 U615 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U616 ( .A1(n562), .A2(n561), .ZN(G171) );
  INV_X1 U617 ( .A(G171), .ZN(G301) );
  NAND2_X1 U618 ( .A1(n805), .A2(G89), .ZN(n563) );
  XNOR2_X1 U619 ( .A(n563), .B(KEYINPUT4), .ZN(n565) );
  NAND2_X1 U620 ( .A1(G76), .A2(n802), .ZN(n564) );
  NAND2_X1 U621 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U622 ( .A(n566), .B(KEYINPUT5), .ZN(n571) );
  NAND2_X1 U623 ( .A1(G63), .A2(n801), .ZN(n568) );
  NAND2_X1 U624 ( .A1(G51), .A2(n806), .ZN(n567) );
  NAND2_X1 U625 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U626 ( .A(KEYINPUT6), .B(n569), .Z(n570) );
  NAND2_X1 U627 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U628 ( .A(n572), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U629 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U630 ( .A1(G62), .A2(n801), .ZN(n574) );
  NAND2_X1 U631 ( .A1(G50), .A2(n806), .ZN(n573) );
  NAND2_X1 U632 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U633 ( .A(KEYINPUT81), .B(n575), .ZN(n579) );
  NAND2_X1 U634 ( .A1(G75), .A2(n802), .ZN(n577) );
  NAND2_X1 U635 ( .A1(G88), .A2(n805), .ZN(n576) );
  AND2_X1 U636 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U637 ( .A1(n579), .A2(n578), .ZN(G303) );
  INV_X1 U638 ( .A(G303), .ZN(G166) );
  NAND2_X1 U639 ( .A1(G49), .A2(n806), .ZN(n581) );
  NAND2_X1 U640 ( .A1(G74), .A2(G651), .ZN(n580) );
  NAND2_X1 U641 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U642 ( .A1(n801), .A2(n582), .ZN(n585) );
  NAND2_X1 U643 ( .A1(G87), .A2(n583), .ZN(n584) );
  NAND2_X1 U644 ( .A1(n585), .A2(n584), .ZN(G288) );
  NAND2_X1 U645 ( .A1(G61), .A2(n801), .ZN(n587) );
  NAND2_X1 U646 ( .A1(G86), .A2(n805), .ZN(n586) );
  NAND2_X1 U647 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U648 ( .A1(n802), .A2(G73), .ZN(n588) );
  XOR2_X1 U649 ( .A(KEYINPUT2), .B(n588), .Z(n589) );
  NOR2_X1 U650 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U651 ( .A1(n806), .A2(G48), .ZN(n591) );
  NAND2_X1 U652 ( .A1(n592), .A2(n591), .ZN(G305) );
  AND2_X1 U653 ( .A1(n801), .A2(G60), .ZN(n596) );
  NAND2_X1 U654 ( .A1(G72), .A2(n802), .ZN(n594) );
  NAND2_X1 U655 ( .A1(G85), .A2(n805), .ZN(n593) );
  NAND2_X1 U656 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U657 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U658 ( .A1(n806), .A2(G47), .ZN(n597) );
  NAND2_X1 U659 ( .A1(n598), .A2(n597), .ZN(G290) );
  XOR2_X1 U660 ( .A(KEYINPUT68), .B(KEYINPUT14), .Z(n600) );
  NAND2_X1 U661 ( .A1(G56), .A2(n801), .ZN(n599) );
  XNOR2_X1 U662 ( .A(n600), .B(n599), .ZN(n608) );
  NAND2_X1 U663 ( .A1(n802), .A2(G68), .ZN(n601) );
  XNOR2_X1 U664 ( .A(KEYINPUT69), .B(n601), .ZN(n604) );
  NAND2_X1 U665 ( .A1(n805), .A2(G81), .ZN(n602) );
  XOR2_X1 U666 ( .A(n602), .B(KEYINPUT12), .Z(n603) );
  NOR2_X1 U667 ( .A1(n604), .A2(n603), .ZN(n606) );
  NOR2_X1 U668 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U669 ( .A1(n806), .A2(G43), .ZN(n609) );
  NAND2_X1 U670 ( .A1(n610), .A2(n609), .ZN(n989) );
  XOR2_X1 U671 ( .A(G1996), .B(KEYINPUT96), .Z(n963) );
  INV_X1 U672 ( .A(KEYINPUT90), .ZN(n612) );
  NAND2_X1 U673 ( .A1(G40), .A2(G160), .ZN(n611) );
  XNOR2_X1 U674 ( .A(n611), .B(KEYINPUT84), .ZN(n720) );
  XNOR2_X1 U675 ( .A(n612), .B(n720), .ZN(n613) );
  NOR2_X1 U676 ( .A1(G164), .A2(G1384), .ZN(n719) );
  NAND2_X2 U677 ( .A1(n613), .A2(n719), .ZN(n675) );
  NOR2_X1 U678 ( .A1(n963), .A2(n675), .ZN(n614) );
  XNOR2_X1 U679 ( .A(n614), .B(KEYINPUT26), .ZN(n615) );
  NOR2_X1 U680 ( .A1(n989), .A2(n615), .ZN(n617) );
  NAND2_X1 U681 ( .A1(G1341), .A2(n675), .ZN(n616) );
  NAND2_X1 U682 ( .A1(n617), .A2(n616), .ZN(n633) );
  NAND2_X1 U683 ( .A1(n801), .A2(G66), .ZN(n618) );
  NAND2_X1 U684 ( .A1(n805), .A2(G92), .ZN(n619) );
  NAND2_X1 U685 ( .A1(n525), .A2(n619), .ZN(n621) );
  XNOR2_X1 U686 ( .A(n621), .B(n620), .ZN(n625) );
  NAND2_X1 U687 ( .A1(G79), .A2(n802), .ZN(n623) );
  NAND2_X1 U688 ( .A1(G54), .A2(n806), .ZN(n622) );
  NAND2_X1 U689 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U690 ( .A(KEYINPUT15), .B(n626), .ZN(n1003) );
  NOR2_X1 U691 ( .A1(n633), .A2(n1003), .ZN(n627) );
  XNOR2_X1 U692 ( .A(n627), .B(KEYINPUT97), .ZN(n632) );
  INV_X1 U693 ( .A(KEYINPUT95), .ZN(n628) );
  NAND2_X1 U694 ( .A1(G2067), .A2(n524), .ZN(n630) );
  NAND2_X1 U695 ( .A1(G1348), .A2(n675), .ZN(n629) );
  NAND2_X1 U696 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U697 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U698 ( .A1(n633), .A2(n1003), .ZN(n634) );
  NAND2_X1 U699 ( .A1(n635), .A2(n634), .ZN(n641) );
  INV_X1 U700 ( .A(G299), .ZN(n988) );
  NAND2_X1 U701 ( .A1(n524), .A2(G2072), .ZN(n637) );
  XNOR2_X1 U702 ( .A(n637), .B(KEYINPUT27), .ZN(n639) );
  INV_X1 U703 ( .A(G1956), .ZN(n1021) );
  NOR2_X1 U704 ( .A1(n1021), .A2(n524), .ZN(n638) );
  NOR2_X1 U705 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U706 ( .A1(n988), .A2(n642), .ZN(n640) );
  NAND2_X1 U707 ( .A1(n641), .A2(n640), .ZN(n645) );
  XOR2_X1 U708 ( .A(n643), .B(KEYINPUT28), .Z(n644) );
  NAND2_X1 U709 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U710 ( .A(n646), .B(KEYINPUT29), .ZN(n653) );
  INV_X1 U711 ( .A(n675), .ZN(n647) );
  NOR2_X1 U712 ( .A1(n647), .A2(G1961), .ZN(n648) );
  XNOR2_X1 U713 ( .A(n648), .B(KEYINPUT94), .ZN(n651) );
  INV_X1 U714 ( .A(n524), .ZN(n649) );
  XOR2_X1 U715 ( .A(G2078), .B(KEYINPUT25), .Z(n972) );
  NOR2_X1 U716 ( .A1(n649), .A2(n972), .ZN(n650) );
  NOR2_X1 U717 ( .A1(n651), .A2(n650), .ZN(n659) );
  NOR2_X1 U718 ( .A1(G301), .A2(n659), .ZN(n652) );
  NOR2_X1 U719 ( .A1(n653), .A2(n652), .ZN(n664) );
  NAND2_X1 U720 ( .A1(n675), .A2(G8), .ZN(n713) );
  NOR2_X1 U721 ( .A1(G1966), .A2(n713), .ZN(n654) );
  XOR2_X1 U722 ( .A(KEYINPUT93), .B(n654), .Z(n665) );
  NOR2_X1 U723 ( .A1(G2084), .A2(n675), .ZN(n655) );
  XOR2_X1 U724 ( .A(KEYINPUT92), .B(n655), .Z(n666) );
  NAND2_X1 U725 ( .A1(G8), .A2(n666), .ZN(n656) );
  NOR2_X1 U726 ( .A1(n665), .A2(n656), .ZN(n657) );
  XOR2_X1 U727 ( .A(KEYINPUT30), .B(n657), .Z(n658) );
  NOR2_X1 U728 ( .A1(G168), .A2(n658), .ZN(n661) );
  AND2_X1 U729 ( .A1(G301), .A2(n659), .ZN(n660) );
  NOR2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n662), .B(KEYINPUT31), .ZN(n663) );
  OR2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n674) );
  INV_X1 U733 ( .A(n674), .ZN(n671) );
  INV_X1 U734 ( .A(n665), .ZN(n669) );
  INV_X1 U735 ( .A(n666), .ZN(n667) );
  NAND2_X1 U736 ( .A1(G8), .A2(n667), .ZN(n668) );
  NAND2_X1 U737 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U738 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U739 ( .A(KEYINPUT98), .B(n672), .ZN(n687) );
  AND2_X1 U740 ( .A1(G286), .A2(G8), .ZN(n673) );
  NAND2_X1 U741 ( .A1(n674), .A2(n673), .ZN(n683) );
  INV_X1 U742 ( .A(G8), .ZN(n681) );
  NOR2_X1 U743 ( .A1(G2090), .A2(n675), .ZN(n676) );
  XNOR2_X1 U744 ( .A(KEYINPUT99), .B(n676), .ZN(n679) );
  NOR2_X1 U745 ( .A1(G1971), .A2(n713), .ZN(n677) );
  NOR2_X1 U746 ( .A1(G166), .A2(n677), .ZN(n678) );
  NAND2_X1 U747 ( .A1(n679), .A2(n678), .ZN(n680) );
  OR2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n682) );
  AND2_X1 U749 ( .A1(n683), .A2(n682), .ZN(n685) );
  INV_X1 U750 ( .A(KEYINPUT32), .ZN(n684) );
  XNOR2_X1 U751 ( .A(n685), .B(n684), .ZN(n686) );
  NOR2_X2 U752 ( .A1(n687), .A2(n686), .ZN(n709) );
  NOR2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n692) );
  NOR2_X1 U754 ( .A1(G1971), .A2(G303), .ZN(n688) );
  NOR2_X1 U755 ( .A1(n692), .A2(n688), .ZN(n997) );
  XOR2_X1 U756 ( .A(n997), .B(KEYINPUT100), .Z(n689) );
  NOR2_X1 U757 ( .A1(n709), .A2(n689), .ZN(n690) );
  NOR2_X1 U758 ( .A1(n690), .A2(n713), .ZN(n699) );
  NAND2_X1 U759 ( .A1(G1976), .A2(G288), .ZN(n996) );
  INV_X1 U760 ( .A(KEYINPUT33), .ZN(n701) );
  INV_X1 U761 ( .A(n713), .ZN(n691) );
  NAND2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U763 ( .A1(n701), .A2(n693), .ZN(n694) );
  XNOR2_X1 U764 ( .A(n694), .B(KEYINPUT101), .ZN(n700) );
  AND2_X1 U765 ( .A1(n996), .A2(n700), .ZN(n697) );
  OR2_X1 U766 ( .A1(G1981), .A2(G305), .ZN(n706) );
  NAND2_X1 U767 ( .A1(G1981), .A2(G305), .ZN(n695) );
  NAND2_X1 U768 ( .A1(n706), .A2(n695), .ZN(n986) );
  INV_X1 U769 ( .A(n986), .ZN(n696) );
  AND2_X1 U770 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U771 ( .A1(n699), .A2(n698), .ZN(n705) );
  INV_X1 U772 ( .A(n700), .ZN(n702) );
  OR2_X1 U773 ( .A1(n702), .A2(n701), .ZN(n703) );
  OR2_X1 U774 ( .A1(n986), .A2(n703), .ZN(n704) );
  NAND2_X1 U775 ( .A1(n705), .A2(n704), .ZN(n718) );
  XNOR2_X1 U776 ( .A(n706), .B(KEYINPUT24), .ZN(n707) );
  NOR2_X1 U777 ( .A1(n713), .A2(n707), .ZN(n708) );
  XNOR2_X1 U778 ( .A(n708), .B(KEYINPUT91), .ZN(n716) );
  INV_X1 U779 ( .A(n709), .ZN(n712) );
  NOR2_X1 U780 ( .A1(G2090), .A2(G303), .ZN(n710) );
  NAND2_X1 U781 ( .A1(G8), .A2(n710), .ZN(n711) );
  NAND2_X1 U782 ( .A1(n712), .A2(n711), .ZN(n714) );
  NAND2_X1 U783 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U784 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U785 ( .A1(n718), .A2(n717), .ZN(n750) );
  NOR2_X1 U786 ( .A1(n720), .A2(n719), .ZN(n765) );
  XNOR2_X1 U787 ( .A(KEYINPUT87), .B(KEYINPUT36), .ZN(n732) );
  NAND2_X1 U788 ( .A1(G104), .A2(n890), .ZN(n722) );
  NAND2_X1 U789 ( .A1(G140), .A2(n891), .ZN(n721) );
  NAND2_X1 U790 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U791 ( .A(n723), .B(KEYINPUT85), .ZN(n724) );
  XNOR2_X1 U792 ( .A(n724), .B(KEYINPUT34), .ZN(n730) );
  XNOR2_X1 U793 ( .A(KEYINPUT86), .B(KEYINPUT35), .ZN(n728) );
  NAND2_X1 U794 ( .A1(G116), .A2(n886), .ZN(n726) );
  NAND2_X1 U795 ( .A1(G128), .A2(n887), .ZN(n725) );
  NAND2_X1 U796 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U797 ( .A(n728), .B(n727), .ZN(n729) );
  NAND2_X1 U798 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U799 ( .A(n732), .B(n731), .ZN(n907) );
  XNOR2_X1 U800 ( .A(G2067), .B(KEYINPUT37), .ZN(n762) );
  NOR2_X1 U801 ( .A1(n907), .A2(n762), .ZN(n940) );
  NAND2_X1 U802 ( .A1(n765), .A2(n940), .ZN(n760) );
  NAND2_X1 U803 ( .A1(G105), .A2(n890), .ZN(n733) );
  XNOR2_X1 U804 ( .A(n733), .B(KEYINPUT38), .ZN(n740) );
  NAND2_X1 U805 ( .A1(G141), .A2(n891), .ZN(n735) );
  NAND2_X1 U806 ( .A1(G117), .A2(n886), .ZN(n734) );
  NAND2_X1 U807 ( .A1(n735), .A2(n734), .ZN(n738) );
  NAND2_X1 U808 ( .A1(n887), .A2(G129), .ZN(n736) );
  XOR2_X1 U809 ( .A(KEYINPUT88), .B(n736), .Z(n737) );
  NOR2_X1 U810 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U811 ( .A1(n740), .A2(n739), .ZN(n900) );
  NAND2_X1 U812 ( .A1(n900), .A2(G1996), .ZN(n741) );
  XNOR2_X1 U813 ( .A(n741), .B(KEYINPUT89), .ZN(n939) );
  NAND2_X1 U814 ( .A1(G131), .A2(n891), .ZN(n743) );
  NAND2_X1 U815 ( .A1(G119), .A2(n887), .ZN(n742) );
  NAND2_X1 U816 ( .A1(n743), .A2(n742), .ZN(n747) );
  NAND2_X1 U817 ( .A1(G95), .A2(n890), .ZN(n745) );
  NAND2_X1 U818 ( .A1(G107), .A2(n886), .ZN(n744) );
  NAND2_X1 U819 ( .A1(n745), .A2(n744), .ZN(n746) );
  OR2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n903) );
  AND2_X1 U821 ( .A1(n903), .A2(G1991), .ZN(n934) );
  OR2_X1 U822 ( .A1(n939), .A2(n934), .ZN(n748) );
  NAND2_X1 U823 ( .A1(n765), .A2(n748), .ZN(n754) );
  NAND2_X1 U824 ( .A1(n760), .A2(n754), .ZN(n749) );
  NOR2_X1 U825 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U826 ( .A(n751), .B(KEYINPUT102), .ZN(n753) );
  XNOR2_X1 U827 ( .A(G1986), .B(G290), .ZN(n995) );
  NAND2_X1 U828 ( .A1(n995), .A2(n765), .ZN(n752) );
  NAND2_X1 U829 ( .A1(n753), .A2(n752), .ZN(n768) );
  NOR2_X1 U830 ( .A1(G1996), .A2(n900), .ZN(n949) );
  INV_X1 U831 ( .A(n754), .ZN(n757) );
  NOR2_X1 U832 ( .A1(G1991), .A2(n903), .ZN(n933) );
  NOR2_X1 U833 ( .A1(G1986), .A2(G290), .ZN(n755) );
  NOR2_X1 U834 ( .A1(n933), .A2(n755), .ZN(n756) );
  NOR2_X1 U835 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U836 ( .A1(n949), .A2(n758), .ZN(n759) );
  XNOR2_X1 U837 ( .A(n759), .B(KEYINPUT39), .ZN(n761) );
  NAND2_X1 U838 ( .A1(n761), .A2(n760), .ZN(n763) );
  NAND2_X1 U839 ( .A1(n907), .A2(n762), .ZN(n954) );
  NAND2_X1 U840 ( .A1(n763), .A2(n954), .ZN(n764) );
  XOR2_X1 U841 ( .A(KEYINPUT103), .B(n764), .Z(n766) );
  NAND2_X1 U842 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U843 ( .A1(n768), .A2(n767), .ZN(n770) );
  XNOR2_X1 U844 ( .A(KEYINPUT40), .B(KEYINPUT104), .ZN(n769) );
  XNOR2_X1 U845 ( .A(n770), .B(n769), .ZN(G329) );
  AND2_X1 U846 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U847 ( .A(G57), .ZN(G237) );
  INV_X1 U848 ( .A(G132), .ZN(G219) );
  INV_X1 U849 ( .A(G82), .ZN(G220) );
  NAND2_X1 U850 ( .A1(G7), .A2(G661), .ZN(n771) );
  XNOR2_X1 U851 ( .A(n771), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U852 ( .A(G223), .ZN(n836) );
  NAND2_X1 U853 ( .A1(n836), .A2(G567), .ZN(n772) );
  XOR2_X1 U854 ( .A(KEYINPUT11), .B(n772), .Z(G234) );
  INV_X1 U855 ( .A(G860), .ZN(n778) );
  OR2_X1 U856 ( .A1(n989), .A2(n778), .ZN(G153) );
  INV_X1 U857 ( .A(G868), .ZN(n819) );
  NAND2_X1 U858 ( .A1(n1003), .A2(n819), .ZN(n773) );
  XNOR2_X1 U859 ( .A(n773), .B(KEYINPUT74), .ZN(n775) );
  NAND2_X1 U860 ( .A1(G868), .A2(G301), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n775), .A2(n774), .ZN(G284) );
  NAND2_X1 U862 ( .A1(G286), .A2(G868), .ZN(n777) );
  NAND2_X1 U863 ( .A1(G299), .A2(n819), .ZN(n776) );
  NAND2_X1 U864 ( .A1(n777), .A2(n776), .ZN(G297) );
  NAND2_X1 U865 ( .A1(n778), .A2(G559), .ZN(n779) );
  INV_X1 U866 ( .A(n1003), .ZN(n799) );
  NAND2_X1 U867 ( .A1(n779), .A2(n799), .ZN(n780) );
  XNOR2_X1 U868 ( .A(n780), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U869 ( .A1(n1003), .A2(n819), .ZN(n781) );
  XOR2_X1 U870 ( .A(KEYINPUT76), .B(n781), .Z(n782) );
  NOR2_X1 U871 ( .A1(G559), .A2(n782), .ZN(n785) );
  NOR2_X1 U872 ( .A1(G868), .A2(n989), .ZN(n783) );
  XOR2_X1 U873 ( .A(KEYINPUT75), .B(n783), .Z(n784) );
  NOR2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U875 ( .A(KEYINPUT77), .B(n786), .Z(G282) );
  NAND2_X1 U876 ( .A1(G123), .A2(n887), .ZN(n787) );
  XNOR2_X1 U877 ( .A(n787), .B(KEYINPUT78), .ZN(n788) );
  XNOR2_X1 U878 ( .A(n788), .B(KEYINPUT18), .ZN(n790) );
  NAND2_X1 U879 ( .A1(G135), .A2(n891), .ZN(n789) );
  NAND2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U881 ( .A(n791), .B(KEYINPUT79), .ZN(n793) );
  NAND2_X1 U882 ( .A1(G99), .A2(n890), .ZN(n792) );
  NAND2_X1 U883 ( .A1(n793), .A2(n792), .ZN(n796) );
  NAND2_X1 U884 ( .A1(n886), .A2(G111), .ZN(n794) );
  XOR2_X1 U885 ( .A(KEYINPUT80), .B(n794), .Z(n795) );
  NOR2_X1 U886 ( .A1(n796), .A2(n795), .ZN(n938) );
  XNOR2_X1 U887 ( .A(n938), .B(G2096), .ZN(n798) );
  INV_X1 U888 ( .A(G2100), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n798), .A2(n797), .ZN(G156) );
  NAND2_X1 U890 ( .A1(G559), .A2(n799), .ZN(n800) );
  XNOR2_X1 U891 ( .A(n800), .B(n989), .ZN(n817) );
  NOR2_X1 U892 ( .A1(n817), .A2(G860), .ZN(n811) );
  NAND2_X1 U893 ( .A1(G67), .A2(n801), .ZN(n804) );
  NAND2_X1 U894 ( .A1(G80), .A2(n802), .ZN(n803) );
  NAND2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n810) );
  NAND2_X1 U896 ( .A1(G93), .A2(n805), .ZN(n808) );
  NAND2_X1 U897 ( .A1(G55), .A2(n806), .ZN(n807) );
  NAND2_X1 U898 ( .A1(n808), .A2(n807), .ZN(n809) );
  OR2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n820) );
  XOR2_X1 U900 ( .A(n811), .B(n820), .Z(G145) );
  XNOR2_X1 U901 ( .A(KEYINPUT19), .B(G288), .ZN(n812) );
  XNOR2_X1 U902 ( .A(n812), .B(G305), .ZN(n813) );
  XOR2_X1 U903 ( .A(n820), .B(n813), .Z(n815) );
  XNOR2_X1 U904 ( .A(G290), .B(n988), .ZN(n814) );
  XNOR2_X1 U905 ( .A(n815), .B(n814), .ZN(n816) );
  XNOR2_X1 U906 ( .A(G166), .B(n816), .ZN(n911) );
  XNOR2_X1 U907 ( .A(n817), .B(n911), .ZN(n818) );
  NAND2_X1 U908 ( .A1(n818), .A2(G868), .ZN(n822) );
  NAND2_X1 U909 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U910 ( .A1(n822), .A2(n821), .ZN(G295) );
  NAND2_X1 U911 ( .A1(G2078), .A2(G2084), .ZN(n823) );
  XOR2_X1 U912 ( .A(KEYINPUT20), .B(n823), .Z(n824) );
  NAND2_X1 U913 ( .A1(G2090), .A2(n824), .ZN(n825) );
  XNOR2_X1 U914 ( .A(KEYINPUT21), .B(n825), .ZN(n826) );
  NAND2_X1 U915 ( .A1(n826), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U916 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U917 ( .A1(G220), .A2(G219), .ZN(n827) );
  XOR2_X1 U918 ( .A(KEYINPUT22), .B(n827), .Z(n828) );
  NOR2_X1 U919 ( .A1(G218), .A2(n828), .ZN(n829) );
  NAND2_X1 U920 ( .A1(G96), .A2(n829), .ZN(n840) );
  NAND2_X1 U921 ( .A1(n840), .A2(G2106), .ZN(n833) );
  NAND2_X1 U922 ( .A1(G69), .A2(G120), .ZN(n830) );
  NOR2_X1 U923 ( .A1(G237), .A2(n830), .ZN(n831) );
  NAND2_X1 U924 ( .A1(G108), .A2(n831), .ZN(n841) );
  NAND2_X1 U925 ( .A1(n841), .A2(G567), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(n842) );
  NAND2_X1 U927 ( .A1(G661), .A2(G483), .ZN(n834) );
  XNOR2_X1 U928 ( .A(KEYINPUT82), .B(n834), .ZN(n835) );
  NOR2_X1 U929 ( .A1(n842), .A2(n835), .ZN(n839) );
  NAND2_X1 U930 ( .A1(n839), .A2(G36), .ZN(G176) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n836), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U933 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U935 ( .A1(n839), .A2(n838), .ZN(G188) );
  XOR2_X1 U936 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  INV_X1 U938 ( .A(G120), .ZN(G236) );
  INV_X1 U939 ( .A(G69), .ZN(G235) );
  NOR2_X1 U940 ( .A1(n841), .A2(n840), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  INV_X1 U942 ( .A(n842), .ZN(G319) );
  XOR2_X1 U943 ( .A(KEYINPUT43), .B(KEYINPUT108), .Z(n844) );
  XNOR2_X1 U944 ( .A(KEYINPUT42), .B(G2678), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U946 ( .A(KEYINPUT107), .B(G2072), .Z(n846) );
  XNOR2_X1 U947 ( .A(G2067), .B(G2090), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U949 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U950 ( .A(G2096), .B(G2100), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n852) );
  XOR2_X1 U952 ( .A(G2078), .B(G2084), .Z(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(G227) );
  XOR2_X1 U954 ( .A(G1981), .B(G1966), .Z(n854) );
  XNOR2_X1 U955 ( .A(G1986), .B(G1971), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U957 ( .A(G1956), .B(G1976), .Z(n856) );
  XNOR2_X1 U958 ( .A(G1996), .B(G1991), .ZN(n855) );
  XNOR2_X1 U959 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U960 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U961 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(n862) );
  XOR2_X1 U963 ( .A(G1961), .B(G2474), .Z(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(G229) );
  XOR2_X1 U965 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n864) );
  NAND2_X1 U966 ( .A1(G124), .A2(n887), .ZN(n863) );
  XNOR2_X1 U967 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U968 ( .A(KEYINPUT110), .B(n865), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n891), .A2(G136), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U971 ( .A(KEYINPUT112), .B(n868), .Z(n870) );
  NAND2_X1 U972 ( .A1(n886), .A2(G112), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n873) );
  NAND2_X1 U974 ( .A1(G100), .A2(n890), .ZN(n871) );
  XNOR2_X1 U975 ( .A(KEYINPUT113), .B(n871), .ZN(n872) );
  NOR2_X1 U976 ( .A1(n873), .A2(n872), .ZN(G162) );
  NAND2_X1 U977 ( .A1(G115), .A2(n886), .ZN(n875) );
  NAND2_X1 U978 ( .A1(G127), .A2(n887), .ZN(n874) );
  NAND2_X1 U979 ( .A1(n875), .A2(n874), .ZN(n877) );
  XOR2_X1 U980 ( .A(KEYINPUT47), .B(KEYINPUT116), .Z(n876) );
  XNOR2_X1 U981 ( .A(n877), .B(n876), .ZN(n883) );
  NAND2_X1 U982 ( .A1(n891), .A2(G139), .ZN(n878) );
  XNOR2_X1 U983 ( .A(n878), .B(KEYINPUT114), .ZN(n880) );
  NAND2_X1 U984 ( .A1(G103), .A2(n890), .ZN(n879) );
  NAND2_X1 U985 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U986 ( .A(KEYINPUT115), .B(n881), .Z(n882) );
  NOR2_X1 U987 ( .A1(n883), .A2(n882), .ZN(n944) );
  XOR2_X1 U988 ( .A(KEYINPUT118), .B(KEYINPUT46), .Z(n885) );
  XNOR2_X1 U989 ( .A(KEYINPUT117), .B(KEYINPUT48), .ZN(n884) );
  XNOR2_X1 U990 ( .A(n885), .B(n884), .ZN(n898) );
  NAND2_X1 U991 ( .A1(G118), .A2(n886), .ZN(n889) );
  NAND2_X1 U992 ( .A1(G130), .A2(n887), .ZN(n888) );
  NAND2_X1 U993 ( .A1(n889), .A2(n888), .ZN(n896) );
  NAND2_X1 U994 ( .A1(G106), .A2(n890), .ZN(n893) );
  NAND2_X1 U995 ( .A1(G142), .A2(n891), .ZN(n892) );
  NAND2_X1 U996 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U997 ( .A(n894), .B(KEYINPUT45), .Z(n895) );
  NOR2_X1 U998 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U999 ( .A(n898), .B(n897), .Z(n902) );
  XOR2_X1 U1000 ( .A(G164), .B(n938), .Z(n899) );
  XNOR2_X1 U1001 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U1002 ( .A(n902), .B(n901), .Z(n905) );
  XOR2_X1 U1003 ( .A(G160), .B(n903), .Z(n904) );
  XNOR2_X1 U1004 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n944), .B(n906), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n907), .B(G162), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n910), .ZN(G395) );
  XNOR2_X1 U1009 ( .A(G171), .B(n989), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(n912), .B(n911), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n1003), .B(G286), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n915), .ZN(n916) );
  XOR2_X1 U1014 ( .A(KEYINPUT119), .B(n916), .Z(G397) );
  XOR2_X1 U1015 ( .A(G2454), .B(G2430), .Z(n918) );
  XNOR2_X1 U1016 ( .A(G2451), .B(G2446), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(n918), .B(n917), .ZN(n925) );
  XOR2_X1 U1018 ( .A(G2443), .B(G2427), .Z(n920) );
  XNOR2_X1 U1019 ( .A(G2438), .B(KEYINPUT105), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(n920), .B(n919), .ZN(n921) );
  XOR2_X1 U1021 ( .A(n921), .B(G2435), .Z(n923) );
  XNOR2_X1 U1022 ( .A(G1341), .B(G1348), .ZN(n922) );
  XNOR2_X1 U1023 ( .A(n923), .B(n922), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(n925), .B(n924), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n926), .A2(G14), .ZN(n932) );
  NAND2_X1 U1026 ( .A1(G319), .A2(n932), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(G227), .A2(G229), .ZN(n927) );
  XNOR2_X1 U1028 ( .A(KEYINPUT49), .B(n927), .ZN(n928) );
  NOR2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n931) );
  NOR2_X1 U1030 ( .A1(G395), .A2(G397), .ZN(n930) );
  NAND2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(G225) );
  INV_X1 U1032 ( .A(G225), .ZN(G308) );
  INV_X1 U1033 ( .A(G108), .ZN(G238) );
  INV_X1 U1034 ( .A(n932), .ZN(G401) );
  XNOR2_X1 U1035 ( .A(G160), .B(G2084), .ZN(n936) );
  NOR2_X1 U1036 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n942) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1041 ( .A(KEYINPUT120), .B(n943), .ZN(n957) );
  XOR2_X1 U1042 ( .A(G2072), .B(n944), .Z(n946) );
  XOR2_X1 U1043 ( .A(G164), .B(G2078), .Z(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1045 ( .A(KEYINPUT50), .B(n947), .Z(n953) );
  XOR2_X1 U1046 ( .A(G2090), .B(G162), .Z(n948) );
  NOR2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1048 ( .A(KEYINPUT121), .B(n950), .Z(n951) );
  XNOR2_X1 U1049 ( .A(KEYINPUT51), .B(n951), .ZN(n952) );
  NOR2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(KEYINPUT52), .B(n958), .ZN(n959) );
  INV_X1 U1054 ( .A(KEYINPUT55), .ZN(n981) );
  NAND2_X1 U1055 ( .A1(n959), .A2(n981), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n960), .A2(G29), .ZN(n1040) );
  XNOR2_X1 U1057 ( .A(KEYINPUT54), .B(KEYINPUT123), .ZN(n961) );
  XNOR2_X1 U1058 ( .A(n961), .B(G34), .ZN(n962) );
  XNOR2_X1 U1059 ( .A(G2084), .B(n962), .ZN(n979) );
  XNOR2_X1 U1060 ( .A(G2090), .B(G35), .ZN(n977) );
  XNOR2_X1 U1061 ( .A(n963), .B(G32), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(G1991), .B(G25), .ZN(n965) );
  XNOR2_X1 U1063 ( .A(G2072), .B(G33), .ZN(n964) );
  NOR2_X1 U1064 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1065 ( .A1(G28), .A2(n966), .ZN(n969) );
  XNOR2_X1 U1066 ( .A(KEYINPUT122), .B(G2067), .ZN(n967) );
  XNOR2_X1 U1067 ( .A(G26), .B(n967), .ZN(n968) );
  NOR2_X1 U1068 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1069 ( .A1(n971), .A2(n970), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(G27), .B(n972), .ZN(n973) );
  NOR2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1072 ( .A(KEYINPUT53), .B(n975), .ZN(n976) );
  NOR2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(n981), .B(n980), .ZN(n983) );
  INV_X1 U1076 ( .A(G29), .ZN(n982) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(G11), .A2(n984), .ZN(n1038) );
  XNOR2_X1 U1079 ( .A(G16), .B(KEYINPUT56), .ZN(n1009) );
  XOR2_X1 U1080 ( .A(G1966), .B(G168), .Z(n985) );
  NOR2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1082 ( .A(KEYINPUT57), .B(n987), .Z(n1007) );
  XNOR2_X1 U1083 ( .A(n988), .B(G1956), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(G301), .B(G1961), .ZN(n991) );
  XNOR2_X1 U1085 ( .A(n989), .B(G1341), .ZN(n990) );
  NOR2_X1 U1086 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n1002) );
  AND2_X1 U1089 ( .A1(G303), .A2(G1971), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1092 ( .A(n1000), .B(KEYINPUT124), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(G1348), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1036) );
  INV_X1 U1098 ( .A(G16), .ZN(n1034) );
  XNOR2_X1 U1099 ( .A(G1976), .B(G23), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(G1971), .B(G22), .ZN(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1102 ( .A(KEYINPUT126), .B(n1012), .Z(n1014) );
  XNOR2_X1 U1103 ( .A(G1986), .B(G24), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(KEYINPUT58), .B(n1015), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(G1961), .B(G5), .ZN(n1017) );
  XNOR2_X1 U1107 ( .A(G21), .B(G1966), .ZN(n1016) );
  NOR2_X1 U1108 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1109 ( .A1(n1019), .A2(n1018), .ZN(n1031) );
  XNOR2_X1 U1110 ( .A(KEYINPUT59), .B(G1348), .ZN(n1020) );
  XNOR2_X1 U1111 ( .A(n1020), .B(G4), .ZN(n1027) );
  XOR2_X1 U1112 ( .A(G1341), .B(G19), .Z(n1023) );
  XNOR2_X1 U1113 ( .A(n1021), .B(G20), .ZN(n1022) );
  NAND2_X1 U1114 ( .A1(n1023), .A2(n1022), .ZN(n1025) );
  XNOR2_X1 U1115 ( .A(G6), .B(G1981), .ZN(n1024) );
  NOR2_X1 U1116 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1117 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1118 ( .A(KEYINPUT125), .B(n1028), .Z(n1029) );
  XNOR2_X1 U1119 ( .A(KEYINPUT60), .B(n1029), .ZN(n1030) );
  NOR2_X1 U1120 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1121 ( .A(KEYINPUT61), .B(n1032), .ZN(n1033) );
  NAND2_X1 U1122 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1123 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NOR2_X1 U1124 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NAND2_X1 U1125 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XOR2_X1 U1126 ( .A(KEYINPUT62), .B(n1041), .Z(G311) );
  INV_X1 U1127 ( .A(G311), .ZN(G150) );
endmodule

