//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n580, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT66), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n454), .A2(G567), .ZN(new_n457));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n457), .B1(new_n451), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(KEYINPUT68), .A3(new_n463), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(G125), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n461), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n468), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n469), .A2(new_n463), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n461), .ZN(new_n477));
  INV_X1    g052(.A(G137), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT69), .ZN(G160));
  INV_X1    g056(.A(new_n477), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n476), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n483), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND3_X1  g065(.A1(new_n476), .A2(G126), .A3(G2105), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n461), .A2(G138), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n476), .A2(KEYINPUT4), .A3(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n466), .A2(new_n470), .A3(new_n492), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  XNOR2_X1  g076(.A(KEYINPUT6), .B(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G50), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n503), .A2(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(G62), .B1(new_n506), .B2(new_n505), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(KEYINPUT70), .B1(G75), .B2(G543), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT5), .B(G543), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(new_n515), .A3(G62), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n511), .B1(new_n517), .B2(G651), .ZN(G166));
  INV_X1    g093(.A(new_n505), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  OR2_X1    g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT71), .B(G89), .Z(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n528));
  INV_X1    g103(.A(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n529), .B1(new_n521), .B2(new_n522), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G51), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n525), .A2(new_n527), .A3(new_n528), .A4(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n514), .A2(G64), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(KEYINPUT72), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n503), .A2(new_n542), .B1(new_n509), .B2(new_n543), .ZN(new_n544));
  NOR3_X1   g119(.A1(new_n540), .A2(new_n541), .A3(new_n544), .ZN(G171));
  NAND3_X1  g120(.A1(new_n502), .A2(G43), .A3(G543), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n514), .A2(new_n502), .A3(G81), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  OAI211_X1 g123(.A(new_n546), .B(new_n547), .C1(new_n548), .C2(new_n534), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(new_n555));
  XOR2_X1   g130(.A(new_n555), .B(KEYINPUT73), .Z(G188));
  OAI211_X1 g131(.A(G53), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n557));
  AND2_X1   g132(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n558));
  NOR2_X1   g133(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n502), .A2(G53), .A3(G543), .A4(new_n558), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n514), .A2(new_n502), .A3(G91), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT76), .ZN(new_n565));
  XNOR2_X1  g140(.A(KEYINPUT75), .B(G65), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n514), .A2(new_n566), .B1(G78), .B2(G543), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n565), .B1(new_n567), .B2(new_n534), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(KEYINPUT75), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G65), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n506), .A2(new_n505), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n569), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n576), .A2(KEYINPUT76), .A3(G651), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n564), .B1(new_n568), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G299));
  NOR2_X1   g154(.A1(new_n541), .A2(new_n544), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n580), .B1(new_n539), .B2(new_n538), .ZN(G301));
  INV_X1    g156(.A(G166), .ZN(G303));
  NAND2_X1  g157(.A1(G74), .A2(G651), .ZN(new_n583));
  OAI211_X1 g158(.A(KEYINPUT77), .B(new_n583), .C1(new_n575), .C2(new_n534), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT77), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n585), .B(G651), .C1(new_n514), .C2(G74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n523), .A2(G87), .B1(new_n530), .B2(G49), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G288));
  AOI22_X1  g164(.A1(new_n514), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT78), .B1(new_n590), .B2(new_n534), .ZN(new_n591));
  OAI21_X1  g166(.A(G61), .B1(new_n506), .B2(new_n505), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n534), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n523), .A2(G86), .B1(new_n530), .B2(G48), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n591), .A2(new_n596), .A3(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n523), .A2(G85), .B1(new_n530), .B2(G47), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n534), .B2(new_n600), .ZN(G290));
  NAND3_X1  g176(.A1(new_n523), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n509), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n575), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(G54), .B2(new_n530), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G171), .B2(new_n612), .ZN(G284));
  OAI21_X1  g189(.A(new_n613), .B1(G171), .B2(new_n612), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(new_n578), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n616), .B1(new_n578), .B2(G868), .ZN(G280));
  INV_X1    g193(.A(new_n611), .ZN(new_n619));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G860), .ZN(G148));
  OR3_X1    g196(.A1(new_n611), .A2(KEYINPUT79), .A3(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(KEYINPUT79), .B1(new_n611), .B2(G559), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  MUX2_X1   g199(.A(new_n549), .B(new_n624), .S(G868), .Z(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g201(.A1(new_n466), .A2(new_n470), .A3(new_n474), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  INV_X1    g204(.A(G2100), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n485), .A2(G123), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n482), .A2(G135), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT80), .ZN(new_n635));
  OR3_X1    g210(.A1(new_n635), .A2(new_n461), .A3(G111), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n461), .B2(G111), .ZN(new_n637));
  OR2_X1    g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  NAND4_X1  g213(.A1(new_n636), .A2(G2104), .A3(new_n637), .A4(new_n638), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n633), .A2(new_n634), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  NAND3_X1  g216(.A1(new_n631), .A2(new_n632), .A3(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT82), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2430), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(KEYINPUT14), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G1341), .B(G1348), .Z(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(G14), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n653), .ZN(G401));
  XOR2_X1   g233(.A(KEYINPUT83), .B(KEYINPUT18), .Z(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g237(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n659), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n662), .B2(new_n659), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n665), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2096), .B(G2100), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XOR2_X1   g245(.A(G1991), .B(G1996), .Z(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT19), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  AND2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT85), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n675), .A2(new_n676), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n674), .A2(new_n677), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n674), .B2(new_n683), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n681), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n686), .A2(new_n688), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n671), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n691), .ZN(new_n693));
  INV_X1    g268(.A(new_n671), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n693), .A2(new_n694), .A3(new_n689), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  AND3_X1   g271(.A1(new_n692), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n696), .B1(new_n692), .B2(new_n695), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(G229));
  INV_X1    g274(.A(G11), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n700), .A2(KEYINPUT31), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(KEYINPUT31), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT30), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n703), .A2(G28), .ZN(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n703), .B2(G28), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n701), .B(new_n702), .C1(new_n704), .C2(new_n706), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n640), .A2(new_n705), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT97), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n709), .B2(new_n708), .ZN(new_n711));
  INV_X1    g286(.A(G2078), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n705), .A2(G27), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT98), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n500), .B2(G29), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n711), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n717), .A2(G21), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G286), .B2(G16), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT95), .B(G1966), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n717), .A2(G19), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n550), .B2(new_n717), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(G1341), .Z(new_n724));
  AND3_X1   g299(.A1(new_n716), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n705), .A2(G26), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT28), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n482), .A2(G140), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n485), .A2(G128), .ZN(new_n729));
  OR2_X1    g304(.A1(G104), .A2(G2105), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n730), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n728), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n727), .B1(new_n733), .B2(new_n705), .ZN(new_n734));
  INV_X1    g309(.A(G2067), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G1348), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n619), .A2(G16), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G4), .B2(G16), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n736), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n715), .A2(new_n712), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n739), .A2(new_n737), .ZN(new_n742));
  NOR3_X1   g317(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n705), .A2(G35), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n489), .B2(G29), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT29), .ZN(new_n746));
  INV_X1    g321(.A(G2090), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT99), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n725), .A2(new_n743), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n482), .A2(G141), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT92), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n474), .A2(G105), .ZN(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT26), .ZN(new_n756));
  AOI211_X1 g331(.A(new_n754), .B(new_n756), .C1(new_n485), .C2(G129), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  OR3_X1    g333(.A1(new_n758), .A2(KEYINPUT93), .A3(new_n705), .ZN(new_n759));
  OR2_X1    g334(.A1(G29), .A2(G32), .ZN(new_n760));
  OAI211_X1 g335(.A(KEYINPUT93), .B(new_n760), .C1(new_n758), .C2(new_n705), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT27), .B(G1996), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT94), .Z(new_n764));
  OR2_X1    g339(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n717), .A2(G5), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G171), .B2(new_n717), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(G1961), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n762), .B2(new_n764), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n705), .A2(G33), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT25), .Z(new_n772));
  INV_X1    g347(.A(G139), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n477), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n466), .A2(G127), .A3(new_n470), .ZN(new_n775));
  NAND2_X1  g350(.A1(G115), .A2(G2104), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n461), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n770), .B1(new_n778), .B2(new_n705), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n779), .A2(G2072), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G1961), .B2(new_n767), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n719), .A2(new_n720), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT96), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G2072), .B2(new_n779), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n765), .A2(new_n769), .A3(new_n781), .A4(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(G34), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n786), .A2(KEYINPUT24), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(KEYINPUT24), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n705), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G160), .B2(new_n705), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2084), .ZN(new_n791));
  OR3_X1    g366(.A1(new_n750), .A2(new_n785), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n746), .A2(new_n747), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT100), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n717), .A2(G20), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT23), .Z(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G299), .B2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1956), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT101), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n794), .A2(KEYINPUT101), .A3(new_n798), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n792), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n705), .A2(G25), .ZN(new_n805));
  NOR2_X1   g380(.A1(G95), .A2(G2105), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT86), .Z(new_n807));
  OAI21_X1  g382(.A(G2104), .B1(new_n461), .B2(G107), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(G119), .ZN(new_n810));
  INV_X1    g385(.A(G131), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n810), .A2(new_n484), .B1(new_n477), .B2(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n805), .B1(new_n814), .B2(new_n705), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT35), .B(G1991), .Z(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n815), .B(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(KEYINPUT91), .B2(KEYINPUT36), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n717), .A2(G24), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n600), .A2(new_n534), .ZN(new_n821));
  INV_X1    g396(.A(G47), .ZN(new_n822));
  INV_X1    g397(.A(G85), .ZN(new_n823));
  OAI22_X1  g398(.A1(new_n503), .A2(new_n822), .B1(new_n509), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n820), .B1(new_n825), .B2(new_n717), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT87), .B(G1986), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n819), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n587), .A2(new_n588), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(new_n717), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n717), .B2(G23), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT88), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT33), .B(G1976), .Z(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  MUX2_X1   g413(.A(G6), .B(G305), .S(G16), .Z(new_n839));
  XOR2_X1   g414(.A(KEYINPUT32), .B(G1981), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(G166), .A2(G16), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(G16), .B2(G22), .ZN(new_n844));
  XNOR2_X1  g419(.A(KEYINPUT89), .B(G1971), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT90), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n844), .B(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n835), .B2(new_n837), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n842), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT34), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n830), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(KEYINPUT34), .B1(new_n842), .B2(new_n848), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n848), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n856), .A2(new_n850), .A3(new_n838), .A4(new_n841), .ZN(new_n857));
  INV_X1    g432(.A(new_n854), .ZN(new_n858));
  INV_X1    g433(.A(new_n830), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n857), .A2(new_n852), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n804), .A2(new_n855), .A3(KEYINPUT102), .A4(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n750), .A2(new_n785), .A3(new_n791), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n863), .A2(new_n860), .A3(new_n801), .A4(new_n802), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n858), .B1(new_n851), .B2(new_n852), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n861), .A2(new_n866), .ZN(G311));
  NAND3_X1  g442(.A1(new_n804), .A2(new_n855), .A3(new_n860), .ZN(G150));
  NOR2_X1   g443(.A1(new_n611), .A2(new_n620), .ZN(new_n869));
  XNOR2_X1  g444(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n547), .A2(new_n546), .ZN(new_n872));
  AOI22_X1  g447(.A1(new_n523), .A2(G93), .B1(new_n530), .B2(G55), .ZN(new_n873));
  NAND2_X1  g448(.A1(G68), .A2(G543), .ZN(new_n874));
  INV_X1    g449(.A(G56), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n874), .B1(new_n575), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(G651), .ZN(new_n877));
  OAI21_X1  g452(.A(G67), .B1(new_n506), .B2(new_n505), .ZN(new_n878));
  NAND2_X1  g453(.A1(G80), .A2(G543), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n534), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n872), .A2(new_n873), .A3(new_n877), .A4(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n502), .A2(G55), .A3(G543), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n514), .A2(new_n502), .A3(G93), .ZN(new_n884));
  INV_X1    g459(.A(new_n879), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(new_n514), .B2(G67), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n883), .B(new_n884), .C1(new_n886), .C2(new_n534), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n549), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n882), .A2(new_n888), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n871), .B(new_n889), .Z(new_n890));
  AND2_X1   g465(.A1(new_n890), .A2(KEYINPUT39), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(KEYINPUT39), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n891), .A2(new_n892), .A3(G860), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n887), .A2(G860), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT37), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n893), .A2(new_n895), .ZN(G145));
  AND2_X1   g471(.A1(new_n753), .A2(new_n757), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n897), .A2(new_n778), .ZN(new_n898));
  NOR3_X1   g473(.A1(new_n758), .A2(new_n777), .A3(new_n774), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n482), .A2(G142), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n485), .A2(G130), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n461), .A2(G118), .ZN(new_n902));
  OAI21_X1  g477(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n900), .B(new_n901), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n628), .ZN(new_n905));
  OR3_X1    g480(.A1(new_n898), .A2(new_n899), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n905), .B1(new_n898), .B2(new_n899), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n500), .B(new_n732), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(new_n813), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(G160), .B(new_n640), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(G162), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n906), .A2(new_n910), .A3(new_n907), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n912), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G37), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n914), .B1(new_n912), .B2(new_n915), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n920), .B(new_n921), .ZN(G395));
  XNOR2_X1  g497(.A(new_n624), .B(new_n889), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n578), .A2(new_n611), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT41), .B1(new_n578), .B2(new_n611), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(KEYINPUT105), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n578), .A2(new_n929), .A3(new_n611), .ZN(new_n930));
  NAND2_X1  g505(.A1(G299), .A2(new_n619), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT41), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n927), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OR3_X1    g509(.A1(new_n923), .A2(new_n934), .A3(KEYINPUT106), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n931), .A2(new_n924), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n923), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT106), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n923), .A2(new_n934), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OR2_X1    g515(.A1(new_n940), .A2(KEYINPUT42), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n942));
  XNOR2_X1  g517(.A(G166), .B(G305), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n825), .B(G288), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n502), .A2(G48), .A3(G543), .ZN(new_n946));
  INV_X1    g521(.A(G86), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n946), .B1(new_n947), .B2(new_n509), .ZN(new_n948));
  INV_X1    g523(.A(new_n594), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n948), .B1(KEYINPUT78), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(G166), .A2(new_n950), .A3(new_n596), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n534), .B1(new_n513), .B2(new_n516), .ZN(new_n952));
  OAI21_X1  g527(.A(G305), .B1(new_n952), .B2(new_n511), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n831), .A2(new_n825), .ZN(new_n955));
  NAND2_X1  g530(.A1(G290), .A2(G288), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(KEYINPUT107), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT108), .B1(new_n954), .B2(new_n957), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n944), .A2(new_n960), .A3(new_n953), .A4(new_n951), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n945), .A2(new_n958), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n940), .A2(KEYINPUT42), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n941), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n962), .B1(new_n941), .B2(new_n963), .ZN(new_n965));
  OAI21_X1  g540(.A(G868), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n887), .A2(new_n612), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(G295));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n967), .ZN(G331));
  AND3_X1   g544(.A1(new_n882), .A2(new_n888), .A3(G286), .ZN(new_n970));
  AOI21_X1  g545(.A(G286), .B1(new_n882), .B2(new_n888), .ZN(new_n971));
  OAI21_X1  g546(.A(G301), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AOI22_X1  g547(.A1(new_n877), .A2(new_n872), .B1(new_n873), .B2(new_n881), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n549), .A2(new_n887), .ZN(new_n974));
  OAI21_X1  g549(.A(G168), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n882), .A2(new_n888), .A3(G286), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n975), .A2(G171), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n936), .B1(new_n972), .B2(new_n977), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n972), .A2(new_n977), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n978), .B1(new_n934), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n917), .B1(new_n980), .B2(new_n962), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n934), .A2(new_n979), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n972), .A2(new_n977), .ZN(new_n983));
  INV_X1    g558(.A(new_n936), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n982), .A2(new_n962), .A3(new_n985), .ZN(new_n986));
  OR3_X1    g561(.A1(new_n981), .A2(new_n986), .A3(KEYINPUT43), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n988));
  INV_X1    g563(.A(new_n927), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n578), .A2(new_n929), .A3(new_n611), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n929), .B1(new_n578), .B2(new_n611), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n578), .A2(new_n611), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n989), .B1(new_n993), .B2(KEYINPUT41), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n985), .B1(new_n994), .B2(new_n983), .ZN(new_n995));
  INV_X1    g570(.A(new_n962), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n984), .B1(new_n983), .B2(new_n933), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n932), .A2(new_n972), .A3(KEYINPUT41), .A4(new_n977), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n962), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n997), .A2(new_n917), .A3(new_n1000), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n987), .B(KEYINPUT44), .C1(new_n988), .C2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT43), .B1(new_n981), .B2(new_n986), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n997), .A2(new_n988), .A3(new_n917), .A4(new_n1000), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT109), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n1008));
  AOI211_X1 g583(.A(new_n1008), .B(KEYINPUT44), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1002), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT110), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1002), .B(new_n1012), .C1(new_n1007), .C2(new_n1009), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(G397));
  NOR2_X1   g589(.A1(G305), .A2(G1981), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n949), .B1(new_n597), .B2(KEYINPUT115), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n948), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(G1981), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT49), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT116), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1024));
  NOR3_X1   g599(.A1(G305), .A2(KEYINPUT114), .A3(G1981), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1021), .B(new_n1023), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G40), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n473), .A2(new_n479), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1384), .B1(new_n496), .B2(new_n499), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(G8), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1023), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OR2_X1    g608(.A1(G288), .A2(G1976), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1017), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1030), .A2(G8), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1036), .B(KEYINPUT117), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n831), .A2(G1976), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1030), .A2(G8), .A3(new_n1039), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1040), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT113), .B1(new_n1040), .B2(KEYINPUT52), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1043), .B1(new_n831), .B2(G1976), .ZN(new_n1044));
  OAI22_X1  g619(.A1(new_n1041), .A2(new_n1042), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1033), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  NOR2_X1   g622(.A1(G166), .A2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1048), .B(KEYINPUT55), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1029), .A2(KEYINPUT45), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1050), .A2(new_n1028), .ZN(new_n1051));
  INV_X1    g626(.A(G1384), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n500), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT45), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(G1971), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1029), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1028), .B1(new_n1029), .B2(new_n1057), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1059), .A2(new_n1060), .A3(G2090), .ZN(new_n1061));
  OAI211_X1 g636(.A(G8), .B(new_n1049), .C1(new_n1056), .C2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT112), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1050), .A2(new_n1028), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1029), .A2(KEYINPUT45), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1053), .A2(KEYINPUT50), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(new_n1028), .A3(new_n1058), .ZN(new_n1068));
  OAI22_X1  g643(.A1(new_n1066), .A2(G1971), .B1(new_n1068), .B2(G2090), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT112), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1069), .A2(new_n1070), .A3(G8), .A4(new_n1049), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1046), .A2(new_n1063), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1038), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1049), .B1(new_n1069), .B2(G8), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1074), .B1(new_n1063), .B2(new_n1071), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1050), .A2(KEYINPUT118), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1029), .A2(new_n1077), .A3(KEYINPUT45), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1076), .A2(new_n1078), .A3(new_n1028), .A4(new_n1055), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1080));
  INV_X1    g655(.A(G2084), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1079), .A2(new_n720), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1082), .A2(new_n1047), .A3(G286), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1075), .A2(new_n1046), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT63), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1075), .A2(KEYINPUT63), .A3(new_n1046), .A4(new_n1083), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1073), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1055), .A2(new_n712), .A3(new_n1050), .A4(new_n1028), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G1961), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1068), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1090), .A2(G2078), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1091), .B(new_n1093), .C1(new_n1095), .C2(new_n1079), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(G171), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n1098));
  NOR2_X1   g673(.A1(G168), .A2(new_n1047), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1079), .A2(new_n720), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g680(.A(G8), .B(new_n1102), .C1(new_n1105), .C2(G286), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1099), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1107), .B(new_n1101), .C1(new_n1082), .C2(new_n1047), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1105), .A2(new_n1099), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1106), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1097), .B1(new_n1110), .B2(KEYINPUT62), .ZN(new_n1111));
  INV_X1    g686(.A(G1956), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1068), .A2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n578), .B(KEYINPUT57), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT56), .B(G2072), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(KEYINPUT119), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1055), .A2(new_n1050), .A3(new_n1028), .A4(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1113), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1030), .A2(G2067), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n1068), .B2(new_n737), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1120), .A2(new_n611), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1114), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1118), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT120), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1125), .B(new_n1118), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n611), .B1(new_n1120), .B2(KEYINPUT60), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(KEYINPUT60), .B2(new_n1120), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1113), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1129), .B1(new_n1130), .B2(new_n1122), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1114), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(KEYINPUT61), .A3(new_n1118), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1128), .A2(new_n1131), .A3(new_n1135), .ZN(new_n1136));
  XOR2_X1   g711(.A(KEYINPUT58), .B(G1341), .Z(new_n1137));
  NAND2_X1  g712(.A1(new_n1030), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT121), .B(G1996), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n550), .ZN(new_n1142));
  NAND2_X1  g717(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1141), .A2(KEYINPUT122), .A3(KEYINPUT59), .A4(new_n550), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1120), .A2(KEYINPUT60), .A3(new_n611), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1124), .B(new_n1126), .C1(new_n1136), .C2(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1029), .A2(KEYINPUT111), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1054), .B1(new_n1029), .B2(KEYINPUT111), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1051), .B(new_n1094), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1151), .A2(new_n1091), .A3(G301), .A4(new_n1093), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT54), .B1(new_n1097), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT54), .B1(new_n1096), .B2(G171), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1151), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1155), .B1(new_n1156), .B2(G171), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1156), .A2(new_n1155), .A3(G171), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1153), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1111), .B1(new_n1148), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1096), .A2(KEYINPUT62), .A3(G171), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1106), .A2(new_n1108), .A3(new_n1162), .A4(new_n1109), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1075), .A2(new_n1164), .A3(new_n1046), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n1075), .B2(new_n1046), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1163), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1088), .B1(new_n1161), .B2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1028), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n897), .B(G1996), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n732), .B(new_n735), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n814), .A2(new_n816), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n813), .A2(new_n817), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(G290), .B(G1986), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1171), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1168), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n897), .A2(new_n1173), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1171), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1170), .A2(G1996), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1182), .A2(KEYINPUT126), .A3(KEYINPUT46), .ZN(new_n1183));
  AOI21_X1  g758(.A(KEYINPUT126), .B1(new_n1182), .B2(KEYINPUT46), .ZN(new_n1184));
  OAI221_X1 g759(.A(new_n1181), .B1(KEYINPUT46), .B2(new_n1182), .C1(new_n1183), .C2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT47), .ZN(new_n1186));
  OR3_X1    g761(.A1(new_n1170), .A2(G1986), .A3(G290), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1187), .ZN(new_n1188));
  OR2_X1    g763(.A1(new_n1188), .A2(KEYINPUT48), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1176), .A2(new_n1171), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1188), .A2(KEYINPUT48), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1193));
  OAI22_X1  g768(.A1(new_n1193), .A2(new_n1174), .B1(G2067), .B2(new_n732), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(new_n1171), .ZN(new_n1195));
  AND3_X1   g770(.A1(new_n1186), .A2(new_n1192), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1179), .A2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g772(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1199));
  OAI21_X1  g773(.A(new_n1199), .B1(new_n697), .B2(new_n698), .ZN(new_n1200));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n1201));
  NAND2_X1  g775(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  OAI211_X1 g776(.A(KEYINPUT127), .B(new_n1199), .C1(new_n697), .C2(new_n698), .ZN(new_n1203));
  AOI21_X1  g777(.A(new_n920), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g778(.A1(new_n1204), .A2(new_n1005), .ZN(G225));
  INV_X1    g779(.A(G225), .ZN(G308));
endmodule


