//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n192), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT77), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n192), .A2(new_n194), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n199), .B1(G143), .B2(new_n191), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n198), .B1(new_n200), .B2(new_n189), .ZN(new_n201));
  XNOR2_X1  g015(.A(G143), .B(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT77), .A3(new_n190), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n197), .A2(new_n201), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(new_n205), .B2(G107), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G104), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(G107), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n206), .A2(new_n209), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n205), .A2(G107), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n208), .A2(G104), .ZN(new_n214));
  OAI21_X1  g028(.A(G101), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n204), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT10), .ZN(new_n218));
  AND2_X1   g032(.A1(KEYINPUT66), .A2(G128), .ZN(new_n219));
  NOR2_X1   g033(.A1(KEYINPUT66), .A2(G128), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n198), .B1(new_n221), .B2(new_n200), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n218), .B1(new_n222), .B2(new_n195), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n217), .A2(new_n218), .B1(new_n216), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n206), .A2(new_n209), .A3(new_n211), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT76), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT76), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n206), .A2(new_n209), .A3(new_n227), .A4(new_n211), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(G101), .A3(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n212), .A2(KEYINPUT4), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  XOR2_X1   g045(.A(KEYINPUT0), .B(G128), .Z(new_n232));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(new_n233), .A3(new_n198), .ZN(new_n234));
  OAI211_X1 g048(.A(KEYINPUT0), .B(G128), .C1(new_n202), .C2(KEYINPUT64), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n226), .A2(new_n237), .A3(G101), .A4(new_n228), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n231), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT11), .ZN(new_n240));
  INV_X1    g054(.A(G134), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(G137), .ZN(new_n242));
  INV_X1    g056(.A(G137), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(KEYINPUT11), .A3(G134), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(G137), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G131), .ZN(new_n247));
  INV_X1    g061(.A(G131), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n242), .A2(new_n244), .A3(new_n248), .A4(new_n245), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n247), .A2(KEYINPUT68), .A3(new_n249), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n224), .A2(new_n239), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT78), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n224), .A2(new_n239), .A3(KEYINPUT78), .A4(new_n254), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT69), .B(G953), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G227), .ZN(new_n261));
  XOR2_X1   g075(.A(G110), .B(G140), .Z(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n212), .A2(new_n215), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n222), .A3(new_n195), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n217), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT79), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n254), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n217), .A2(new_n266), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(KEYINPUT79), .B2(KEYINPUT12), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n250), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n269), .A2(new_n271), .B1(KEYINPUT12), .B2(new_n272), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n259), .A2(new_n264), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n224), .A2(new_n239), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n253), .A3(new_n252), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n264), .B1(new_n259), .B2(new_n276), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n187), .B(new_n188), .C1(new_n274), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n259), .A2(new_n273), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n263), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n263), .B1(new_n257), .B2(new_n258), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n276), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n280), .A2(G469), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(G469), .A2(G902), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n278), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT9), .B(G234), .ZN(new_n286));
  OAI21_X1  g100(.A(G221), .B1(new_n286), .B2(G902), .ZN(new_n287));
  OAI21_X1  g101(.A(G214), .B1(G237), .B2(G902), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(G116), .B(G119), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT2), .B(G113), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n290), .B(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n231), .A2(new_n293), .A3(new_n238), .ZN(new_n294));
  INV_X1    g108(.A(G119), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G116), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT80), .B1(new_n296), .B2(KEYINPUT5), .ZN(new_n297));
  INV_X1    g111(.A(G116), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G119), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n296), .A2(new_n299), .A3(KEYINPUT5), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT80), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT5), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n301), .A2(new_n302), .A3(new_n295), .A4(G116), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n297), .A2(new_n300), .A3(G113), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n296), .A2(new_n299), .ZN(new_n305));
  OR2_X1    g119(.A1(new_n305), .A2(new_n291), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(new_n265), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n294), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(G110), .B(G122), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n292), .B1(new_n229), .B2(new_n230), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n308), .B1(new_n314), .B2(new_n238), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n311), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n313), .A2(KEYINPUT6), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G125), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT72), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G125), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n234), .A2(new_n235), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n322), .B1(new_n222), .B2(new_n195), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G224), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n326), .A2(G953), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n325), .B(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT6), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n310), .A2(new_n329), .A3(new_n312), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n317), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n327), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n325), .A2(KEYINPUT7), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(KEYINPUT7), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n334), .B1(new_n323), .B2(new_n324), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n307), .B(new_n265), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n311), .B(KEYINPUT8), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n333), .A2(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(G902), .B1(new_n338), .B2(new_n316), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n331), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(G210), .B1(G237), .B2(G902), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n331), .A2(new_n341), .A3(new_n339), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n289), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n285), .A2(new_n287), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT95), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT16), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n320), .A2(G125), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n318), .A2(KEYINPUT72), .ZN(new_n350));
  OAI21_X1  g164(.A(G140), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(G125), .A2(G140), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n348), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G140), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n322), .A2(new_n348), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n191), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G953), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT69), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT69), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G953), .ZN(new_n362));
  INV_X1    g176(.A(G237), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n360), .A2(new_n362), .A3(G214), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n193), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n260), .A2(G143), .A3(G214), .A4(new_n363), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(KEYINPUT17), .A3(G131), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n352), .B1(new_n322), .B2(G140), .ZN(new_n369));
  OAI211_X1 g183(.A(G146), .B(new_n356), .C1(new_n369), .C2(new_n348), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n358), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT85), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT81), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n374), .B1(new_n367), .B2(G131), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT17), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n365), .A2(new_n366), .A3(KEYINPUT81), .A4(new_n248), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n367), .A2(G131), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n375), .A2(new_n376), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n358), .A2(new_n368), .A3(KEYINPUT85), .A4(new_n370), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n373), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(G113), .B(G122), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT84), .B(G104), .ZN(new_n383));
  XOR2_X1   g197(.A(new_n382), .B(new_n383), .Z(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n367), .A2(KEYINPUT18), .A3(G131), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n369), .A2(G146), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n318), .A2(new_n355), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n191), .B1(new_n388), .B2(new_n352), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(KEYINPUT18), .A2(G131), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n365), .A2(new_n366), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n386), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n381), .A2(new_n385), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT86), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n381), .A2(KEYINPUT86), .A3(new_n385), .A4(new_n393), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n375), .A2(new_n377), .A3(new_n378), .ZN(new_n399));
  XOR2_X1   g213(.A(KEYINPUT83), .B(KEYINPUT19), .Z(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(new_n352), .B2(new_n388), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n369), .A2(KEYINPUT19), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n402), .A2(KEYINPUT82), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(KEYINPUT82), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n401), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n370), .B(new_n399), .C1(new_n405), .C2(G146), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n385), .B1(new_n406), .B2(new_n393), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n398), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT20), .ZN(new_n410));
  NOR2_X1   g224(.A1(G475), .A2(G902), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT87), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n409), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n407), .B1(new_n396), .B2(new_n397), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT20), .B1(new_n415), .B2(new_n412), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n381), .A2(new_n393), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n384), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n398), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n188), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n414), .A2(new_n416), .B1(new_n420), .B2(G475), .ZN(new_n421));
  INV_X1    g235(.A(G217), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n286), .A2(new_n422), .A3(G953), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  OR2_X1    g238(.A1(KEYINPUT66), .A2(G128), .ZN(new_n425));
  NAND2_X1  g239(.A1(KEYINPUT66), .A2(G128), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(G143), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n193), .A2(G128), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n241), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n298), .A2(G122), .ZN(new_n430));
  INV_X1    g244(.A(G122), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G116), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n430), .A2(new_n432), .A3(new_n208), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n431), .A2(G116), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n298), .A2(G122), .ZN(new_n435));
  OAI21_X1  g249(.A(G107), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n429), .A2(KEYINPUT90), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT90), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n427), .A2(new_n438), .A3(new_n241), .A4(new_n428), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n428), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT13), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n442), .A2(KEYINPUT88), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(KEYINPUT88), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n441), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT88), .B(KEYINPUT13), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n428), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(new_n447), .A3(new_n427), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G134), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT89), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n448), .A2(KEYINPUT89), .A3(G134), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n440), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n433), .ZN(new_n454));
  OR3_X1    g268(.A1(new_n430), .A2(KEYINPUT91), .A3(KEYINPUT14), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n435), .B1(KEYINPUT14), .B2(new_n430), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT91), .B1(new_n430), .B2(KEYINPUT14), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n454), .B1(new_n458), .B2(G107), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n427), .A2(new_n428), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G134), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n429), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n453), .A2(new_n464), .A3(KEYINPUT92), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT92), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n448), .A2(KEYINPUT89), .A3(G134), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT89), .B1(new_n448), .B2(G134), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n439), .B(new_n437), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n466), .B1(new_n469), .B2(new_n463), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n424), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT92), .B1(new_n453), .B2(new_n464), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n469), .A2(new_n466), .A3(new_n463), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n423), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n471), .A2(new_n188), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G478), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(KEYINPUT15), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G952), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n479), .A2(KEYINPUT93), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n479), .A2(KEYINPUT93), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n359), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(G234), .B2(G237), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n260), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n188), .B1(G234), .B2(G237), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  XOR2_X1   g301(.A(new_n487), .B(KEYINPUT94), .Z(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT21), .B(G898), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n484), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n477), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n471), .A2(new_n188), .A3(new_n474), .A4(new_n492), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n478), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n346), .A2(new_n347), .A3(new_n421), .A4(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n260), .A2(G221), .A3(G234), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT22), .B(G137), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n496), .B(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT24), .B(G110), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n219), .A2(new_n220), .A3(new_n295), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n189), .A2(G119), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT23), .B1(new_n189), .B2(G119), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(new_n502), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n425), .A2(KEYINPUT23), .A3(G119), .A4(new_n426), .ZN(new_n506));
  INV_X1    g320(.A(G110), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n503), .A2(new_n508), .A3(KEYINPUT73), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n370), .A3(new_n389), .ZN(new_n510));
  AOI21_X1  g324(.A(KEYINPUT73), .B1(new_n503), .B2(new_n508), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n501), .A2(new_n502), .ZN(new_n513));
  INV_X1    g327(.A(new_n500), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n505), .A2(new_n506), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G110), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n518), .B1(new_n358), .B2(new_n370), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n499), .B1(new_n512), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n358), .A2(new_n370), .ZN(new_n521));
  INV_X1    g335(.A(new_n518), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n503), .A2(new_n508), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT73), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n526), .A2(new_n370), .A3(new_n509), .A4(new_n389), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n523), .A2(new_n527), .A3(new_n498), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n520), .A2(new_n188), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT25), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n520), .A2(KEYINPUT25), .A3(new_n528), .A4(new_n188), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(KEYINPUT74), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n422), .B1(G234), .B2(new_n188), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT74), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n529), .A2(new_n535), .A3(new_n530), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT75), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n533), .A2(KEYINPUT75), .A3(new_n534), .A4(new_n536), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n520), .A2(new_n528), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n534), .A2(G902), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n539), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n252), .A2(new_n236), .A3(new_n253), .ZN(new_n546));
  XNOR2_X1  g360(.A(G134), .B(G137), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT65), .B1(new_n547), .B2(new_n248), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT65), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n241), .A2(G137), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n243), .A2(G134), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n549), .B(G131), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  AOI22_X1  g367(.A1(new_n425), .A2(new_n426), .B1(new_n192), .B2(KEYINPUT1), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n195), .B1(new_n554), .B2(new_n202), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n555), .A3(new_n249), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n546), .A2(KEYINPUT30), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n250), .A2(new_n235), .A3(new_n234), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n556), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT30), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT67), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT67), .ZN(new_n562));
  AOI211_X1 g376(.A(new_n562), .B(KEYINPUT30), .C1(new_n558), .C2(new_n556), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n293), .B(new_n557), .C1(new_n561), .C2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n546), .A2(new_n292), .A3(new_n556), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n260), .A2(G210), .A3(new_n363), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT27), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT26), .B(G101), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n564), .A2(new_n565), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT31), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n564), .A2(KEYINPUT31), .A3(new_n565), .A4(new_n569), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n565), .A2(KEYINPUT28), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT28), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n546), .A2(new_n575), .A3(new_n292), .A4(new_n556), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n559), .A2(new_n293), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n569), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n572), .A2(new_n573), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(G472), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(new_n188), .A3(KEYINPUT70), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT70), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n584), .B1(G472), .B2(G902), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT71), .B1(new_n579), .B2(new_n580), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n564), .A2(new_n565), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n580), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT29), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT71), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n577), .A2(new_n593), .A3(new_n578), .A4(new_n569), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n589), .A2(new_n591), .A3(new_n592), .A4(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n292), .B1(new_n546), .B2(new_n556), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n574), .B2(new_n576), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n580), .A2(new_n592), .ZN(new_n598));
  AOI21_X1  g412(.A(G902), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n588), .A2(KEYINPUT32), .B1(new_n600), .B2(G472), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT32), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n602), .B1(new_n581), .B2(new_n587), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n545), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n396), .A2(new_n397), .B1(new_n384), .B2(new_n417), .ZN(new_n605));
  OAI21_X1  g419(.A(G475), .B1(new_n605), .B2(G902), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n410), .B1(new_n409), .B2(new_n413), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n415), .A2(KEYINPUT20), .A3(new_n412), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n606), .B(new_n494), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n285), .A2(new_n287), .A3(new_n345), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT95), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n495), .A2(new_n604), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(G101), .ZN(G3));
  NAND2_X1  g427(.A1(new_n572), .A2(new_n573), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n579), .A2(new_n580), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n586), .ZN(new_n617));
  AOI21_X1  g431(.A(G902), .B1(new_n614), .B2(new_n615), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n617), .B1(new_n582), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n285), .A2(new_n287), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n619), .A2(new_n620), .A3(new_n545), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT96), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  INV_X1    g437(.A(new_n474), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n423), .B1(new_n472), .B2(new_n473), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n471), .A2(KEYINPUT33), .A3(new_n474), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n476), .A2(G902), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n628), .A2(new_n629), .B1(new_n476), .B2(new_n475), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n345), .A2(new_n491), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n421), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n622), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT34), .B(G104), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  NAND2_X1  g450(.A1(new_n478), .A2(new_n493), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n606), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT97), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n639), .B1(new_n607), .B2(new_n608), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n414), .A2(KEYINPUT97), .A3(new_n416), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n631), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n622), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT35), .B(G107), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  NAND2_X1  g462(.A1(new_n523), .A2(new_n527), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n499), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n543), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n539), .A2(new_n540), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n619), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n495), .A2(new_n611), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  AOI21_X1  g471(.A(new_n653), .B1(new_n601), .B2(new_n603), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n484), .B1(new_n488), .B2(G900), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n658), .A2(new_n346), .A3(new_n642), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  INV_X1    g475(.A(new_n344), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n341), .B1(new_n331), .B2(new_n339), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n664), .B(KEYINPUT38), .Z(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n637), .ZN(new_n667));
  NOR4_X1   g481(.A1(new_n666), .A2(new_n421), .A3(new_n667), .A4(new_n289), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n659), .B(KEYINPUT39), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n285), .A2(new_n287), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT40), .Z(new_n671));
  NAND3_X1  g485(.A1(new_n616), .A2(KEYINPUT32), .A3(new_n586), .ZN(new_n672));
  INV_X1    g486(.A(new_n570), .ZN(new_n673));
  INV_X1    g487(.A(new_n596), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n569), .B1(new_n674), .B2(new_n565), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n188), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(G472), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n672), .A2(new_n603), .A3(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n668), .A2(new_n653), .A3(new_n671), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G143), .ZN(G45));
  NAND2_X1  g494(.A1(new_n414), .A2(new_n416), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n630), .B1(new_n681), .B2(new_n606), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n658), .A2(new_n346), .A3(new_n682), .A4(new_n659), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G146), .ZN(G48));
  AND2_X1   g498(.A1(new_n278), .A2(new_n287), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n188), .B1(new_n274), .B2(new_n277), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n686), .A2(KEYINPUT98), .A3(G469), .ZN(new_n687));
  AOI21_X1  g501(.A(KEYINPUT98), .B1(new_n686), .B2(G469), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n685), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT99), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n686), .A2(G469), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT98), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n686), .A2(KEYINPUT98), .A3(G469), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(KEYINPUT99), .A3(new_n685), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n604), .A2(new_n632), .A3(new_n691), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  NAND2_X1  g514(.A1(new_n691), .A2(new_n697), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(new_n644), .A3(new_n604), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  INV_X1    g518(.A(new_n609), .ZN(new_n705));
  INV_X1    g519(.A(new_n345), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n689), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n658), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  OAI21_X1  g523(.A(KEYINPUT103), .B1(new_n421), .B2(new_n667), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT103), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n712), .A3(new_n637), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n586), .B(KEYINPUT100), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n577), .A2(new_n674), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT101), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n569), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n597), .A2(KEYINPUT101), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n715), .B1(new_n614), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n616), .A2(new_n188), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n721), .B1(new_n722), .B2(G472), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n539), .A2(new_n540), .A3(new_n544), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT102), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n572), .A2(new_n573), .B1(new_n718), .B2(new_n719), .ZN(new_n727));
  OAI22_X1  g541(.A1(new_n618), .A2(new_n582), .B1(new_n727), .B2(new_n715), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT102), .B1(new_n728), .B2(new_n545), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n702), .A2(new_n643), .A3(new_n714), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  INV_X1    g546(.A(new_n630), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n711), .A2(new_n733), .A3(new_n659), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT104), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n682), .A2(KEYINPUT104), .A3(new_n659), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n653), .A2(new_n728), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n736), .A2(new_n737), .A3(new_n707), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G125), .ZN(G27));
  AOI21_X1  g554(.A(KEYINPUT104), .B1(new_n682), .B2(new_n659), .ZN(new_n741));
  INV_X1    g555(.A(new_n659), .ZN(new_n742));
  NOR4_X1   g556(.A1(new_n421), .A2(new_n735), .A3(new_n630), .A4(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n617), .A2(KEYINPUT108), .A3(new_n602), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT108), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n603), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n601), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n748), .A2(new_n724), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n662), .A2(new_n663), .A3(new_n289), .ZN(new_n750));
  INV_X1    g564(.A(new_n287), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n284), .B(KEYINPUT105), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  AOI22_X1  g567(.A1(new_n279), .A2(new_n263), .B1(new_n281), .B2(new_n276), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n753), .B1(new_n754), .B2(G469), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n751), .B1(new_n755), .B2(new_n278), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT106), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n750), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AOI211_X1 g572(.A(KEYINPUT106), .B(new_n751), .C1(new_n755), .C2(new_n278), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n744), .A2(KEYINPUT42), .A3(new_n749), .A4(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT42), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n736), .A2(new_n760), .A3(new_n737), .A4(new_n604), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n762), .B1(new_n763), .B2(KEYINPUT107), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n600), .A2(G472), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n672), .A3(new_n603), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n724), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n768), .A2(new_n759), .A3(new_n758), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n765), .B1(new_n744), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n761), .B1(new_n764), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G131), .ZN(G33));
  NAND3_X1  g586(.A1(new_n769), .A2(new_n642), .A3(new_n659), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G134), .ZN(G36));
  NAND2_X1  g588(.A1(new_n421), .A2(new_n733), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT43), .Z(new_n776));
  INV_X1    g590(.A(new_n619), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n653), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n754), .A2(KEYINPUT45), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n754), .A2(KEYINPUT45), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(G469), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT46), .B1(new_n784), .B2(new_n752), .ZN(new_n785));
  INV_X1    g599(.A(new_n278), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n752), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n751), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n750), .B(KEYINPUT109), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n789), .A2(new_n669), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n776), .A2(KEYINPUT44), .A3(new_n778), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n781), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  INV_X1    g608(.A(new_n750), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n734), .A2(new_n767), .A3(new_n724), .A4(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n789), .A2(KEYINPUT47), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n789), .A2(KEYINPUT47), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  AND2_X1   g614(.A1(new_n776), .A2(new_n483), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n801), .A2(new_n730), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n665), .A2(new_n288), .A3(new_n689), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n802), .A2(KEYINPUT50), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT50), .B1(new_n802), .B2(new_n803), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n797), .A2(new_n798), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n696), .A2(new_n278), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n287), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n802), .B(new_n790), .C1(new_n807), .C2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n689), .A2(new_n795), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n801), .A2(new_n811), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n812), .A2(new_n653), .A3(new_n728), .ZN(new_n813));
  INV_X1    g627(.A(new_n811), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n814), .A2(new_n545), .A3(new_n484), .A4(new_n678), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n421), .A2(new_n630), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n813), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n806), .A2(new_n810), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n806), .A2(KEYINPUT51), .A3(new_n810), .A4(new_n818), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n802), .A2(new_n707), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n482), .B1(new_n815), .B2(new_n682), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n749), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT48), .B1(new_n812), .B2(new_n826), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n827), .B(KEYINPUT116), .Z(new_n828));
  NOR3_X1   g642(.A1(new_n812), .A2(KEYINPUT48), .A3(new_n826), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT115), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n825), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n821), .A2(new_n822), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT112), .ZN(new_n834));
  AOI211_X1 g648(.A(new_n751), .B(new_n742), .C1(new_n755), .C2(new_n278), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n678), .A2(new_n835), .A3(new_n653), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n834), .A2(new_n714), .A3(new_n345), .A4(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n706), .B1(new_n710), .B2(new_n713), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n834), .B1(new_n838), .B2(new_n836), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n739), .A2(new_n660), .A3(new_n683), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT52), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n841), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n843), .B(new_n844), .C1(new_n839), .C2(new_n837), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n604), .A2(new_n643), .A3(new_n642), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n698), .B(new_n708), .C1(new_n847), .C2(new_n701), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n725), .B1(new_n723), .B2(new_n724), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n728), .A2(new_n545), .A3(KEYINPUT102), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n421), .A2(KEYINPUT103), .A3(new_n667), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n712), .B1(new_n711), .B2(new_n637), .ZN(new_n852));
  OAI22_X1  g666(.A1(new_n849), .A2(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n691), .A2(new_n697), .A3(new_n643), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n606), .B(new_n637), .C1(new_n607), .C2(new_n608), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n856), .B1(new_n421), .B2(new_n630), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n621), .A2(new_n857), .A3(new_n643), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n612), .A2(new_n655), .A3(new_n858), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n848), .A2(new_n855), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n640), .A2(new_n641), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n667), .A2(new_n606), .A3(new_n659), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n620), .A2(new_n862), .A3(new_n795), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n658), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n760), .A2(new_n604), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n642), .A2(new_n659), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT111), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n736), .A2(new_n737), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n760), .A2(new_n738), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR4_X1   g685(.A1(new_n758), .A2(new_n759), .A3(new_n653), .A4(new_n728), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n744), .A2(KEYINPUT111), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n867), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n771), .A2(new_n860), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n833), .B1(new_n846), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT113), .ZN(new_n877));
  INV_X1    g691(.A(new_n846), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n844), .B1(new_n739), .B2(new_n660), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n879), .A2(new_n833), .A3(new_n859), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n771), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT114), .B1(new_n848), .B2(new_n855), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n698), .A2(new_n708), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT114), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n883), .A2(new_n731), .A3(new_n884), .A4(new_n703), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n882), .A2(new_n885), .A3(new_n874), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  AOI22_X1  g701(.A1(new_n876), .A2(new_n877), .B1(new_n878), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n889));
  OAI211_X1 g703(.A(KEYINPUT113), .B(new_n833), .C1(new_n846), .C2(new_n875), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n876), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n879), .A2(KEYINPUT53), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n846), .A2(new_n875), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT54), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  OAI22_X1  g710(.A1(new_n832), .A2(new_n896), .B1(G952), .B2(G953), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n808), .B(KEYINPUT49), .Z(new_n898));
  NAND3_X1  g712(.A1(new_n724), .A2(new_n287), .A3(new_n288), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT110), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n665), .A2(new_n775), .A3(new_n678), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n897), .A2(new_n902), .ZN(G75));
  NAND2_X1  g717(.A1(new_n876), .A2(new_n877), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n887), .A2(new_n878), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n905), .A3(new_n890), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(G210), .A3(G902), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n317), .A2(new_n330), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT117), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n328), .B(KEYINPUT55), .Z(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n907), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n912), .B1(new_n907), .B2(new_n908), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n260), .A2(G952), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(G51));
  XOR2_X1   g730(.A(new_n752), .B(KEYINPUT57), .Z(new_n917));
  AND4_X1   g731(.A1(new_n889), .A2(new_n904), .A3(new_n890), .A4(new_n905), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n889), .B1(new_n888), .B2(new_n890), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n259), .A2(new_n276), .ZN(new_n921));
  AOI22_X1  g735(.A1(new_n921), .A2(new_n263), .B1(new_n281), .B2(new_n273), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n906), .A2(G902), .ZN(new_n925));
  OR2_X1    g739(.A1(new_n925), .A2(new_n784), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n915), .B1(new_n924), .B2(new_n926), .ZN(G54));
  AND2_X1   g741(.A1(KEYINPUT58), .A2(G475), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n906), .A2(G902), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT118), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n929), .A2(new_n930), .A3(new_n415), .ZN(new_n931));
  INV_X1    g745(.A(new_n915), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n929), .B2(new_n415), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n930), .B1(new_n929), .B2(new_n415), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(G60));
  NAND2_X1  g749(.A1(G478), .A2(G902), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT59), .Z(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n628), .B1(new_n896), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n628), .A2(new_n938), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n906), .A2(KEYINPUT54), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n940), .B1(new_n941), .B2(new_n891), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n939), .A2(new_n915), .A3(new_n942), .ZN(G63));
  INV_X1    g757(.A(KEYINPUT61), .ZN(new_n944));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT60), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n888), .B2(new_n890), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n932), .B1(new_n947), .B2(new_n542), .ZN(new_n948));
  INV_X1    g762(.A(new_n946), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n651), .B(KEYINPUT119), .Z(new_n950));
  AND3_X1   g764(.A1(new_n906), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n944), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n906), .A2(new_n949), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n915), .B1(new_n953), .B2(new_n541), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n947), .A2(new_n950), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n954), .A2(KEYINPUT61), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n952), .A2(new_n956), .ZN(G66));
  OAI21_X1  g771(.A(G953), .B1(new_n489), .B2(new_n326), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT120), .ZN(new_n959));
  INV_X1    g773(.A(new_n860), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n959), .B1(new_n960), .B2(new_n260), .ZN(new_n961));
  INV_X1    g775(.A(G898), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n910), .B1(new_n962), .B2(new_n485), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n961), .B(new_n963), .ZN(G69));
  NAND2_X1  g778(.A1(new_n793), .A2(new_n799), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n768), .A2(new_n670), .A3(new_n795), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n857), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n679), .A2(new_n843), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n967), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n557), .B1(new_n561), .B2(new_n563), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT121), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(new_n405), .Z(new_n974));
  NOR2_X1   g788(.A1(new_n974), .A2(new_n485), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n260), .A2(G900), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT122), .Z(new_n978));
  NAND4_X1  g792(.A1(new_n789), .A2(new_n669), .A3(new_n749), .A4(new_n838), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n843), .A2(new_n773), .A3(new_n979), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n980), .A2(new_n793), .A3(new_n771), .A4(new_n799), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n978), .B1(new_n981), .B2(new_n260), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT123), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n974), .B1(new_n982), .B2(new_n983), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n976), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n260), .B1(G227), .B2(G900), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n986), .B(new_n987), .Z(G72));
  XOR2_X1   g802(.A(new_n590), .B(KEYINPUT126), .Z(new_n989));
  NAND4_X1  g803(.A1(new_n967), .A2(new_n860), .A3(new_n969), .A4(new_n970), .ZN(new_n990));
  XNOR2_X1  g804(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n991));
  NAND2_X1  g805(.A1(G472), .A2(G902), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT125), .Z(new_n994));
  AOI211_X1 g808(.A(new_n580), .B(new_n989), .C1(new_n990), .C2(new_n994), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n892), .A2(new_n894), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n591), .B(KEYINPUT127), .Z(new_n997));
  OAI21_X1  g811(.A(new_n993), .B1(new_n997), .B2(new_n673), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n994), .B1(new_n981), .B2(new_n960), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n1000), .A2(new_n580), .A3(new_n989), .ZN(new_n1001));
  NOR4_X1   g815(.A1(new_n995), .A2(new_n999), .A3(new_n915), .A4(new_n1001), .ZN(G57));
endmodule


