

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594;

  NAND2_X1 U325 ( .A1(n539), .A2(n549), .ZN(n293) );
  XOR2_X1 U326 ( .A(n357), .B(KEYINPUT9), .Z(n294) );
  INV_X1 U327 ( .A(KEYINPUT92), .ZN(n464) );
  XNOR2_X1 U328 ( .A(n464), .B(KEYINPUT25), .ZN(n465) );
  XNOR2_X1 U329 ( .A(n466), .B(n465), .ZN(n467) );
  INV_X1 U330 ( .A(n386), .ZN(n387) );
  XNOR2_X1 U331 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U332 ( .A(n322), .B(n321), .ZN(n328) );
  XNOR2_X1 U333 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U334 ( .A(n328), .B(n327), .ZN(n566) );
  INV_X1 U335 ( .A(G204GAT), .ZN(n455) );
  XOR2_X1 U336 ( .A(n397), .B(n396), .Z(n518) );
  XNOR2_X1 U337 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U338 ( .A(n478), .B(KEYINPUT102), .ZN(n479) );
  XNOR2_X1 U339 ( .A(n481), .B(G43GAT), .ZN(n482) );
  XNOR2_X1 U340 ( .A(n458), .B(n457), .ZN(G1353GAT) );
  XNOR2_X1 U341 ( .A(n480), .B(n479), .ZN(G1331GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n296) );
  XNOR2_X1 U343 ( .A(KEYINPUT31), .B(KEYINPUT73), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n310) );
  XOR2_X1 U345 ( .A(G176GAT), .B(G64GAT), .Z(n386) );
  XOR2_X1 U346 ( .A(KEYINPUT71), .B(n386), .Z(n298) );
  XOR2_X1 U347 ( .A(G148GAT), .B(G78GAT), .Z(n423) );
  XNOR2_X1 U348 ( .A(G204GAT), .B(n423), .ZN(n297) );
  XNOR2_X1 U349 ( .A(n298), .B(n297), .ZN(n303) );
  XNOR2_X1 U350 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n299), .B(KEYINPUT70), .ZN(n332) );
  XOR2_X1 U352 ( .A(KEYINPUT74), .B(n332), .Z(n301) );
  NAND2_X1 U353 ( .A1(G230GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U354 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U355 ( .A(n303), .B(n302), .Z(n308) );
  XOR2_X1 U356 ( .A(G120GAT), .B(G71GAT), .Z(n433) );
  XOR2_X1 U357 ( .A(KEYINPUT72), .B(G92GAT), .Z(n305) );
  XNOR2_X1 U358 ( .A(G99GAT), .B(G85GAT), .ZN(n304) );
  XNOR2_X1 U359 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U360 ( .A(G106GAT), .B(n306), .Z(n326) );
  XNOR2_X1 U361 ( .A(n433), .B(n326), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n310), .B(n309), .ZN(n459) );
  INV_X1 U364 ( .A(n459), .ZN(n454) );
  INV_X1 U365 ( .A(G43GAT), .ZN(n311) );
  NAND2_X1 U366 ( .A1(G29GAT), .A2(n311), .ZN(n314) );
  INV_X1 U367 ( .A(G29GAT), .ZN(n312) );
  NAND2_X1 U368 ( .A1(n312), .A2(G43GAT), .ZN(n313) );
  NAND2_X1 U369 ( .A1(n314), .A2(n313), .ZN(n316) );
  XNOR2_X1 U370 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n315) );
  XNOR2_X1 U371 ( .A(n316), .B(n315), .ZN(n357) );
  NAND2_X1 U372 ( .A1(G232GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U373 ( .A(n294), .B(n317), .ZN(n322) );
  XOR2_X1 U374 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n320) );
  XOR2_X1 U375 ( .A(G50GAT), .B(G162GAT), .Z(n429) );
  XNOR2_X1 U376 ( .A(G36GAT), .B(G190GAT), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n318), .B(G218GAT), .ZN(n380) );
  XNOR2_X1 U378 ( .A(n429), .B(n380), .ZN(n319) );
  XNOR2_X1 U379 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U380 ( .A(KEYINPUT76), .B(KEYINPUT10), .Z(n324) );
  XNOR2_X1 U381 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n323) );
  XNOR2_X1 U382 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U384 ( .A(n566), .B(KEYINPUT79), .Z(n549) );
  XNOR2_X1 U385 ( .A(KEYINPUT36), .B(n549), .ZN(n591) );
  XOR2_X1 U386 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n334) );
  XOR2_X1 U387 ( .A(KEYINPUT80), .B(KEYINPUT15), .Z(n330) );
  XNOR2_X1 U388 ( .A(G8GAT), .B(G64GAT), .ZN(n329) );
  XNOR2_X1 U389 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U390 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U391 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U392 ( .A(G22GAT), .B(G155GAT), .Z(n424) );
  XOR2_X1 U393 ( .A(G15GAT), .B(G127GAT), .Z(n434) );
  XOR2_X1 U394 ( .A(n424), .B(n434), .Z(n336) );
  NAND2_X1 U395 ( .A1(G231GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U397 ( .A(n338), .B(n337), .Z(n343) );
  XOR2_X1 U398 ( .A(G1GAT), .B(KEYINPUT69), .Z(n360) );
  XOR2_X1 U399 ( .A(G78GAT), .B(G211GAT), .Z(n340) );
  XNOR2_X1 U400 ( .A(G183GAT), .B(G71GAT), .ZN(n339) );
  XNOR2_X1 U401 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n360), .B(n341), .ZN(n342) );
  XOR2_X1 U403 ( .A(n343), .B(n342), .Z(n491) );
  INV_X1 U404 ( .A(n491), .ZN(n587) );
  NAND2_X1 U405 ( .A1(n591), .A2(n587), .ZN(n345) );
  XNOR2_X1 U406 ( .A(KEYINPUT45), .B(KEYINPUT108), .ZN(n344) );
  XNOR2_X1 U407 ( .A(n345), .B(n344), .ZN(n346) );
  NOR2_X1 U408 ( .A1(n454), .A2(n346), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n347), .B(KEYINPUT109), .ZN(n366) );
  XOR2_X1 U410 ( .A(KEYINPUT68), .B(G141GAT), .Z(n349) );
  XNOR2_X1 U411 ( .A(G197GAT), .B(G22GAT), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U413 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n351) );
  XNOR2_X1 U414 ( .A(KEYINPUT29), .B(KEYINPUT66), .ZN(n350) );
  XNOR2_X1 U415 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U416 ( .A(n353), .B(n352), .ZN(n365) );
  XOR2_X1 U417 ( .A(G113GAT), .B(G15GAT), .Z(n355) );
  XNOR2_X1 U418 ( .A(G36GAT), .B(G50GAT), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U420 ( .A(G169GAT), .B(G8GAT), .Z(n385) );
  XOR2_X1 U421 ( .A(n356), .B(n385), .Z(n363) );
  XOR2_X1 U422 ( .A(n357), .B(KEYINPUT67), .Z(n359) );
  NAND2_X1 U423 ( .A1(G229GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U424 ( .A(n359), .B(n358), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n365), .B(n364), .ZN(n582) );
  NOR2_X1 U428 ( .A1(n366), .A2(n582), .ZN(n367) );
  XOR2_X1 U429 ( .A(KEYINPUT110), .B(n367), .Z(n375) );
  XOR2_X1 U430 ( .A(KEYINPUT46), .B(KEYINPUT106), .Z(n369) );
  XOR2_X1 U431 ( .A(KEYINPUT41), .B(n454), .Z(n576) );
  NAND2_X1 U432 ( .A1(n576), .A2(n582), .ZN(n368) );
  XNOR2_X1 U433 ( .A(n369), .B(n368), .ZN(n370) );
  NOR2_X1 U434 ( .A1(n370), .A2(n587), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n371), .B(KEYINPUT107), .ZN(n372) );
  NOR2_X1 U436 ( .A1(n566), .A2(n372), .ZN(n373) );
  XNOR2_X1 U437 ( .A(KEYINPUT47), .B(n373), .ZN(n374) );
  NAND2_X1 U438 ( .A1(n375), .A2(n374), .ZN(n377) );
  XNOR2_X1 U439 ( .A(KEYINPUT111), .B(KEYINPUT48), .ZN(n376) );
  XNOR2_X1 U440 ( .A(n377), .B(n376), .ZN(n555) );
  XOR2_X1 U441 ( .A(KEYINPUT87), .B(KEYINPUT89), .Z(n379) );
  XNOR2_X1 U442 ( .A(G92GAT), .B(KEYINPUT86), .ZN(n378) );
  XNOR2_X1 U443 ( .A(n379), .B(n378), .ZN(n392) );
  XOR2_X1 U444 ( .A(n380), .B(KEYINPUT88), .Z(n382) );
  NAND2_X1 U445 ( .A1(G226GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n382), .B(n381), .ZN(n390) );
  XOR2_X1 U447 ( .A(G183GAT), .B(KEYINPUT18), .Z(n384) );
  XNOR2_X1 U448 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n383) );
  XNOR2_X1 U449 ( .A(n384), .B(n383), .ZN(n437) );
  XNOR2_X1 U450 ( .A(n385), .B(n437), .ZN(n388) );
  XNOR2_X1 U451 ( .A(n392), .B(n391), .ZN(n397) );
  XOR2_X1 U452 ( .A(KEYINPUT21), .B(G211GAT), .Z(n394) );
  XNOR2_X1 U453 ( .A(KEYINPUT84), .B(G204GAT), .ZN(n393) );
  XNOR2_X1 U454 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U455 ( .A(G197GAT), .B(n395), .ZN(n430) );
  INV_X1 U456 ( .A(n430), .ZN(n396) );
  NOR2_X1 U457 ( .A1(n555), .A2(n518), .ZN(n398) );
  XNOR2_X1 U458 ( .A(n398), .B(KEYINPUT54), .ZN(n416) );
  XOR2_X1 U459 ( .A(G57GAT), .B(G155GAT), .Z(n400) );
  XNOR2_X1 U460 ( .A(G120GAT), .B(G148GAT), .ZN(n399) );
  XNOR2_X1 U461 ( .A(n400), .B(n399), .ZN(n415) );
  XOR2_X1 U462 ( .A(G85GAT), .B(G162GAT), .Z(n402) );
  XNOR2_X1 U463 ( .A(G29GAT), .B(G127GAT), .ZN(n401) );
  XNOR2_X1 U464 ( .A(n402), .B(n401), .ZN(n407) );
  XNOR2_X1 U465 ( .A(G113GAT), .B(G134GAT), .ZN(n403) );
  XNOR2_X1 U466 ( .A(n403), .B(KEYINPUT0), .ZN(n435) );
  XOR2_X1 U467 ( .A(n435), .B(KEYINPUT6), .Z(n405) );
  NAND2_X1 U468 ( .A1(G225GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U470 ( .A(n407), .B(n406), .Z(n413) );
  XNOR2_X1 U471 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n408) );
  XNOR2_X1 U472 ( .A(n408), .B(KEYINPUT2), .ZN(n417) );
  XOR2_X1 U473 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n410) );
  XNOR2_X1 U474 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n409) );
  XNOR2_X1 U475 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U476 ( .A(n417), .B(n411), .ZN(n412) );
  XNOR2_X1 U477 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U478 ( .A(n415), .B(n414), .Z(n530) );
  INV_X1 U479 ( .A(n530), .ZN(n556) );
  NAND2_X1 U480 ( .A1(n416), .A2(n556), .ZN(n484) );
  XOR2_X1 U481 ( .A(n417), .B(KEYINPUT23), .Z(n422) );
  XOR2_X1 U482 ( .A(KEYINPUT22), .B(KEYINPUT85), .Z(n419) );
  XNOR2_X1 U483 ( .A(G218GAT), .B(G106GAT), .ZN(n418) );
  XNOR2_X1 U484 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U485 ( .A(n420), .B(KEYINPUT24), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n422), .B(n421), .ZN(n428) );
  XOR2_X1 U487 ( .A(n424), .B(n423), .Z(n426) );
  NAND2_X1 U488 ( .A1(G228GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U490 ( .A(n428), .B(n427), .Z(n432) );
  XOR2_X1 U491 ( .A(n430), .B(n429), .Z(n431) );
  XNOR2_X1 U492 ( .A(n432), .B(n431), .ZN(n485) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n436) );
  XNOR2_X1 U494 ( .A(n436), .B(n435), .ZN(n441) );
  XOR2_X1 U495 ( .A(G169GAT), .B(n437), .Z(n439) );
  NAND2_X1 U496 ( .A1(G227GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U497 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U498 ( .A(n441), .B(n440), .Z(n449) );
  XOR2_X1 U499 ( .A(KEYINPUT82), .B(G99GAT), .Z(n443) );
  XNOR2_X1 U500 ( .A(G43GAT), .B(G190GAT), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n443), .B(n442), .ZN(n447) );
  XOR2_X1 U502 ( .A(G176GAT), .B(KEYINPUT64), .Z(n445) );
  XNOR2_X1 U503 ( .A(KEYINPUT83), .B(KEYINPUT20), .ZN(n444) );
  XNOR2_X1 U504 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U506 ( .A(n449), .B(n448), .Z(n539) );
  INV_X1 U507 ( .A(n539), .ZN(n571) );
  NAND2_X1 U508 ( .A1(n485), .A2(n571), .ZN(n450) );
  XNOR2_X1 U509 ( .A(n450), .B(KEYINPUT90), .ZN(n451) );
  XNOR2_X1 U510 ( .A(KEYINPUT26), .B(n451), .ZN(n461) );
  NOR2_X1 U511 ( .A1(n484), .A2(n461), .ZN(n453) );
  INV_X1 U512 ( .A(KEYINPUT123), .ZN(n452) );
  XNOR2_X1 U513 ( .A(n453), .B(n452), .ZN(n590) );
  NAND2_X1 U514 ( .A1(n590), .A2(n454), .ZN(n458) );
  XOR2_X1 U515 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n456) );
  XNOR2_X1 U516 ( .A(n485), .B(KEYINPUT28), .ZN(n536) );
  INV_X1 U517 ( .A(n536), .ZN(n524) );
  XNOR2_X1 U518 ( .A(KEYINPUT38), .B(KEYINPUT97), .ZN(n477) );
  NAND2_X1 U519 ( .A1(n459), .A2(n582), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n460), .B(KEYINPUT75), .ZN(n496) );
  INV_X1 U521 ( .A(n518), .ZN(n532) );
  XOR2_X1 U522 ( .A(KEYINPUT27), .B(n532), .Z(n471) );
  NOR2_X1 U523 ( .A1(n471), .A2(n461), .ZN(n557) );
  NOR2_X1 U524 ( .A1(n571), .A2(n518), .ZN(n462) );
  XOR2_X1 U525 ( .A(KEYINPUT91), .B(n462), .Z(n463) );
  NOR2_X1 U526 ( .A1(n485), .A2(n463), .ZN(n466) );
  NOR2_X1 U527 ( .A1(n557), .A2(n467), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n468), .B(KEYINPUT93), .ZN(n469) );
  NAND2_X1 U529 ( .A1(n469), .A2(n556), .ZN(n473) );
  NAND2_X1 U530 ( .A1(n530), .A2(n524), .ZN(n470) );
  NOR2_X1 U531 ( .A1(n471), .A2(n470), .ZN(n540) );
  NAND2_X1 U532 ( .A1(n571), .A2(n540), .ZN(n472) );
  NAND2_X1 U533 ( .A1(n473), .A2(n472), .ZN(n495) );
  AND2_X1 U534 ( .A1(n491), .A2(n591), .ZN(n474) );
  AND2_X1 U535 ( .A1(n495), .A2(n474), .ZN(n475) );
  XOR2_X1 U536 ( .A(KEYINPUT37), .B(n475), .Z(n527) );
  AND2_X1 U537 ( .A1(n496), .A2(n527), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n477), .B(n476), .ZN(n510) );
  NOR2_X1 U539 ( .A1(n524), .A2(n510), .ZN(n480) );
  INV_X1 U540 ( .A(G50GAT), .ZN(n478) );
  NOR2_X1 U541 ( .A1(n571), .A2(n510), .ZN(n483) );
  XNOR2_X1 U542 ( .A(KEYINPUT40), .B(KEYINPUT101), .ZN(n481) );
  XNOR2_X1 U543 ( .A(n483), .B(n482), .ZN(G1330GAT) );
  NOR2_X1 U544 ( .A1(n485), .A2(n484), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n486), .B(KEYINPUT55), .ZN(n570) );
  NOR2_X1 U546 ( .A1(n570), .A2(n293), .ZN(n488) );
  XNOR2_X1 U547 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(n490) );
  INV_X1 U549 ( .A(G190GAT), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(G1351GAT) );
  NOR2_X1 U551 ( .A1(n549), .A2(n491), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n492), .B(KEYINPUT81), .ZN(n493) );
  XOR2_X1 U553 ( .A(KEYINPUT16), .B(n493), .Z(n494) );
  AND2_X1 U554 ( .A1(n495), .A2(n494), .ZN(n515) );
  NAND2_X1 U555 ( .A1(n496), .A2(n515), .ZN(n504) );
  NOR2_X1 U556 ( .A1(n556), .A2(n504), .ZN(n497) );
  XOR2_X1 U557 ( .A(KEYINPUT34), .B(n497), .Z(n498) );
  XNOR2_X1 U558 ( .A(G1GAT), .B(n498), .ZN(G1324GAT) );
  NOR2_X1 U559 ( .A1(n518), .A2(n504), .ZN(n499) );
  XOR2_X1 U560 ( .A(KEYINPUT94), .B(n499), .Z(n500) );
  XNOR2_X1 U561 ( .A(G8GAT), .B(n500), .ZN(G1325GAT) );
  NOR2_X1 U562 ( .A1(n571), .A2(n504), .ZN(n502) );
  XNOR2_X1 U563 ( .A(KEYINPUT95), .B(KEYINPUT35), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U565 ( .A(G15GAT), .B(n503), .Z(G1326GAT) );
  NOR2_X1 U566 ( .A1(n524), .A2(n504), .ZN(n505) );
  XOR2_X1 U567 ( .A(G22GAT), .B(n505), .Z(G1327GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT96), .B(KEYINPUT39), .Z(n507) );
  XNOR2_X1 U569 ( .A(G29GAT), .B(KEYINPUT98), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n507), .B(n506), .ZN(n509) );
  NOR2_X1 U571 ( .A1(n510), .A2(n556), .ZN(n508) );
  XOR2_X1 U572 ( .A(n509), .B(n508), .Z(G1328GAT) );
  NOR2_X1 U573 ( .A1(n510), .A2(n518), .ZN(n512) );
  XNOR2_X1 U574 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U576 ( .A(G36GAT), .B(n513), .ZN(G1329GAT) );
  INV_X1 U577 ( .A(n576), .ZN(n514) );
  NOR2_X1 U578 ( .A1(n582), .A2(n514), .ZN(n528) );
  NAND2_X1 U579 ( .A1(n528), .A2(n515), .ZN(n523) );
  NOR2_X1 U580 ( .A1(n556), .A2(n523), .ZN(n516) );
  XOR2_X1 U581 ( .A(G57GAT), .B(n516), .Z(n517) );
  XNOR2_X1 U582 ( .A(KEYINPUT42), .B(n517), .ZN(G1332GAT) );
  NOR2_X1 U583 ( .A1(n518), .A2(n523), .ZN(n520) );
  XNOR2_X1 U584 ( .A(G64GAT), .B(KEYINPUT103), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(G1333GAT) );
  NOR2_X1 U586 ( .A1(n571), .A2(n523), .ZN(n521) );
  XOR2_X1 U587 ( .A(KEYINPUT104), .B(n521), .Z(n522) );
  XNOR2_X1 U588 ( .A(G71GAT), .B(n522), .ZN(G1334GAT) );
  NOR2_X1 U589 ( .A1(n524), .A2(n523), .ZN(n526) );
  XNOR2_X1 U590 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(G1335GAT) );
  NAND2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n529), .B(KEYINPUT105), .ZN(n535) );
  NAND2_X1 U594 ( .A1(n530), .A2(n535), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G85GAT), .B(n531), .ZN(G1336GAT) );
  NAND2_X1 U596 ( .A1(n532), .A2(n535), .ZN(n533) );
  XNOR2_X1 U597 ( .A(G92GAT), .B(n533), .ZN(G1337GAT) );
  NAND2_X1 U598 ( .A1(n539), .A2(n535), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n534), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n537), .B(KEYINPUT44), .ZN(n538) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(n538), .ZN(G1339GAT) );
  NAND2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U604 ( .A1(n555), .A2(n541), .ZN(n550) );
  NAND2_X1 U605 ( .A1(n550), .A2(n582), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n542), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT112), .B(KEYINPUT49), .Z(n544) );
  NAND2_X1 U608 ( .A1(n550), .A2(n576), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G120GAT), .B(n545), .ZN(G1341GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n547) );
  NAND2_X1 U612 ( .A1(n550), .A2(n587), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n552) );
  NAND2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n554) );
  XOR2_X1 U618 ( .A(G134GAT), .B(KEYINPUT115), .Z(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1343GAT) );
  XOR2_X1 U620 ( .A(G141GAT), .B(KEYINPUT117), .Z(n561) );
  NOR2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U623 ( .A(KEYINPUT116), .B(n559), .Z(n567) );
  NAND2_X1 U624 ( .A1(n582), .A2(n567), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n561), .B(n560), .ZN(G1344GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n563) );
  NAND2_X1 U627 ( .A1(n576), .A2(n567), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U629 ( .A(G148GAT), .B(n564), .ZN(G1345GAT) );
  NAND2_X1 U630 ( .A1(n567), .A2(n587), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n568), .B(KEYINPUT118), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G162GAT), .B(n569), .ZN(G1347GAT) );
  NOR2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n579) );
  NAND2_X1 U636 ( .A1(n579), .A2(n582), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT57), .B(KEYINPUT120), .Z(n574) );
  XNOR2_X1 U639 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U641 ( .A(KEYINPUT119), .B(n575), .Z(n578) );
  NAND2_X1 U642 ( .A1(n579), .A2(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1349GAT) );
  XOR2_X1 U644 ( .A(G183GAT), .B(KEYINPUT121), .Z(n581) );
  NAND2_X1 U645 ( .A1(n579), .A2(n587), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1350GAT) );
  NAND2_X1 U647 ( .A1(n590), .A2(n582), .ZN(n586) );
  XOR2_X1 U648 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n584) );
  XNOR2_X1 U649 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1352GAT) );
  NAND2_X1 U652 ( .A1(n590), .A2(n587), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(KEYINPUT126), .ZN(n589) );
  XNOR2_X1 U654 ( .A(G211GAT), .B(n589), .ZN(G1354GAT) );
  NAND2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n593) );
  XOR2_X1 U656 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(n594), .B(G218GAT), .ZN(G1355GAT) );
endmodule

