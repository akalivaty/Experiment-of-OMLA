

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777;

  XNOR2_X1 U373 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U374 ( .A(n649), .B(n651), .ZN(n652) );
  BUF_X1 U375 ( .A(n636), .Z(n665) );
  XNOR2_X1 U376 ( .A(n625), .B(n624), .ZN(n721) );
  XNOR2_X1 U377 ( .A(G137), .B(G113), .ZN(n503) );
  XNOR2_X1 U378 ( .A(G140), .B(G143), .ZN(n471) );
  XOR2_X1 U379 ( .A(KEYINPUT84), .B(G110), .Z(n531) );
  AND2_X1 U380 ( .A1(n721), .A2(n656), .ZN(n350) );
  AND2_X2 U381 ( .A1(n389), .A2(n390), .ZN(n381) );
  NOR2_X1 U382 ( .A1(n758), .A2(n623), .ZN(n405) );
  XNOR2_X2 U383 ( .A(n368), .B(n361), .ZN(n757) );
  INV_X2 U384 ( .A(G953), .ZN(n770) );
  XNOR2_X1 U385 ( .A(n637), .B(KEYINPUT69), .ZN(n364) );
  NAND2_X1 U386 ( .A1(n407), .A2(n406), .ZN(n728) );
  NOR2_X1 U387 ( .A1(n358), .A2(n425), .ZN(n407) );
  XNOR2_X1 U388 ( .A(n496), .B(n423), .ZN(n672) );
  BUF_X1 U389 ( .A(n357), .Z(n374) );
  NAND2_X1 U390 ( .A1(n435), .A2(n441), .ZN(n367) );
  NAND2_X1 U391 ( .A1(n364), .A2(n639), .ZN(n363) );
  XNOR2_X1 U392 ( .A(n713), .B(G128), .ZN(G30) );
  XNOR2_X1 U393 ( .A(n582), .B(KEYINPUT40), .ZN(n351) );
  NAND2_X1 U394 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U395 ( .A(n579), .B(KEYINPUT39), .ZN(n581) );
  XNOR2_X1 U396 ( .A(n621), .B(KEYINPUT104), .ZN(n706) );
  NAND2_X1 U397 ( .A1(n609), .A2(n355), .ZN(n656) );
  INV_X1 U398 ( .A(n630), .ZN(n609) );
  XNOR2_X1 U399 ( .A(n352), .B(KEYINPUT81), .ZN(n578) );
  NOR2_X1 U400 ( .A1(n420), .A2(n628), .ZN(n419) );
  NAND2_X1 U401 ( .A1(n353), .A2(n542), .ZN(n352) );
  XNOR2_X1 U402 ( .A(n617), .B(n541), .ZN(n353) );
  NAND2_X1 U403 ( .A1(n434), .A2(n555), .ZN(n617) );
  XNOR2_X1 U404 ( .A(n470), .B(KEYINPUT72), .ZN(n551) );
  NAND2_X2 U405 ( .A1(n412), .A2(n408), .ZN(n735) );
  AND2_X1 U406 ( .A1(n398), .A2(KEYINPUT1), .ZN(n358) );
  XNOR2_X1 U407 ( .A(n458), .B(n457), .ZN(n540) );
  XOR2_X1 U408 ( .A(KEYINPUT62), .B(n666), .Z(n667) );
  OR2_X1 U409 ( .A1(n701), .A2(n428), .ZN(n427) );
  XNOR2_X1 U410 ( .A(n537), .B(n536), .ZN(n701) );
  XNOR2_X1 U411 ( .A(n672), .B(G146), .ZN(n415) );
  XNOR2_X1 U412 ( .A(n424), .B(G131), .ZN(n496) );
  XNOR2_X1 U413 ( .A(G128), .B(KEYINPUT24), .ZN(n446) );
  XNOR2_X1 U414 ( .A(G134), .B(KEYINPUT71), .ZN(n423) );
  NAND2_X1 U415 ( .A1(n351), .A2(n661), .ZN(n584) );
  XNOR2_X1 U416 ( .A(n351), .B(n664), .ZN(G33) );
  XNOR2_X2 U417 ( .A(G146), .B(G125), .ZN(n513) );
  XNOR2_X1 U418 ( .A(n590), .B(n569), .ZN(n745) );
  XNOR2_X1 U419 ( .A(n419), .B(KEYINPUT33), .ZN(n758) );
  XNOR2_X1 U420 ( .A(n688), .B(n354), .ZN(n689) );
  AND2_X1 U421 ( .A1(n372), .A2(G478), .ZN(n354) );
  AND2_X1 U422 ( .A1(n629), .A2(n628), .ZN(n355) );
  NAND2_X1 U423 ( .A1(n365), .A2(n363), .ZN(n356) );
  NAND2_X1 U424 ( .A1(n365), .A2(n363), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n512), .B(n514), .ZN(n386) );
  XNOR2_X1 U426 ( .A(n416), .B(n415), .ZN(n537) );
  XNOR2_X1 U427 ( .A(n356), .B(KEYINPUT45), .ZN(n357) );
  XNOR2_X1 U428 ( .A(n362), .B(KEYINPUT45), .ZN(n645) );
  AND2_X1 U429 ( .A1(n556), .A2(n555), .ZN(n574) );
  NAND2_X1 U430 ( .A1(n401), .A2(n400), .ZN(n638) );
  INV_X1 U431 ( .A(n658), .ZN(n400) );
  INV_X2 U432 ( .A(KEYINPUT70), .ZN(n424) );
  INV_X1 U433 ( .A(G237), .ZN(n525) );
  XNOR2_X1 U434 ( .A(n478), .B(n477), .ZN(n479) );
  OR2_X1 U435 ( .A1(n666), .A2(n409), .ZN(n408) );
  AND2_X1 U436 ( .A1(n414), .A2(n413), .ZN(n412) );
  NAND2_X1 U437 ( .A1(n411), .A2(n410), .ZN(n409) );
  NAND2_X1 U438 ( .A1(n432), .A2(n431), .ZN(n398) );
  NAND2_X1 U439 ( .A1(G902), .A2(G469), .ZN(n431) );
  INV_X1 U440 ( .A(KEYINPUT94), .ZN(n633) );
  NAND2_X1 U441 ( .A1(n429), .A2(n410), .ZN(n428) );
  INV_X1 U442 ( .A(G469), .ZN(n429) );
  XNOR2_X1 U443 ( .A(G116), .B(G119), .ZN(n499) );
  XNOR2_X1 U444 ( .A(KEYINPUT73), .B(KEYINPUT3), .ZN(n519) );
  XNOR2_X1 U445 ( .A(G116), .B(G107), .ZN(n520) );
  AND2_X1 U446 ( .A1(n644), .A2(n391), .ZN(n390) );
  NOR2_X1 U447 ( .A1(n641), .A2(n640), .ZN(n392) );
  NOR2_X1 U448 ( .A1(G953), .A2(G237), .ZN(n502) );
  INV_X1 U449 ( .A(G101), .ZN(n498) );
  XNOR2_X1 U450 ( .A(n513), .B(n385), .ZN(n384) );
  INV_X1 U451 ( .A(KEYINPUT97), .ZN(n385) );
  INV_X1 U452 ( .A(KEYINPUT48), .ZN(n436) );
  NAND2_X1 U453 ( .A1(G234), .A2(G237), .ZN(n459) );
  OR2_X1 U454 ( .A1(n540), .A2(n469), .ZN(n470) );
  INV_X1 U455 ( .A(KEYINPUT113), .ZN(n369) );
  NAND2_X1 U456 ( .A1(n745), .A2(n744), .ZN(n370) );
  NAND2_X1 U457 ( .A1(n728), .A2(n727), .ZN(n420) );
  INV_X1 U458 ( .A(n510), .ZN(n411) );
  NAND2_X1 U459 ( .A1(n510), .A2(G902), .ZN(n413) );
  XNOR2_X1 U460 ( .A(KEYINPUT99), .B(KEYINPUT23), .ZN(n447) );
  XNOR2_X1 U461 ( .A(G122), .B(G134), .ZN(n485) );
  XNOR2_X1 U462 ( .A(G104), .B(G107), .ZN(n530) );
  XNOR2_X1 U463 ( .A(G137), .B(G140), .ZN(n533) );
  BUF_X1 U464 ( .A(n758), .Z(n397) );
  XNOR2_X1 U465 ( .A(n614), .B(KEYINPUT35), .ZN(n615) );
  BUF_X1 U466 ( .A(n540), .Z(n732) );
  XNOR2_X1 U467 ( .A(n484), .B(n483), .ZN(n570) );
  XNOR2_X1 U468 ( .A(n482), .B(n481), .ZN(n483) );
  BUF_X1 U469 ( .A(n728), .Z(n399) );
  INV_X1 U470 ( .A(KEYINPUT42), .ZN(n403) );
  XNOR2_X1 U471 ( .A(n421), .B(n606), .ZN(n663) );
  AND2_X1 U472 ( .A1(n605), .A2(n602), .ZN(n422) );
  NAND2_X1 U473 ( .A1(n599), .A2(n396), .ZN(n625) );
  INV_X1 U474 ( .A(n738), .ZN(n396) );
  INV_X1 U475 ( .A(KEYINPUT56), .ZN(n394) );
  NAND2_X1 U476 ( .A1(n638), .A2(KEYINPUT44), .ZN(n359) );
  INV_X1 U477 ( .A(G902), .ZN(n410) );
  AND2_X1 U478 ( .A1(n427), .A2(n426), .ZN(n360) );
  INV_X1 U479 ( .A(KEYINPUT1), .ZN(n426) );
  XOR2_X1 U480 ( .A(n573), .B(KEYINPUT41), .Z(n361) );
  INV_X1 U481 ( .A(n722), .ZN(n433) );
  XNOR2_X2 U482 ( .A(n366), .B(KEYINPUT93), .ZN(n365) );
  NAND2_X1 U483 ( .A1(n635), .A2(n359), .ZN(n366) );
  NOR2_X1 U484 ( .A1(n367), .A2(n725), .ZN(n646) );
  XNOR2_X2 U485 ( .A(n367), .B(n592), .ZN(n678) );
  NOR2_X2 U486 ( .A1(n743), .A2(n746), .ZN(n368) );
  XNOR2_X2 U487 ( .A(n370), .B(n369), .ZN(n743) );
  XNOR2_X1 U488 ( .A(n424), .B(G131), .ZN(n371) );
  BUF_X1 U489 ( .A(n546), .Z(n590) );
  XNOR2_X1 U490 ( .A(n378), .B(n647), .ZN(n372) );
  NAND2_X2 U491 ( .A1(n379), .A2(n388), .ZN(n378) );
  INV_X1 U492 ( .A(n393), .ZN(n373) );
  INV_X1 U493 ( .A(n724), .ZN(n393) );
  NAND2_X1 U494 ( .A1(n374), .A2(n646), .ZN(n375) );
  NAND2_X1 U495 ( .A1(n357), .A2(n646), .ZN(n382) );
  BUF_X1 U496 ( .A(n557), .Z(n376) );
  XNOR2_X1 U497 ( .A(n386), .B(n384), .ZN(n383) );
  XNOR2_X1 U498 ( .A(n375), .B(KEYINPUT80), .ZN(n377) );
  XNOR2_X1 U499 ( .A(n382), .B(KEYINPUT80), .ZN(n388) );
  XNOR2_X2 U500 ( .A(n378), .B(n647), .ZN(n698) );
  NAND2_X1 U501 ( .A1(n393), .A2(n392), .ZN(n380) );
  XNOR2_X1 U502 ( .A(n416), .B(n383), .ZN(n523) );
  NAND2_X1 U503 ( .A1(n381), .A2(n380), .ZN(n379) );
  XNOR2_X2 U504 ( .A(n671), .B(n498), .ZN(n416) );
  XNOR2_X2 U505 ( .A(n497), .B(n387), .ZN(n671) );
  XNOR2_X2 U506 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n387) );
  XNOR2_X2 U507 ( .A(G143), .B(G128), .ZN(n497) );
  NAND2_X1 U508 ( .A1(n377), .A2(n726), .ZN(n762) );
  NAND2_X1 U509 ( .A1(n724), .A2(n640), .ZN(n389) );
  NAND2_X1 U510 ( .A1(n641), .A2(n640), .ZN(n391) );
  NAND2_X1 U511 ( .A1(n645), .A2(n678), .ZN(n724) );
  XNOR2_X1 U512 ( .A(n395), .B(n394), .ZN(G51) );
  NAND2_X1 U513 ( .A1(n655), .A2(n694), .ZN(n395) );
  XNOR2_X2 U514 ( .A(n616), .B(n615), .ZN(n636) );
  NAND2_X1 U515 ( .A1(n350), .A2(n706), .ZN(n439) );
  XNOR2_X1 U516 ( .A(n451), .B(n676), .ZN(n686) );
  INV_X1 U517 ( .A(n610), .ZN(n434) );
  XNOR2_X1 U518 ( .A(n405), .B(KEYINPUT34), .ZN(n613) );
  INV_X1 U519 ( .A(n398), .ZN(n430) );
  INV_X1 U520 ( .A(n663), .ZN(n401) );
  NAND2_X1 U521 ( .A1(n609), .A2(n422), .ZN(n421) );
  XNOR2_X1 U522 ( .A(n402), .B(n450), .ZN(n451) );
  XNOR2_X1 U523 ( .A(n449), .B(n448), .ZN(n402) );
  XNOR2_X2 U524 ( .A(n404), .B(n403), .ZN(n661) );
  NOR2_X2 U525 ( .A1(n757), .A2(n575), .ZN(n404) );
  NOR2_X1 U526 ( .A1(n648), .A2(n524), .ZN(n526) );
  NAND2_X1 U527 ( .A1(n360), .A2(n430), .ZN(n406) );
  NAND2_X1 U528 ( .A1(n666), .A2(n510), .ZN(n414) );
  XNOR2_X2 U529 ( .A(n735), .B(KEYINPUT6), .ZN(n628) );
  NAND2_X1 U530 ( .A1(n701), .A2(G469), .ZN(n432) );
  XNOR2_X2 U531 ( .A(n417), .B(KEYINPUT0), .ZN(n599) );
  NOR2_X2 U532 ( .A1(n597), .A2(n596), .ZN(n417) );
  XNOR2_X2 U533 ( .A(n557), .B(KEYINPUT19), .ZN(n597) );
  AND2_X2 U534 ( .A1(n546), .A2(n744), .ZN(n557) );
  XNOR2_X2 U535 ( .A(n418), .B(G104), .ZN(n518) );
  XNOR2_X2 U536 ( .A(G122), .B(G113), .ZN(n418) );
  INV_X1 U537 ( .A(n420), .ZN(n622) );
  XNOR2_X1 U538 ( .A(n537), .B(n507), .ZN(n666) );
  XNOR2_X1 U539 ( .A(n526), .B(n444), .ZN(n546) );
  NAND2_X1 U540 ( .A1(n430), .A2(n427), .ZN(n555) );
  NOR2_X1 U541 ( .A1(n427), .A2(n426), .ZN(n425) );
  NAND2_X1 U542 ( .A1(n581), .A2(n433), .ZN(n657) );
  XNOR2_X1 U543 ( .A(n437), .B(n436), .ZN(n435) );
  NAND2_X1 U544 ( .A1(n585), .A2(n586), .ZN(n437) );
  NAND2_X1 U545 ( .A1(n439), .A2(n438), .ZN(n631) );
  NAND2_X1 U546 ( .A1(n656), .A2(n742), .ZN(n438) );
  INV_X1 U547 ( .A(n599), .ZN(n623) );
  NAND2_X1 U548 ( .A1(n599), .A2(n440), .ZN(n618) );
  INV_X1 U549 ( .A(n617), .ZN(n440) );
  XNOR2_X2 U550 ( .A(G119), .B(G110), .ZN(n516) );
  AND2_X1 U551 ( .A1(n659), .A2(n657), .ZN(n441) );
  AND2_X1 U552 ( .A1(n598), .A2(n731), .ZN(n442) );
  XOR2_X1 U553 ( .A(n583), .B(KEYINPUT64), .Z(n443) );
  NAND2_X1 U554 ( .A1(n527), .A2(G210), .ZN(n444) );
  INV_X1 U555 ( .A(KEYINPUT88), .ZN(n640) );
  BUF_X1 U556 ( .A(n671), .Z(n674) );
  XNOR2_X1 U557 ( .A(n371), .B(n471), .ZN(n472) );
  INV_X1 U558 ( .A(KEYINPUT90), .ZN(n592) );
  XNOR2_X1 U559 ( .A(n480), .B(n479), .ZN(n691) );
  XNOR2_X1 U560 ( .A(n513), .B(KEYINPUT10), .ZN(n474) );
  XNOR2_X1 U561 ( .A(n474), .B(n533), .ZN(n676) );
  NAND2_X1 U562 ( .A1(n770), .A2(G234), .ZN(n445) );
  XNOR2_X1 U563 ( .A(n445), .B(KEYINPUT8), .ZN(n489) );
  INV_X1 U564 ( .A(G221), .ZN(n465) );
  OR2_X1 U565 ( .A1(n489), .A2(n465), .ZN(n450) );
  XNOR2_X1 U566 ( .A(n446), .B(KEYINPUT74), .ZN(n449) );
  XNOR2_X1 U567 ( .A(n516), .B(n447), .ZN(n448) );
  NAND2_X1 U568 ( .A1(n686), .A2(n410), .ZN(n458) );
  XNOR2_X2 U569 ( .A(KEYINPUT15), .B(G902), .ZN(n641) );
  NAND2_X1 U570 ( .A1(n641), .A2(G234), .ZN(n452) );
  XNOR2_X1 U571 ( .A(n452), .B(KEYINPUT20), .ZN(n464) );
  NAND2_X1 U572 ( .A1(n464), .A2(G217), .ZN(n456) );
  XNOR2_X1 U573 ( .A(KEYINPUT83), .B(KEYINPUT100), .ZN(n454) );
  XNOR2_X1 U574 ( .A(KEYINPUT25), .B(KEYINPUT82), .ZN(n453) );
  XNOR2_X1 U575 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U576 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U577 ( .A(n459), .B(KEYINPUT14), .ZN(n462) );
  NAND2_X1 U578 ( .A1(G902), .A2(n462), .ZN(n460) );
  XOR2_X1 U579 ( .A(KEYINPUT98), .B(n460), .Z(n461) );
  NAND2_X1 U580 ( .A1(G953), .A2(n461), .ZN(n593) );
  OR2_X1 U581 ( .A1(n593), .A2(G900), .ZN(n463) );
  NAND2_X1 U582 ( .A1(G952), .A2(n462), .ZN(n755) );
  OR2_X1 U583 ( .A1(n755), .A2(G953), .ZN(n594) );
  NAND2_X1 U584 ( .A1(n463), .A2(n594), .ZN(n542) );
  INV_X1 U585 ( .A(n464), .ZN(n466) );
  OR2_X1 U586 ( .A1(n466), .A2(n465), .ZN(n468) );
  INV_X1 U587 ( .A(KEYINPUT21), .ZN(n467) );
  XNOR2_X1 U588 ( .A(n468), .B(n467), .ZN(n731) );
  NAND2_X1 U589 ( .A1(n542), .A2(n731), .ZN(n469) );
  NAND2_X1 U590 ( .A1(G214), .A2(n502), .ZN(n473) );
  XNOR2_X1 U591 ( .A(n473), .B(n472), .ZN(n480) );
  XNOR2_X1 U592 ( .A(n474), .B(n518), .ZN(n478) );
  XOR2_X1 U593 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n476) );
  XNOR2_X1 U594 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n475) );
  XNOR2_X1 U595 ( .A(n476), .B(n475), .ZN(n477) );
  NOR2_X1 U596 ( .A1(G902), .A2(n691), .ZN(n484) );
  XNOR2_X1 U597 ( .A(KEYINPUT107), .B(KEYINPUT13), .ZN(n482) );
  INV_X1 U598 ( .A(G475), .ZN(n481) );
  XNOR2_X1 U599 ( .A(n497), .B(n520), .ZN(n487) );
  XNOR2_X1 U600 ( .A(n485), .B(KEYINPUT7), .ZN(n486) );
  XNOR2_X1 U601 ( .A(n487), .B(n486), .ZN(n493) );
  INV_X1 U602 ( .A(G217), .ZN(n488) );
  OR2_X1 U603 ( .A1(n489), .A2(n488), .ZN(n491) );
  XOR2_X1 U604 ( .A(KEYINPUT9), .B(KEYINPUT108), .Z(n490) );
  XNOR2_X1 U605 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U606 ( .A(n493), .B(n492), .ZN(n688) );
  NAND2_X1 U607 ( .A1(n688), .A2(n410), .ZN(n495) );
  INV_X1 U608 ( .A(G478), .ZN(n494) );
  XNOR2_X1 U609 ( .A(n495), .B(n494), .ZN(n571) );
  NAND2_X1 U610 ( .A1(n570), .A2(n571), .ZN(n718) );
  XOR2_X1 U611 ( .A(KEYINPUT5), .B(KEYINPUT102), .Z(n500) );
  XNOR2_X1 U612 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U613 ( .A(n501), .B(n519), .ZN(n506) );
  NAND2_X1 U614 ( .A1(n502), .A2(G210), .ZN(n504) );
  XNOR2_X1 U615 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U616 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U617 ( .A(G472), .B(KEYINPUT103), .Z(n509) );
  INV_X1 U618 ( .A(KEYINPUT75), .ZN(n508) );
  XNOR2_X1 U619 ( .A(n509), .B(n508), .ZN(n510) );
  OR2_X1 U620 ( .A1(n718), .A2(n628), .ZN(n511) );
  NOR2_X1 U621 ( .A1(n551), .A2(n511), .ZN(n587) );
  XNOR2_X1 U622 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n512) );
  NAND2_X1 U623 ( .A1(n770), .A2(G224), .ZN(n514) );
  XNOR2_X1 U624 ( .A(KEYINPUT77), .B(KEYINPUT16), .ZN(n515) );
  XNOR2_X1 U625 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U626 ( .A(n518), .B(n517), .ZN(n522) );
  XNOR2_X1 U627 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U628 ( .A(n522), .B(n521), .ZN(n769) );
  XNOR2_X1 U629 ( .A(n523), .B(n769), .ZN(n648) );
  INV_X1 U630 ( .A(n641), .ZN(n524) );
  NAND2_X1 U631 ( .A1(n410), .A2(n525), .ZN(n527) );
  NAND2_X1 U632 ( .A1(n527), .A2(G214), .ZN(n744) );
  NAND2_X1 U633 ( .A1(n587), .A2(n376), .ZN(n529) );
  INV_X1 U634 ( .A(KEYINPUT36), .ZN(n528) );
  XNOR2_X1 U635 ( .A(n529), .B(n528), .ZN(n538) );
  XNOR2_X1 U636 ( .A(n531), .B(n530), .ZN(n535) );
  NAND2_X1 U637 ( .A1(n770), .A2(G227), .ZN(n532) );
  XNOR2_X1 U638 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U639 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U640 ( .A(n728), .B(KEYINPUT96), .ZN(n603) );
  NAND2_X1 U641 ( .A1(n538), .A2(n603), .ZN(n539) );
  XNOR2_X1 U642 ( .A(n539), .B(KEYINPUT115), .ZN(n776) );
  NAND2_X1 U643 ( .A1(n540), .A2(n731), .ZN(n610) );
  INV_X1 U644 ( .A(KEYINPUT110), .ZN(n541) );
  NAND2_X1 U645 ( .A1(n735), .A2(n744), .ZN(n544) );
  XNOR2_X1 U646 ( .A(KEYINPUT111), .B(KEYINPUT30), .ZN(n543) );
  XNOR2_X1 U647 ( .A(n544), .B(n543), .ZN(n576) );
  INV_X1 U648 ( .A(n571), .ZN(n545) );
  NAND2_X1 U649 ( .A1(n570), .A2(n545), .ZN(n611) );
  INV_X1 U650 ( .A(n590), .ZN(n547) );
  NOR2_X1 U651 ( .A1(n611), .A2(n547), .ZN(n548) );
  AND2_X1 U652 ( .A1(n576), .A2(n548), .ZN(n549) );
  NAND2_X1 U653 ( .A1(n578), .A2(n549), .ZN(n714) );
  OR2_X1 U654 ( .A1(n570), .A2(n571), .ZN(n722) );
  NAND2_X1 U655 ( .A1(n722), .A2(n718), .ZN(n626) );
  INV_X1 U656 ( .A(n626), .ZN(n742) );
  NAND2_X1 U657 ( .A1(KEYINPUT47), .A2(n742), .ZN(n550) );
  XOR2_X1 U658 ( .A(KEYINPUT87), .B(n550), .Z(n561) );
  INV_X1 U659 ( .A(n551), .ZN(n552) );
  NAND2_X1 U660 ( .A1(n552), .A2(n735), .ZN(n554) );
  XOR2_X1 U661 ( .A(KEYINPUT112), .B(KEYINPUT28), .Z(n553) );
  XNOR2_X1 U662 ( .A(n554), .B(n553), .ZN(n556) );
  BUF_X1 U663 ( .A(n597), .Z(n558) );
  INV_X1 U664 ( .A(n558), .ZN(n559) );
  NAND2_X1 U665 ( .A1(n574), .A2(n559), .ZN(n710) );
  NAND2_X1 U666 ( .A1(n710), .A2(KEYINPUT47), .ZN(n560) );
  AND2_X1 U667 ( .A1(n561), .A2(n560), .ZN(n562) );
  AND2_X1 U668 ( .A1(n714), .A2(n562), .ZN(n567) );
  INV_X1 U669 ( .A(KEYINPUT47), .ZN(n563) );
  NAND2_X1 U670 ( .A1(n626), .A2(n563), .ZN(n564) );
  OR2_X1 U671 ( .A1(n710), .A2(n564), .ZN(n565) );
  XNOR2_X1 U672 ( .A(n565), .B(KEYINPUT78), .ZN(n566) );
  NAND2_X1 U673 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U674 ( .A1(n776), .A2(n568), .ZN(n586) );
  XNOR2_X1 U675 ( .A(KEYINPUT79), .B(KEYINPUT38), .ZN(n569) );
  INV_X1 U676 ( .A(n570), .ZN(n572) );
  NAND2_X1 U677 ( .A1(n572), .A2(n571), .ZN(n746) );
  INV_X1 U678 ( .A(KEYINPUT114), .ZN(n573) );
  INV_X1 U679 ( .A(n574), .ZN(n575) );
  AND2_X1 U680 ( .A1(n576), .A2(n745), .ZN(n577) );
  NAND2_X1 U681 ( .A1(n578), .A2(n577), .ZN(n579) );
  INV_X1 U682 ( .A(n718), .ZN(n580) );
  XNOR2_X1 U683 ( .A(KEYINPUT92), .B(KEYINPUT46), .ZN(n583) );
  XNOR2_X1 U684 ( .A(n584), .B(n443), .ZN(n585) );
  NAND2_X1 U685 ( .A1(n587), .A2(n744), .ZN(n588) );
  NOR2_X1 U686 ( .A1(n588), .A2(n399), .ZN(n589) );
  XNOR2_X1 U687 ( .A(n589), .B(KEYINPUT43), .ZN(n591) );
  OR2_X1 U688 ( .A1(n591), .A2(n590), .ZN(n659) );
  OR2_X1 U689 ( .A1(n593), .A2(G898), .ZN(n595) );
  AND2_X1 U690 ( .A1(n595), .A2(n594), .ZN(n596) );
  INV_X1 U691 ( .A(n746), .ZN(n598) );
  NAND2_X1 U692 ( .A1(n599), .A2(n442), .ZN(n601) );
  XNOR2_X1 U693 ( .A(KEYINPUT76), .B(KEYINPUT22), .ZN(n600) );
  XNOR2_X1 U694 ( .A(n601), .B(n600), .ZN(n630) );
  XNOR2_X1 U695 ( .A(n628), .B(KEYINPUT86), .ZN(n602) );
  INV_X1 U696 ( .A(n732), .ZN(n627) );
  NAND2_X1 U697 ( .A1(n603), .A2(n627), .ZN(n604) );
  XNOR2_X1 U698 ( .A(n604), .B(KEYINPUT109), .ZN(n605) );
  XNOR2_X1 U699 ( .A(KEYINPUT85), .B(KEYINPUT32), .ZN(n606) );
  OR2_X1 U700 ( .A1(n735), .A2(n732), .ZN(n607) );
  NOR2_X1 U701 ( .A1(n399), .A2(n607), .ZN(n608) );
  AND2_X1 U702 ( .A1(n609), .A2(n608), .ZN(n658) );
  INV_X1 U703 ( .A(n610), .ZN(n727) );
  INV_X1 U704 ( .A(n611), .ZN(n612) );
  NAND2_X1 U705 ( .A1(n613), .A2(n612), .ZN(n616) );
  INV_X1 U706 ( .A(KEYINPUT91), .ZN(n614) );
  NAND2_X1 U707 ( .A1(n636), .A2(KEYINPUT44), .ZN(n632) );
  XNOR2_X1 U708 ( .A(n618), .B(KEYINPUT101), .ZN(n620) );
  INV_X1 U709 ( .A(n735), .ZN(n619) );
  NAND2_X1 U710 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U711 ( .A1(n622), .A2(n735), .ZN(n738) );
  INV_X1 U712 ( .A(KEYINPUT31), .ZN(n624) );
  NOR2_X1 U713 ( .A1(n399), .A2(n627), .ZN(n629) );
  NAND2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n634) );
  XNOR2_X1 U715 ( .A(n634), .B(n633), .ZN(n635) );
  OR2_X2 U716 ( .A1(n665), .A2(KEYINPUT44), .ZN(n637) );
  INV_X1 U717 ( .A(n638), .ZN(n639) );
  XNOR2_X1 U718 ( .A(n641), .B(KEYINPUT89), .ZN(n642) );
  NAND2_X1 U719 ( .A1(n642), .A2(KEYINPUT2), .ZN(n643) );
  XOR2_X1 U720 ( .A(KEYINPUT67), .B(n643), .Z(n644) );
  INV_X1 U721 ( .A(KEYINPUT2), .ZN(n725) );
  INV_X1 U722 ( .A(KEYINPUT66), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n698), .A2(G210), .ZN(n653) );
  BUF_X1 U724 ( .A(n648), .Z(n649) );
  XNOR2_X1 U725 ( .A(KEYINPUT95), .B(KEYINPUT54), .ZN(n650) );
  XOR2_X1 U726 ( .A(n650), .B(KEYINPUT55), .Z(n651) );
  XNOR2_X1 U727 ( .A(n653), .B(n652), .ZN(n655) );
  INV_X1 U728 ( .A(G952), .ZN(n654) );
  NAND2_X1 U729 ( .A1(n654), .A2(G953), .ZN(n694) );
  XNOR2_X1 U730 ( .A(n656), .B(G101), .ZN(G3) );
  XNOR2_X1 U731 ( .A(n657), .B(G134), .ZN(G36) );
  XOR2_X1 U732 ( .A(G110), .B(n658), .Z(G12) );
  XNOR2_X1 U733 ( .A(n659), .B(G140), .ZN(G42) );
  NOR2_X1 U734 ( .A1(n706), .A2(n718), .ZN(n660) );
  XOR2_X1 U735 ( .A(G104), .B(n660), .Z(G6) );
  XNOR2_X1 U736 ( .A(n661), .B(G137), .ZN(G39) );
  XOR2_X1 U737 ( .A(G119), .B(KEYINPUT126), .Z(n662) );
  XNOR2_X1 U738 ( .A(n663), .B(n662), .ZN(G21) );
  XOR2_X1 U739 ( .A(G131), .B(KEYINPUT127), .Z(n664) );
  XOR2_X1 U740 ( .A(n665), .B(G122), .Z(G24) );
  NAND2_X1 U741 ( .A1(n698), .A2(G472), .ZN(n668) );
  XNOR2_X1 U742 ( .A(n668), .B(n667), .ZN(n669) );
  NAND2_X1 U743 ( .A1(n669), .A2(n694), .ZN(n670) );
  XNOR2_X1 U744 ( .A(n670), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U745 ( .A(n672), .B(KEYINPUT124), .Z(n673) );
  XNOR2_X1 U746 ( .A(n674), .B(n673), .ZN(n675) );
  XOR2_X1 U747 ( .A(n676), .B(n675), .Z(n680) );
  XNOR2_X1 U748 ( .A(n680), .B(KEYINPUT125), .ZN(n677) );
  XNOR2_X1 U749 ( .A(n678), .B(n677), .ZN(n679) );
  NAND2_X1 U750 ( .A1(n679), .A2(n770), .ZN(n684) );
  XNOR2_X1 U751 ( .A(n680), .B(G227), .ZN(n681) );
  NAND2_X1 U752 ( .A1(n681), .A2(G900), .ZN(n682) );
  NAND2_X1 U753 ( .A1(n682), .A2(G953), .ZN(n683) );
  NAND2_X1 U754 ( .A1(n684), .A2(n683), .ZN(G72) );
  NAND2_X1 U755 ( .A1(n372), .A2(G217), .ZN(n685) );
  XOR2_X1 U756 ( .A(n685), .B(n686), .Z(n687) );
  INV_X1 U757 ( .A(n694), .ZN(n704) );
  NOR2_X1 U758 ( .A1(n687), .A2(n704), .ZN(G66) );
  NOR2_X1 U759 ( .A1(n689), .A2(n704), .ZN(G63) );
  NAND2_X1 U760 ( .A1(n698), .A2(G475), .ZN(n693) );
  XOR2_X1 U761 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n690) );
  XNOR2_X1 U762 ( .A(n693), .B(n692), .ZN(n695) );
  NAND2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n697) );
  XOR2_X1 U764 ( .A(KEYINPUT68), .B(KEYINPUT60), .Z(n696) );
  XNOR2_X1 U765 ( .A(n697), .B(n696), .ZN(G60) );
  NAND2_X1 U766 ( .A1(n372), .A2(G469), .ZN(n703) );
  XOR2_X1 U767 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n699) );
  XNOR2_X1 U768 ( .A(n699), .B(KEYINPUT58), .ZN(n700) );
  XNOR2_X1 U769 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U770 ( .A(n703), .B(n702), .ZN(n705) );
  NOR2_X1 U771 ( .A1(n705), .A2(n704), .ZN(G54) );
  NOR2_X1 U772 ( .A1(n706), .A2(n722), .ZN(n708) );
  XNOR2_X1 U773 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n707) );
  XNOR2_X1 U774 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U775 ( .A(G107), .B(n709), .ZN(G9) );
  XOR2_X1 U776 ( .A(KEYINPUT29), .B(KEYINPUT116), .Z(n712) );
  INV_X1 U777 ( .A(n710), .ZN(n716) );
  NAND2_X1 U778 ( .A1(n716), .A2(n433), .ZN(n711) );
  XNOR2_X1 U779 ( .A(n712), .B(n711), .ZN(n713) );
  XOR2_X1 U780 ( .A(G143), .B(n714), .Z(n715) );
  XNOR2_X1 U781 ( .A(n715), .B(KEYINPUT117), .ZN(G45) );
  NAND2_X1 U782 ( .A1(n716), .A2(n580), .ZN(n717) );
  XNOR2_X1 U783 ( .A(n717), .B(G146), .ZN(G48) );
  NOR2_X1 U784 ( .A1(n718), .A2(n721), .ZN(n719) );
  XOR2_X1 U785 ( .A(KEYINPUT118), .B(n719), .Z(n720) );
  XNOR2_X1 U786 ( .A(G113), .B(n720), .ZN(G15) );
  NOR2_X1 U787 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U788 ( .A(G116), .B(n723), .Z(G18) );
  NAND2_X1 U789 ( .A1(n373), .A2(n725), .ZN(n726) );
  NOR2_X1 U790 ( .A1(n399), .A2(n727), .ZN(n729) );
  XNOR2_X1 U791 ( .A(n729), .B(KEYINPUT50), .ZN(n730) );
  XNOR2_X1 U792 ( .A(n730), .B(KEYINPUT119), .ZN(n737) );
  NOR2_X1 U793 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U794 ( .A(KEYINPUT49), .B(n733), .Z(n734) );
  NOR2_X1 U795 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U796 ( .A1(n737), .A2(n736), .ZN(n739) );
  NAND2_X1 U797 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U798 ( .A(KEYINPUT51), .B(n740), .ZN(n741) );
  NOR2_X1 U799 ( .A1(n741), .A2(n757), .ZN(n752) );
  NOR2_X1 U800 ( .A1(n743), .A2(n742), .ZN(n749) );
  NOR2_X1 U801 ( .A1(n745), .A2(n744), .ZN(n747) );
  NOR2_X1 U802 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U803 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U804 ( .A1(n397), .A2(n750), .ZN(n751) );
  NOR2_X1 U805 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U806 ( .A(n753), .B(KEYINPUT52), .ZN(n754) );
  NOR2_X1 U807 ( .A1(n755), .A2(n754), .ZN(n756) );
  OR2_X1 U808 ( .A1(n756), .A2(G953), .ZN(n760) );
  NOR2_X1 U809 ( .A1(n397), .A2(n757), .ZN(n759) );
  NOR2_X1 U810 ( .A1(n760), .A2(n759), .ZN(n761) );
  AND2_X1 U811 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U812 ( .A(KEYINPUT53), .B(n763), .ZN(G75) );
  NAND2_X1 U813 ( .A1(n374), .A2(n770), .ZN(n767) );
  NAND2_X1 U814 ( .A1(G953), .A2(G224), .ZN(n764) );
  XNOR2_X1 U815 ( .A(KEYINPUT61), .B(n764), .ZN(n765) );
  NAND2_X1 U816 ( .A1(n765), .A2(G898), .ZN(n766) );
  NAND2_X1 U817 ( .A1(n767), .A2(n766), .ZN(n774) );
  XNOR2_X1 U818 ( .A(G101), .B(KEYINPUT122), .ZN(n768) );
  XNOR2_X1 U819 ( .A(n769), .B(n768), .ZN(n772) );
  NOR2_X1 U820 ( .A1(n770), .A2(G898), .ZN(n771) );
  NOR2_X1 U821 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U822 ( .A(n774), .B(n773), .ZN(n775) );
  XOR2_X1 U823 ( .A(KEYINPUT123), .B(n775), .Z(G69) );
  XNOR2_X1 U824 ( .A(G125), .B(n776), .ZN(n777) );
  XNOR2_X1 U825 ( .A(n777), .B(KEYINPUT37), .ZN(G27) );
endmodule

