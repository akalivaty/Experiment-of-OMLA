//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n548, new_n550, new_n551, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n597,
    new_n599, new_n600, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1139, new_n1140;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT67), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n467), .A2(new_n473), .A3(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n464), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(G137), .A3(new_n464), .ZN(new_n478));
  INV_X1    g053(.A(G101), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n464), .A2(G2104), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n476), .A2(new_n481), .ZN(G160));
  AND2_X1   g057(.A1(new_n477), .A2(KEYINPUT68), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n477), .A2(KEYINPUT68), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n485), .A2(new_n464), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n464), .A2(G112), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n487), .B(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  XOR2_X1   g067(.A(new_n492), .B(KEYINPUT69), .Z(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  NAND3_X1  g069(.A1(new_n477), .A2(G126), .A3(G2105), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G114), .C2(new_n464), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n499), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n467), .A2(new_n473), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n502));
  OAI211_X1 g077(.A(G138), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n501), .A2(new_n502), .B1(KEYINPUT4), .B2(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n467), .A2(new_n473), .A3(KEYINPUT70), .A4(new_n500), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n498), .B1(new_n504), .B2(new_n505), .ZN(G164));
  OR2_X1    g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI21_X1  g093(.A(G543), .B1(new_n515), .B2(new_n516), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n512), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  XOR2_X1   g098(.A(KEYINPUT71), .B(KEYINPUT7), .Z(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n524), .B(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G89), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n517), .A2(new_n529), .B1(new_n519), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n528), .A2(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  AOI22_X1  g108(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n511), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  INV_X1    g111(.A(G52), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n517), .A2(new_n536), .B1(new_n519), .B2(new_n537), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n535), .A2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  AOI22_X1  g115(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n511), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n517), .A2(new_n543), .B1(new_n519), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT72), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  INV_X1    g127(.A(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(KEYINPUT6), .A2(G651), .ZN(new_n554));
  NAND2_X1  g129(.A1(KEYINPUT6), .A2(G651), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G53), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(new_n509), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n507), .A2(new_n508), .B1(new_n554), .B2(new_n555), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n562), .A2(G651), .B1(new_n563), .B2(G91), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n558), .A2(new_n564), .ZN(G299));
  NAND2_X1  g140(.A1(new_n563), .A2(G87), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n556), .A2(G49), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  INV_X1    g145(.A(G48), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n517), .A2(new_n570), .B1(new_n519), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g147(.A(G61), .B1(new_n514), .B2(new_n513), .ZN(new_n573));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n511), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G305));
  AOI22_X1  g152(.A1(new_n563), .A2(G85), .B1(new_n556), .B2(G47), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT73), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(new_n511), .ZN(new_n581));
  AND2_X1   g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n563), .A2(G92), .ZN(new_n585));
  XOR2_X1   g160(.A(new_n585), .B(KEYINPUT10), .Z(new_n586));
  NAND2_X1  g161(.A1(G79), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G66), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n560), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(G54), .B2(new_n556), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n584), .B1(new_n592), .B2(G868), .ZN(G321));
  XNOR2_X1  g168(.A(G321), .B(KEYINPUT74), .ZN(G284));
  MUX2_X1   g169(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g170(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g171(.A(G559), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n592), .B1(new_n597), .B2(G860), .ZN(G148));
  NAND2_X1  g173(.A1(new_n592), .A2(new_n597), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(G868), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g176(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g177(.A1(new_n467), .A2(new_n473), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(new_n480), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT12), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT13), .ZN(new_n606));
  INV_X1    g181(.A(G2100), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n486), .A2(G135), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n488), .A2(G123), .ZN(new_n611));
  OR2_X1    g186(.A1(G99), .A2(G2105), .ZN(new_n612));
  OAI211_X1 g187(.A(new_n612), .B(G2104), .C1(G111), .C2(new_n464), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(G2096), .Z(new_n615));
  NAND3_X1  g190(.A1(new_n608), .A2(new_n609), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT75), .ZN(G156));
  XNOR2_X1  g192(.A(G1341), .B(G1348), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT77), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n619), .B(new_n620), .Z(new_n621));
  INV_X1    g196(.A(KEYINPUT14), .ZN(new_n622));
  XNOR2_X1  g197(.A(G2427), .B(G2438), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2430), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(new_n625), .B2(new_n624), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n621), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(G2443), .B(G2446), .Z(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n628), .A2(new_n631), .ZN(new_n633));
  AND3_X1   g208(.A1(new_n632), .A2(G14), .A3(new_n633), .ZN(G401));
  XOR2_X1   g209(.A(G2072), .B(G2078), .Z(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT79), .B(KEYINPUT17), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2067), .B(G2678), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT78), .ZN(new_n639));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  NAND3_X1  g215(.A1(new_n637), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT80), .Z(new_n642));
  INV_X1    g217(.A(new_n640), .ZN(new_n643));
  NOR3_X1   g218(.A1(new_n639), .A2(new_n635), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT18), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n640), .B1(new_n639), .B2(new_n635), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n637), .B2(new_n639), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n642), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT81), .ZN(new_n649));
  XOR2_X1   g224(.A(G2096), .B(G2100), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(G227));
  XNOR2_X1  g226(.A(G1971), .B(G1976), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT19), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G1956), .B(G2474), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT82), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1961), .B(G1966), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n654), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT20), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n654), .B1(new_n656), .B2(new_n658), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n656), .A2(new_n658), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n660), .B(new_n663), .C1(new_n653), .C2(new_n662), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1991), .B(G1996), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G229));
  INV_X1    g245(.A(G29), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G35), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT94), .Z(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n493), .B2(G29), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT29), .ZN(new_n675));
  INV_X1    g250(.A(G2090), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G5), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(G171), .B2(new_n679), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n681), .A2(G1961), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT24), .ZN(new_n683));
  INV_X1    g258(.A(G34), .ZN(new_n684));
  AOI21_X1  g259(.A(G29), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(new_n683), .B2(new_n684), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(G160), .B2(new_n671), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT88), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n671), .A2(G32), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n488), .A2(G129), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT89), .Z(new_n691));
  NAND3_X1  g266(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT26), .Z(new_n693));
  INV_X1    g268(.A(G105), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(new_n694), .B2(new_n480), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n486), .B2(G141), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n689), .B1(new_n697), .B2(G29), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT27), .B(G1996), .ZN(new_n699));
  OAI221_X1 g274(.A(new_n682), .B1(new_n688), .B2(G2084), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(KEYINPUT92), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(KEYINPUT92), .ZN(new_n702));
  NAND4_X1  g277(.A1(new_n677), .A2(new_n678), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n679), .A2(G21), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G168), .B2(new_n679), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(G1966), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT90), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT30), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n709), .A2(G28), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n671), .B1(new_n709), .B2(G28), .ZN(new_n711));
  AND2_X1   g286(.A1(KEYINPUT31), .A2(G11), .ZN(new_n712));
  NOR2_X1   g287(.A1(KEYINPUT31), .A2(G11), .ZN(new_n713));
  OAI22_X1  g288(.A1(new_n710), .A2(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n706), .B2(G1966), .ZN(new_n715));
  INV_X1    g290(.A(new_n614), .ZN(new_n716));
  AOI22_X1  g291(.A1(G29), .A2(new_n716), .B1(new_n681), .B2(G1961), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n708), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(KEYINPUT91), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n671), .A2(G33), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT25), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n486), .B2(G139), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT86), .ZN(new_n724));
  INV_X1    g299(.A(new_n603), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n725), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n726), .A2(new_n464), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT87), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n720), .B1(new_n729), .B2(new_n671), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(G2072), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n719), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n671), .A2(G26), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT28), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n486), .A2(G140), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n488), .A2(G128), .ZN(new_n736));
  OR2_X1    g311(.A1(G104), .A2(G2105), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n737), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT85), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n735), .A2(new_n736), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n734), .B1(new_n740), .B2(G29), .ZN(new_n741));
  INV_X1    g316(.A(G2067), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G4), .A2(G16), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT84), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n591), .B2(new_n679), .ZN(new_n746));
  INV_X1    g321(.A(G1348), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n679), .A2(G19), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n546), .B2(new_n679), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G1341), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n679), .A2(G20), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT23), .Z(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G299), .B2(G16), .ZN(new_n754));
  INV_X1    g329(.A(G1956), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  OR3_X1    g331(.A1(new_n748), .A2(new_n751), .A3(new_n756), .ZN(new_n757));
  AOI211_X1 g332(.A(new_n743), .B(new_n757), .C1(new_n698), .C2(new_n699), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n732), .A2(new_n758), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n718), .A2(KEYINPUT91), .B1(G2084), .B2(new_n688), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n671), .A2(G27), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT93), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n501), .A2(new_n502), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n763), .A2(new_n505), .A3(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n498), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n762), .B1(new_n767), .B2(G29), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(G2078), .Z(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n730), .B2(G2072), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n760), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n759), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n704), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(KEYINPUT95), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT95), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n704), .A2(new_n772), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n679), .A2(G22), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G166), .B2(new_n679), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1971), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n679), .A2(G23), .ZN(new_n780));
  INV_X1    g355(.A(G288), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(new_n679), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT33), .B(G1976), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(G6), .A2(G16), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n576), .B2(G16), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT32), .B(G1981), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n779), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT34), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n679), .A2(G24), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n582), .B2(new_n679), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(G1986), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n671), .A2(G25), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n464), .A2(G107), .ZN(new_n797));
  OAI21_X1  g372(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n488), .A2(G119), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n486), .A2(G131), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n796), .B1(new_n803), .B2(new_n671), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT35), .B(G1991), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n792), .A2(new_n795), .A3(new_n806), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT83), .Z(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n791), .B2(new_n790), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(KEYINPUT36), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n809), .A2(KEYINPUT36), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n774), .A2(new_n776), .B1(new_n810), .B2(new_n811), .ZN(G311));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n810), .ZN(new_n813));
  INV_X1    g388(.A(new_n776), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n775), .B1(new_n704), .B2(new_n772), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(G150));
  NAND2_X1  g391(.A1(new_n592), .A2(G559), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT38), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(new_n511), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT96), .B(G93), .ZN(new_n821));
  INV_X1    g396(.A(G55), .ZN(new_n822));
  OAI22_X1  g397(.A1(new_n517), .A2(new_n821), .B1(new_n519), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n546), .B(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n818), .B(new_n825), .Z(new_n826));
  OR2_X1    g401(.A1(new_n826), .A2(KEYINPUT39), .ZN(new_n827));
  INV_X1    g402(.A(G860), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(KEYINPUT39), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n824), .A2(new_n828), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT37), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(G145));
  XNOR2_X1  g408(.A(new_n740), .B(new_n767), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n486), .A2(G142), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n488), .A2(G130), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n464), .A2(G118), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n835), .B(new_n836), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n834), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n729), .A2(new_n691), .A3(new_n696), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n724), .A2(new_n728), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n697), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n803), .A2(KEYINPUT97), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n803), .A2(KEYINPUT97), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n605), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n847), .A2(new_n605), .A3(new_n848), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n846), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n845), .B1(new_n851), .B2(new_n852), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n841), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n614), .B(G160), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n493), .B(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n846), .A2(new_n853), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n845), .A2(new_n851), .A3(new_n852), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n840), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n856), .A2(new_n858), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT98), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n856), .A2(new_n864), .A3(new_n858), .A4(new_n861), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n858), .B1(new_n856), .B2(new_n861), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n867), .A2(G37), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n866), .A2(KEYINPUT40), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT40), .B1(new_n866), .B2(new_n868), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(G395));
  XNOR2_X1  g446(.A(G303), .B(KEYINPUT99), .ZN(new_n872));
  XNOR2_X1  g447(.A(G290), .B(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n781), .B(new_n576), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(KEYINPUT42), .Z(new_n876));
  XNOR2_X1  g451(.A(new_n591), .B(G299), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(KEYINPUT41), .Z(new_n878));
  XOR2_X1   g453(.A(new_n599), .B(new_n825), .Z(new_n879));
  MUX2_X1   g454(.A(new_n877), .B(new_n878), .S(new_n879), .Z(new_n880));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n881), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n876), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n876), .A2(new_n883), .ZN(new_n885));
  OAI21_X1  g460(.A(G868), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(G868), .B2(new_n824), .ZN(G295));
  OAI21_X1  g462(.A(new_n886), .B1(G868), .B2(new_n824), .ZN(G331));
  XNOR2_X1  g463(.A(new_n825), .B(G301), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(G168), .ZN(new_n890));
  INV_X1    g465(.A(new_n877), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n878), .B2(new_n890), .ZN(new_n893));
  INV_X1    g468(.A(new_n875), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n892), .B(new_n875), .C1(new_n878), .C2(new_n890), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT43), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n895), .A2(new_n900), .A3(new_n896), .A4(new_n897), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(KEYINPUT44), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT101), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n899), .A2(new_n903), .A3(new_n901), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n898), .A2(KEYINPUT101), .A3(KEYINPUT43), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n902), .B1(new_n906), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g482(.A(KEYINPUT45), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(G164), .B2(G1384), .ZN(new_n909));
  INV_X1    g484(.A(G1384), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n767), .A2(KEYINPUT45), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(G40), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n476), .A2(new_n912), .A3(new_n481), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n909), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G1966), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(KEYINPUT110), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(G1384), .B1(new_n765), .B2(new_n766), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT50), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n920));
  INV_X1    g495(.A(G2084), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .A4(new_n913), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n916), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT110), .B1(new_n914), .B2(new_n915), .ZN(new_n924));
  OAI21_X1  g499(.A(G8), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT121), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g502(.A(KEYINPUT121), .B(G8), .C1(new_n923), .C2(new_n924), .ZN(new_n928));
  XOR2_X1   g503(.A(KEYINPUT106), .B(G8), .Z(new_n929));
  NOR2_X1   g504(.A1(G168), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n927), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n929), .ZN(new_n933));
  OAI211_X1 g508(.A(KEYINPUT122), .B(new_n933), .C1(new_n923), .C2(new_n924), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n930), .A2(KEYINPUT51), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n933), .B1(new_n923), .B2(new_n924), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT122), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n932), .A2(KEYINPUT51), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n930), .B1(new_n923), .B2(new_n924), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT62), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT62), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n936), .A2(new_n939), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT51), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n930), .B1(new_n925), .B2(new_n926), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n946), .B1(new_n947), .B2(new_n928), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n944), .B(new_n941), .C1(new_n945), .C2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT125), .ZN(new_n950));
  INV_X1    g525(.A(G8), .ZN(new_n951));
  XNOR2_X1  g526(.A(KEYINPUT103), .B(G1971), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n914), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(KEYINPUT104), .B(G2090), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n919), .A2(new_n920), .A3(new_n913), .A4(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n951), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(G303), .A2(G8), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n959), .B(KEYINPUT55), .Z(new_n960));
  NAND3_X1  g535(.A1(new_n953), .A2(new_n955), .A3(KEYINPUT105), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n958), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G1976), .ZN(new_n963));
  NOR2_X1   g538(.A1(G288), .A2(new_n963), .ZN(new_n964));
  AOI211_X1 g539(.A(new_n929), .B(new_n964), .C1(new_n917), .C2(new_n913), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT52), .B1(G288), .B2(new_n963), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT49), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT107), .ZN(new_n968));
  AOI22_X1  g543(.A1(new_n563), .A2(G86), .B1(new_n556), .B2(G48), .ZN(new_n969));
  INV_X1    g544(.A(new_n575), .ZN(new_n970));
  INV_X1    g545(.A(G1981), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(G1981), .B1(new_n572), .B2(new_n575), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n968), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n971), .B1(new_n969), .B2(new_n970), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n572), .A2(new_n575), .A3(G1981), .ZN(new_n976));
  OAI22_X1  g551(.A1(new_n975), .A2(new_n976), .B1(KEYINPUT107), .B2(new_n967), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n974), .B1(new_n977), .B2(new_n968), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n929), .B1(new_n917), .B2(new_n913), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n965), .A2(new_n966), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n767), .A2(new_n913), .A3(new_n910), .ZN(new_n981));
  INV_X1    g556(.A(new_n964), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n981), .A2(new_n933), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT52), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT109), .B1(new_n980), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n979), .A2(new_n982), .A3(new_n966), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n978), .A2(new_n979), .ZN(new_n987));
  AND4_X1   g562(.A1(KEYINPUT109), .A2(new_n984), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n929), .B1(new_n953), .B2(new_n955), .ZN(new_n989));
  OAI22_X1  g564(.A1(new_n985), .A2(new_n988), .B1(new_n960), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n950), .B1(new_n962), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n958), .A2(new_n960), .A3(new_n961), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n989), .A2(new_n960), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n987), .A2(new_n986), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n983), .A2(KEYINPUT52), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n980), .A2(KEYINPUT109), .A3(new_n984), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n992), .A2(KEYINPUT125), .A3(new_n993), .A4(new_n999), .ZN(new_n1000));
  XOR2_X1   g575(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n914), .B2(G2078), .ZN(new_n1002));
  INV_X1    g577(.A(G1961), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n913), .B1(new_n917), .B2(new_n918), .ZN(new_n1004));
  NOR3_X1   g579(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n1008));
  OR3_X1    g583(.A1(new_n914), .A2(new_n1008), .A3(G2078), .ZN(new_n1009));
  AOI21_X1  g584(.A(G301), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n991), .A2(new_n1000), .A3(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n943), .A2(new_n949), .A3(new_n1011), .ZN(new_n1012));
  AOI211_X1 g587(.A(G1976), .B(G288), .C1(new_n978), .C2(new_n979), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n976), .B(KEYINPUT108), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n979), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n995), .A2(new_n996), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1015), .B1(new_n992), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n992), .A2(new_n993), .A3(new_n999), .ZN(new_n1020));
  OAI211_X1 g595(.A(G168), .B(new_n933), .C1(new_n923), .C2(new_n924), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1019), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n990), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1021), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1023), .A2(KEYINPUT111), .A3(new_n992), .A4(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT63), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1022), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n962), .A2(new_n1026), .A3(new_n1017), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n958), .A2(new_n961), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1028), .B(new_n1024), .C1(new_n960), .C2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1018), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n474), .A2(new_n475), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n464), .B1(new_n1033), .B2(KEYINPUT124), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(KEYINPUT124), .B2(new_n1033), .ZN(new_n1035));
  NOR4_X1   g610(.A1(new_n481), .A2(new_n1008), .A3(new_n912), .A4(G2078), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n909), .A2(new_n911), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1002), .A2(new_n1006), .A3(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(G171), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1032), .B1(new_n1010), .B2(new_n1039), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n991), .A2(new_n1000), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(G301), .B1(new_n1038), .B2(KEYINPUT126), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(KEYINPUT126), .B2(new_n1038), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1009), .A2(new_n1006), .A3(new_n1002), .A4(G301), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1044), .A2(KEYINPUT54), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT127), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT127), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1043), .A2(new_n1048), .A3(new_n1045), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n755), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1052), .A2(KEYINPUT112), .ZN(new_n1053));
  NAND2_X1  g628(.A1(G299), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(KEYINPUT112), .ZN(new_n1055));
  XOR2_X1   g630(.A(new_n1055), .B(KEYINPUT113), .Z(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(G299), .A2(new_n1053), .A3(new_n1056), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT56), .B(G2072), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n909), .A2(new_n911), .A3(new_n913), .A4(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1051), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1060), .B1(new_n1051), .B2(new_n1062), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(new_n1064), .B2(KEYINPUT118), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1051), .A2(new_n1066), .A3(new_n1060), .A4(new_n1062), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1065), .A2(KEYINPUT61), .A3(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n592), .A2(KEYINPUT119), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n1071));
  AND4_X1   g646(.A1(new_n1071), .A2(new_n767), .A3(new_n913), .A4(new_n910), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1071), .B1(new_n917), .B2(new_n913), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n742), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n747), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT60), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n592), .B2(KEYINPUT119), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1070), .A2(new_n1074), .A3(new_n1075), .A4(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1069), .B1(new_n1079), .B2(new_n1076), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g657(.A(KEYINPUT117), .B(KEYINPUT61), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1063), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1083), .B1(new_n1084), .B2(new_n1064), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT116), .B1(new_n1086), .B2(KEYINPUT115), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n981), .A2(KEYINPUT114), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n917), .A2(new_n1071), .A3(new_n913), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT58), .B(G1341), .Z(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G1996), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n909), .A2(new_n911), .A3(new_n1092), .A4(new_n913), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1087), .B1(new_n1094), .B2(new_n546), .ZN(new_n1095));
  INV_X1    g670(.A(new_n546), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1087), .B1(KEYINPUT116), .B2(new_n1086), .ZN(new_n1097));
  AOI211_X1 g672(.A(new_n1096), .B(new_n1097), .C1(new_n1091), .C2(new_n1093), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1068), .A2(new_n1082), .A3(new_n1085), .A4(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n591), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1063), .B1(new_n1102), .B2(new_n1064), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1100), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1101), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1041), .B(new_n1050), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n940), .A2(new_n942), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1012), .B(new_n1031), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n909), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n913), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n697), .B(G1996), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n740), .B(new_n742), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n802), .B(new_n805), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1110), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1110), .ZN(new_n1117));
  NOR2_X1   g692(.A1(G290), .A2(G1986), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT102), .ZN(new_n1120));
  NAND2_X1  g695(.A1(G290), .A2(G1986), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1120), .B(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1116), .B1(new_n1117), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1108), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1119), .A2(new_n1110), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1125), .A2(KEYINPUT48), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1125), .A2(KEYINPUT48), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1116), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1117), .A2(new_n1092), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1129), .B(KEYINPUT46), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1117), .B1(new_n1113), .B2(new_n697), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(new_n1132), .B(KEYINPUT47), .Z(new_n1133));
  NAND3_X1  g708(.A1(new_n1114), .A2(new_n805), .A3(new_n803), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(G2067), .B2(new_n740), .ZN(new_n1135));
  AOI211_X1 g710(.A(new_n1128), .B(new_n1133), .C1(new_n1117), .C2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1124), .A2(new_n1136), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g712(.A1(new_n866), .A2(new_n868), .ZN(new_n1139));
  NOR4_X1   g713(.A1(G229), .A2(new_n462), .A3(G401), .A4(G227), .ZN(new_n1140));
  AND4_X1   g714(.A1(new_n1139), .A2(new_n905), .A3(new_n904), .A4(new_n1140), .ZN(G308));
  NAND4_X1  g715(.A1(new_n1139), .A2(new_n905), .A3(new_n904), .A4(new_n1140), .ZN(G225));
endmodule


