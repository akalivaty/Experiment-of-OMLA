//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n628, new_n629, new_n630, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G104), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(KEYINPUT3), .A3(G104), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n191), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G101), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n193), .A2(G107), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT88), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n200), .B1(new_n190), .B2(G104), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n193), .A2(KEYINPUT88), .A3(G107), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n199), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n198), .B1(new_n197), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT89), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT1), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n207), .B1(new_n206), .B2(KEYINPUT1), .ZN(new_n210));
  OAI21_X1  g024(.A(G128), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n206), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT1), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n206), .A2(new_n213), .A3(new_n216), .A4(G128), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n204), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT64), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(new_n205), .A3(G143), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT64), .B1(new_n212), .B2(G146), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n212), .A2(G146), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(G128), .B1(new_n222), .B2(new_n216), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n217), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT10), .ZN(new_n227));
  OAI22_X1  g041(.A1(new_n218), .A2(KEYINPUT10), .B1(new_n204), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT87), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n194), .A2(new_n195), .ZN(new_n230));
  OAI21_X1  g044(.A(G101), .B1(new_n230), .B2(new_n191), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n231), .A2(KEYINPUT86), .A3(KEYINPUT4), .A4(new_n198), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT86), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT4), .B1(new_n196), .B2(new_n197), .ZN(new_n234));
  AOI211_X1 g048(.A(G101), .B(new_n191), .C1(new_n194), .C2(new_n195), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  OR3_X1    g051(.A1(new_n196), .A2(KEYINPUT4), .A3(new_n197), .ZN(new_n238));
  AND2_X1   g052(.A1(KEYINPUT0), .A2(G128), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n206), .A2(new_n213), .A3(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(KEYINPUT0), .A2(G128), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT65), .B1(new_n223), .B2(new_n242), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n223), .A2(KEYINPUT65), .A3(new_n242), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n238), .B(new_n240), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n229), .B1(new_n237), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n245), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n232), .A2(new_n236), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(KEYINPUT87), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n228), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G137), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT11), .B1(new_n251), .B2(G134), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(G134), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT66), .ZN(new_n255));
  INV_X1    g069(.A(G131), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n251), .A2(KEYINPUT11), .A3(G134), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n254), .A2(new_n255), .A3(new_n256), .A4(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT11), .ZN(new_n259));
  INV_X1    g073(.A(G134), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n259), .B1(new_n260), .B2(G137), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(G137), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n261), .A2(new_n257), .A3(new_n256), .A4(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT66), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n254), .A2(new_n257), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n258), .A2(new_n264), .B1(new_n265), .B2(G131), .ZN(new_n266));
  OR2_X1    g080(.A1(new_n250), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n228), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n237), .A2(new_n229), .A3(new_n245), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT87), .B1(new_n247), .B2(new_n248), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n268), .B(new_n266), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(G110), .B(G140), .ZN(new_n273));
  INV_X1    g087(.A(G227), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(G953), .ZN(new_n275));
  XOR2_X1   g089(.A(new_n273), .B(new_n275), .Z(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n218), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n204), .A2(new_n225), .A3(new_n217), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n266), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n281), .B(KEYINPUT12), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n277), .B1(new_n250), .B2(new_n266), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n282), .B1(new_n283), .B2(KEYINPUT90), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n271), .A2(new_n276), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT90), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n284), .A2(new_n287), .A3(KEYINPUT91), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT91), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT12), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n281), .B(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n291), .B1(new_n285), .B2(new_n286), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n283), .A2(KEYINPUT90), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n289), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n278), .B1(new_n288), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G469), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n267), .A2(new_n283), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n282), .A2(new_n271), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n299), .B1(new_n300), .B2(new_n276), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n297), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G469), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n189), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(G113), .B(G122), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n305), .B(new_n193), .ZN(new_n306));
  INV_X1    g120(.A(G140), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(G125), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(KEYINPUT78), .ZN(new_n309));
  INV_X1    g123(.A(G125), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(G140), .ZN(new_n311));
  OR2_X1    g125(.A1(new_n311), .A2(KEYINPUT77), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(KEYINPUT77), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n309), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT16), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n311), .A2(KEYINPUT16), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n315), .A2(new_n205), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n205), .B1(new_n315), .B2(new_n316), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G237), .ZN(new_n320));
  INV_X1    g134(.A(G953), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G214), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(G143), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(new_n256), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n256), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT17), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n324), .A2(KEYINPUT17), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n319), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n314), .A2(G146), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT95), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n311), .A2(new_n308), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(KEYINPUT81), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n205), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n314), .A2(KEYINPUT95), .A3(G146), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n334), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(KEYINPUT18), .A2(G131), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n324), .A2(KEYINPUT18), .B1(new_n323), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n306), .B1(new_n331), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT20), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n315), .A2(new_n316), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G146), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n325), .A2(new_n326), .ZN(new_n348));
  MUX2_X1   g162(.A(new_n336), .B(new_n314), .S(KEYINPUT19), .Z(new_n349));
  OAI211_X1 g163(.A(new_n347), .B(new_n348), .C1(G146), .C2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n306), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n351), .A3(new_n342), .ZN(new_n352));
  NOR2_X1   g166(.A1(G475), .A2(G902), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n344), .A2(new_n345), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n319), .A2(new_n330), .B1(new_n339), .B2(new_n341), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n352), .B(new_n353), .C1(new_n355), .C2(new_n351), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT20), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n306), .A2(KEYINPUT96), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n297), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n355), .A2(new_n359), .ZN(new_n362));
  OAI21_X1  g176(.A(G475), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G128), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G143), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT13), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n212), .A2(G128), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(KEYINPUT97), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT13), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n369), .B1(new_n370), .B2(new_n368), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT97), .B1(new_n367), .B2(new_n368), .ZN(new_n372));
  OAI21_X1  g186(.A(G134), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n368), .A2(new_n366), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n260), .ZN(new_n375));
  INV_X1    g189(.A(G116), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(G122), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(G122), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n190), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n190), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n373), .B(new_n375), .C1(new_n380), .C2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n374), .B(new_n260), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n379), .B1(new_n377), .B2(KEYINPUT14), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(KEYINPUT14), .B2(new_n379), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G107), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n387), .A3(new_n381), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G217), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n187), .A2(new_n390), .A3(G953), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n383), .A2(new_n388), .A3(new_n391), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n297), .ZN(new_n396));
  INV_X1    g210(.A(G478), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n397), .A2(KEYINPUT15), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n396), .B(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n364), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(G234), .A2(G237), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n401), .A2(G952), .A3(new_n321), .ZN(new_n402));
  XOR2_X1   g216(.A(KEYINPUT21), .B(G898), .Z(new_n403));
  XNOR2_X1  g217(.A(new_n403), .B(KEYINPUT98), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n401), .A2(G902), .A3(G953), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n402), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  XOR2_X1   g221(.A(new_n407), .B(KEYINPUT99), .Z(new_n408));
  NAND2_X1  g222(.A1(new_n400), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(G214), .B1(G237), .B2(G902), .ZN(new_n411));
  XOR2_X1   g225(.A(new_n411), .B(KEYINPUT92), .Z(new_n412));
  XOR2_X1   g226(.A(KEYINPUT2), .B(G113), .Z(new_n413));
  XNOR2_X1  g227(.A(G116), .B(G119), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n413), .B(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n238), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n416), .B1(new_n236), .B2(new_n232), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n414), .A2(KEYINPUT5), .ZN(new_n418));
  INV_X1    g232(.A(G119), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G116), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n418), .B(G113), .C1(KEYINPUT5), .C2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n413), .A2(new_n414), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(new_n204), .ZN(new_n424));
  XNOR2_X1  g238(.A(G110), .B(G122), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  OR3_X1    g240(.A1(new_n417), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n426), .B1(new_n417), .B2(new_n424), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(KEYINPUT6), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT6), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n430), .B(new_n426), .C1(new_n417), .C2(new_n424), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT65), .ZN(new_n432));
  NOR3_X1   g246(.A1(new_n212), .A2(KEYINPUT64), .A3(G146), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n219), .B1(new_n205), .B2(G143), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n433), .B1(new_n206), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n242), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n432), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n223), .A2(KEYINPUT65), .A3(new_n242), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(G125), .A3(new_n240), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n226), .A2(new_n310), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G224), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(G953), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n442), .B(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n429), .A2(new_n431), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n442), .ZN(new_n448));
  AND2_X1   g262(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n449));
  NOR2_X1   g263(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n445), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n423), .B(new_n204), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n425), .B(KEYINPUT8), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n448), .A2(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n444), .B1(new_n440), .B2(new_n441), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n455), .A2(KEYINPUT94), .A3(KEYINPUT7), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT94), .B1(new_n455), .B2(KEYINPUT7), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n454), .B(new_n427), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n447), .A2(new_n297), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(G210), .B1(G237), .B2(G902), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n447), .A2(new_n458), .A3(new_n297), .A4(new_n460), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n412), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n304), .A2(new_n410), .A3(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(G472), .A2(G902), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT67), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n258), .A2(new_n264), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n260), .A2(G137), .ZN(new_n469));
  OAI21_X1  g283(.A(G131), .B1(new_n469), .B2(new_n253), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n226), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT30), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n240), .B1(new_n244), .B2(new_n243), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n471), .B(new_n472), .C1(new_n473), .C2(new_n266), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n265), .A2(G131), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n263), .A2(KEYINPUT66), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n263), .A2(KEYINPUT66), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(new_n439), .A3(new_n240), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n472), .B1(new_n480), .B2(new_n471), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n467), .B(new_n415), .C1(new_n475), .C2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n320), .A2(new_n321), .A3(G210), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n483), .B(KEYINPUT27), .Z(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(KEYINPUT68), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT26), .B(G101), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n485), .B(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n415), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n471), .B1(new_n473), .B2(new_n266), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT30), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n488), .B1(new_n490), .B2(new_n474), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n471), .B(new_n488), .C1(new_n473), .C2(new_n266), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(KEYINPUT67), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n482), .B(new_n487), .C1(new_n491), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT31), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n475), .A2(new_n481), .ZN(new_n497));
  OAI22_X1  g311(.A1(new_n497), .A2(new_n488), .B1(KEYINPUT67), .B2(new_n493), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT31), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n498), .A2(new_n499), .A3(new_n482), .A4(new_n487), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n488), .B1(new_n480), .B2(new_n471), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n502), .B1(new_n493), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT28), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n492), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n487), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  AND4_X1   g322(.A1(KEYINPUT70), .A2(new_n496), .A3(new_n500), .A4(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n507), .B1(new_n495), .B2(KEYINPUT31), .ZN(new_n510));
  AOI21_X1  g324(.A(KEYINPUT70), .B1(new_n510), .B2(new_n500), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n466), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT32), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(KEYINPUT71), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT71), .ZN(new_n515));
  INV_X1    g329(.A(new_n466), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n496), .A2(new_n500), .A3(new_n508), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT70), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n510), .A2(KEYINPUT70), .A3(new_n500), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n515), .B1(new_n521), .B2(KEYINPUT32), .ZN(new_n522));
  OAI211_X1 g336(.A(KEYINPUT32), .B(new_n466), .C1(new_n509), .C2(new_n511), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n514), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G472), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n498), .A2(new_n482), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT29), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n487), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT72), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n493), .A2(new_n503), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n530), .B1(new_n531), .B2(new_n505), .ZN(new_n532));
  OAI211_X1 g346(.A(KEYINPUT72), .B(KEYINPUT28), .C1(new_n493), .C2(new_n503), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n506), .B(KEYINPUT73), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n528), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AND4_X1   g350(.A1(new_n528), .A2(new_n504), .A3(new_n487), .A4(new_n506), .ZN(new_n537));
  OR3_X1    g351(.A1(new_n529), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n526), .B1(new_n538), .B2(new_n297), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n525), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n365), .A2(KEYINPUT23), .A3(G119), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT75), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n542), .A2(new_n543), .B1(new_n419), .B2(G128), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n365), .A2(G119), .ZN(new_n545));
  AND2_X1   g359(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n546));
  NOR2_X1   g360(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n544), .B(new_n548), .C1(new_n543), .C2(new_n542), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(G110), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT79), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT24), .B(G110), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n419), .A2(G128), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n545), .A2(new_n553), .A3(KEYINPUT74), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT74), .B1(new_n545), .B2(new_n553), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n552), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n550), .B1(new_n551), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n557), .B1(new_n551), .B2(new_n556), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT80), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT80), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n557), .B(new_n560), .C1(new_n551), .C2(new_n556), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n559), .A2(new_n347), .A3(new_n561), .A4(new_n337), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n554), .A2(new_n555), .A3(new_n552), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(G110), .B2(new_n549), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n564), .B1(new_n317), .B2(new_n318), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n321), .A2(G221), .A3(G234), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT82), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT22), .B(G137), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n562), .A2(new_n565), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n570), .B1(new_n562), .B2(new_n565), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT84), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT25), .B1(new_n575), .B2(KEYINPUT83), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n574), .A2(new_n297), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n390), .B1(G234), .B2(new_n297), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n572), .A2(new_n573), .A3(G902), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n575), .A2(KEYINPUT25), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT83), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n581), .B1(new_n575), .B2(KEYINPUT25), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n577), .B(new_n578), .C1(new_n579), .C2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n578), .A2(G902), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(KEYINPUT85), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n574), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n465), .A2(new_n541), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G101), .ZN(G3));
  INV_X1    g405(.A(new_n304), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n297), .B1(new_n509), .B2(new_n511), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G472), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n512), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n592), .A2(new_n588), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n411), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n462), .B2(new_n463), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n408), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n396), .A2(G478), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n395), .B(KEYINPUT33), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n297), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n600), .B1(new_n602), .B2(G478), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n364), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n596), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT34), .B(G104), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G6));
  AND2_X1   g422(.A1(new_n358), .A2(new_n363), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n399), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n599), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n596), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT100), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT35), .B(G107), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G9));
  INV_X1    g429(.A(new_n595), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n562), .A2(new_n565), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n569), .A2(KEYINPUT36), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n586), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n584), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n465), .A2(new_n616), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT37), .B(G110), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT101), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n622), .B(new_n624), .ZN(G12));
  INV_X1    g439(.A(G900), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n402), .B1(new_n406), .B2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n610), .A2(new_n627), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n628), .A2(new_n621), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n541), .A2(new_n304), .A3(new_n598), .A4(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G128), .ZN(G30));
  XOR2_X1   g445(.A(new_n627), .B(KEYINPUT39), .Z(new_n632));
  NAND2_X1  g446(.A1(new_n304), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(new_n633), .B(KEYINPUT40), .Z(new_n634));
  OAI21_X1  g448(.A(new_n495), .B1(new_n487), .B2(new_n531), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n297), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G472), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n525), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n462), .A2(new_n463), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT38), .ZN(new_n640));
  INV_X1    g454(.A(new_n621), .ZN(new_n641));
  AND4_X1   g455(.A1(new_n364), .A2(new_n641), .A3(new_n399), .A4(new_n411), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n634), .A2(new_n638), .A3(new_n640), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G143), .ZN(G45));
  NOR2_X1   g458(.A1(new_n604), .A2(new_n627), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n541), .A2(new_n304), .A3(new_n598), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G146), .ZN(G48));
  OAI21_X1  g463(.A(KEYINPUT91), .B1(new_n284), .B2(new_n287), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n292), .A2(new_n289), .A3(new_n293), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n650), .A2(new_n651), .B1(new_n272), .B2(new_n277), .ZN(new_n652));
  OAI21_X1  g466(.A(G469), .B1(new_n652), .B2(G902), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n298), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n189), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n541), .A2(new_n589), .A3(new_n605), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT41), .B(G113), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G15));
  NAND4_X1  g472(.A1(new_n541), .A2(new_n589), .A3(new_n611), .A4(new_n655), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G116), .ZN(G18));
  NAND4_X1  g474(.A1(new_n653), .A2(new_n298), .A3(new_n188), .A4(new_n598), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n641), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n541), .A2(new_n662), .A3(new_n410), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G119), .ZN(G21));
  XOR2_X1   g478(.A(new_n466), .B(KEYINPUT102), .Z(new_n665));
  NAND2_X1  g479(.A1(new_n496), .A2(new_n500), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n487), .B1(new_n534), .B2(new_n535), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT103), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n589), .A2(new_n594), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n598), .A2(new_n364), .A3(new_n399), .ZN(new_n671));
  INV_X1    g485(.A(new_n408), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n673), .A2(new_n188), .A3(new_n298), .A4(new_n653), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(G122), .Z(G24));
  NAND3_X1  g490(.A1(new_n669), .A2(new_n594), .A3(new_n645), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n677), .A2(new_n661), .A3(new_n641), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(new_n310), .ZN(G27));
  NAND2_X1  g493(.A1(new_n512), .A2(new_n513), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n523), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n539), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n681), .A2(KEYINPUT105), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n588), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n462), .A2(new_n463), .A3(new_n411), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT104), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n690));
  NOR4_X1   g504(.A1(new_n592), .A2(new_n689), .A3(new_n690), .A4(new_n646), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n298), .A2(new_n303), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n692), .A2(new_n188), .A3(new_n688), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n541), .A2(new_n693), .A3(new_n589), .A4(new_n645), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n686), .A2(new_n691), .B1(new_n694), .B2(new_n690), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(new_n256), .ZN(G33));
  NAND4_X1  g510(.A1(new_n541), .A2(new_n693), .A3(new_n589), .A4(new_n628), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G134), .ZN(G36));
  NAND2_X1  g512(.A1(new_n609), .A2(new_n603), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n595), .A3(new_n621), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(KEYINPUT44), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n701), .A2(new_n704), .A3(new_n595), .A4(new_n621), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n689), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n301), .A2(KEYINPUT45), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n301), .A2(KEYINPUT45), .ZN(new_n708));
  OAI21_X1  g522(.A(G469), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n296), .A2(new_n297), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n709), .A2(KEYINPUT46), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n298), .B1(new_n712), .B2(KEYINPUT106), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n301), .B(KEYINPUT45), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n710), .B1(new_n715), .B2(G469), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n714), .B1(new_n716), .B2(KEYINPUT46), .ZN(new_n717));
  OAI21_X1  g531(.A(KEYINPUT107), .B1(new_n713), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n716), .A2(new_n714), .A3(KEYINPUT46), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n712), .A2(KEYINPUT106), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n719), .A2(new_n720), .A3(new_n721), .A4(new_n298), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n716), .A2(KEYINPUT46), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n718), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n706), .A2(new_n724), .A3(new_n188), .A4(new_n632), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G137), .ZN(G39));
  NOR4_X1   g540(.A1(new_n541), .A2(new_n589), .A3(new_n646), .A4(new_n689), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n724), .A2(KEYINPUT47), .A3(new_n188), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT47), .B1(new_n724), .B2(new_n188), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G140), .ZN(G42));
  OR4_X1    g545(.A1(new_n588), .A2(new_n189), .A3(new_n412), .A4(new_n699), .ZN(new_n732));
  AOI211_X1 g546(.A(new_n640), .B(new_n732), .C1(KEYINPUT49), .C2(new_n654), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n654), .A2(KEYINPUT49), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(KEYINPUT108), .ZN(new_n735));
  INV_X1    g549(.A(new_n638), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n733), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n640), .A2(new_n411), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n655), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT113), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n701), .A2(new_n402), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n670), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n655), .A2(new_n688), .ZN(new_n747));
  INV_X1    g561(.A(new_n402), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n747), .A2(new_n588), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n603), .A2(new_n364), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n736), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n747), .A2(new_n742), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n669), .A2(new_n621), .A3(new_n594), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n755), .A2(KEYINPUT51), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n654), .A2(new_n188), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n728), .A2(new_n729), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n743), .A2(new_n688), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n746), .B(new_n756), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(G952), .ZN(new_n761));
  INV_X1    g575(.A(new_n661), .ZN(new_n762));
  AOI211_X1 g576(.A(new_n761), .B(G953), .C1(new_n743), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n749), .A2(new_n736), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n763), .B1(new_n764), .B2(new_n604), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n686), .A2(new_n752), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n766), .A2(KEYINPUT48), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(KEYINPUT48), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n765), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n760), .A2(new_n769), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n758), .A2(new_n759), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n746), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n744), .B(KEYINPUT50), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT114), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n771), .A2(new_n773), .A3(new_n775), .A4(new_n755), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n770), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n680), .A2(new_n515), .A3(new_n523), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n539), .B1(new_n779), .B2(new_n514), .ZN(new_n780));
  INV_X1    g594(.A(new_n598), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n780), .A2(new_n592), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n678), .B1(new_n782), .B2(new_n629), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n621), .A2(new_n627), .A3(new_n671), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n638), .A2(new_n304), .A3(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n783), .A2(KEYINPUT52), .A3(new_n648), .A4(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n678), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n630), .A2(new_n648), .A3(new_n787), .A4(new_n785), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n627), .ZN(new_n792));
  AND4_X1   g606(.A1(new_n400), .A2(new_n688), .A3(new_n621), .A4(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n541), .A2(new_n793), .A3(new_n304), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n693), .A2(new_n645), .A3(new_n753), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n697), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT110), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n697), .A2(new_n794), .A3(KEYINPUT110), .A4(new_n795), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n695), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n801));
  INV_X1    g615(.A(new_n675), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n656), .A2(new_n659), .A3(new_n802), .A4(new_n663), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n464), .A2(new_n408), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n804), .A2(new_n610), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT109), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n804), .A2(new_n610), .A3(KEYINPUT109), .ZN(new_n808));
  OAI22_X1  g622(.A1(new_n807), .A2(new_n808), .B1(new_n604), .B2(new_n804), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n596), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n590), .A3(new_n622), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n803), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n791), .A2(new_n800), .A3(new_n801), .A4(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n788), .A2(new_n789), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n788), .A2(new_n789), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT111), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT111), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n786), .A2(new_n790), .A3(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n816), .A2(new_n818), .A3(new_n812), .A4(new_n800), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  OAI211_X1 g634(.A(KEYINPUT54), .B(new_n813), .C1(new_n820), .C2(new_n801), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT112), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n803), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n780), .A2(new_n409), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n675), .B1(new_n824), .B2(new_n662), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n825), .A2(KEYINPUT112), .A3(new_n656), .A4(new_n659), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n811), .A2(new_n801), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n791), .A2(new_n800), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n819), .B2(new_n801), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n778), .A2(new_n821), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n834));
  OAI22_X1  g648(.A1(new_n833), .A2(new_n834), .B1(G952), .B2(G953), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n737), .B1(new_n835), .B2(new_n836), .ZN(G75));
  NOR2_X1   g651(.A1(new_n830), .A2(new_n297), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(G210), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT56), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n429), .A2(new_n431), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(new_n446), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT55), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n839), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n843), .B1(new_n839), .B2(new_n840), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n761), .A2(G953), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT116), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n844), .A2(new_n845), .A3(new_n848), .ZN(G51));
  XNOR2_X1  g663(.A(new_n830), .B(KEYINPUT54), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n710), .B(KEYINPUT57), .Z(new_n851));
  OAI21_X1  g665(.A(new_n295), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n838), .A2(G469), .A3(new_n715), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n848), .B1(new_n852), .B2(new_n853), .ZN(G54));
  NAND2_X1  g668(.A1(KEYINPUT58), .A2(G475), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT117), .Z(new_n856));
  NAND2_X1  g670(.A1(new_n838), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n344), .A2(new_n352), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n847), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n858), .B2(new_n857), .ZN(G60));
  XNOR2_X1  g674(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n861));
  NAND2_X1  g675(.A1(G478), .A2(G902), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n861), .B(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n601), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n847), .B1(new_n850), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n832), .A2(new_n821), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n601), .B1(new_n866), .B2(new_n863), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n865), .A2(new_n867), .ZN(G63));
  NAND2_X1  g682(.A1(G217), .A2(G902), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n869), .B(KEYINPUT60), .Z(new_n870));
  NAND2_X1  g684(.A1(new_n798), .A2(new_n799), .ZN(new_n871));
  INV_X1    g685(.A(new_n695), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n872), .A3(new_n812), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n817), .B1(new_n786), .B2(new_n790), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT53), .B1(new_n875), .B2(new_n818), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n870), .B1(new_n876), .B2(new_n829), .ZN(new_n877));
  INV_X1    g691(.A(new_n574), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n848), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g693(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT119), .ZN(new_n881));
  INV_X1    g695(.A(new_n870), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n819), .A2(new_n801), .ZN(new_n883));
  INV_X1    g697(.A(new_n829), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n881), .B1(new_n885), .B2(new_n619), .ZN(new_n886));
  INV_X1    g700(.A(new_n619), .ZN(new_n887));
  NOR4_X1   g701(.A1(new_n830), .A2(KEYINPUT119), .A3(new_n887), .A4(new_n882), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n879), .B(new_n880), .C1(new_n886), .C2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n619), .B(new_n870), .C1(new_n876), .C2(new_n829), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT119), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n883), .A2(new_n884), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n893), .A2(new_n881), .A3(new_n619), .A4(new_n870), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n880), .B1(new_n895), .B2(new_n879), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n890), .A2(new_n896), .ZN(G66));
  OAI21_X1  g711(.A(G953), .B1(new_n405), .B2(new_n443), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n898), .B1(new_n812), .B2(G953), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n841), .B1(G898), .B2(new_n321), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n899), .B(new_n900), .ZN(G69));
  XOR2_X1   g715(.A(new_n497), .B(new_n349), .Z(new_n902));
  AND3_X1   g716(.A1(new_n630), .A2(new_n648), .A3(new_n787), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n643), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT62), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n610), .A2(new_n604), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n688), .A2(new_n906), .ZN(new_n907));
  OR4_X1    g721(.A1(new_n588), .A2(new_n780), .A3(new_n633), .A4(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n730), .A2(new_n725), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n902), .B1(new_n910), .B2(G953), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n321), .A2(G900), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n725), .A2(new_n903), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n913), .B(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n872), .A2(new_n697), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n872), .A2(KEYINPUT125), .A3(new_n697), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI211_X1 g734(.A(new_n588), .B(new_n671), .C1(new_n684), .C2(new_n685), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n921), .A2(new_n724), .A3(new_n188), .A4(new_n632), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n730), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n915), .A2(new_n920), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n912), .B1(new_n924), .B2(new_n321), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n911), .B1(new_n925), .B2(new_n902), .ZN(new_n926));
  OAI21_X1  g740(.A(G953), .B1(new_n274), .B2(new_n626), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT122), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n926), .A2(KEYINPUT126), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT126), .B1(new_n926), .B2(new_n929), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n928), .B(KEYINPUT123), .Z(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n911), .B2(KEYINPUT121), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(KEYINPUT121), .B2(new_n911), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n925), .A2(new_n902), .ZN(new_n935));
  OAI22_X1  g749(.A1(new_n930), .A2(new_n931), .B1(new_n934), .B2(new_n935), .ZN(G72));
  NAND2_X1  g750(.A1(new_n910), .A2(new_n812), .ZN(new_n937));
  XNOR2_X1  g751(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n526), .A2(new_n297), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n938), .B(new_n939), .Z(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n487), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n527), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n848), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n527), .A2(new_n943), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n946), .A2(new_n944), .A3(new_n940), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n813), .B(new_n947), .C1(new_n820), .C2(new_n801), .ZN(new_n948));
  INV_X1    g762(.A(new_n812), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n941), .B1(new_n924), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n946), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n945), .A2(new_n948), .A3(new_n951), .ZN(G57));
endmodule


