//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT64), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT64), .A2(G146), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(G143), .A3(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n192), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT64), .A2(G146), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT64), .A2(G146), .ZN(new_n199));
  OAI211_X1 g013(.A(KEYINPUT65), .B(new_n193), .C1(new_n198), .C2(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(G143), .B1(new_n190), .B2(new_n191), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n202), .B1(new_n193), .B2(G146), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n200), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n195), .B1(new_n192), .B2(KEYINPUT1), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n197), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT68), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT68), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n208), .B(new_n197), .C1(new_n204), .C2(new_n205), .ZN(new_n209));
  XNOR2_X1  g023(.A(G104), .B(G107), .ZN(new_n210));
  INV_X1    g024(.A(G101), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT76), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G104), .ZN(new_n214));
  INV_X1    g028(.A(G104), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G107), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT76), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(G101), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT3), .B1(new_n215), .B2(G107), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(new_n213), .A3(G104), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n220), .A2(new_n222), .A3(new_n211), .A4(new_n216), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n212), .A2(new_n219), .A3(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n207), .A2(KEYINPUT10), .A3(new_n209), .A4(new_n224), .ZN(new_n225));
  XOR2_X1   g039(.A(KEYINPUT0), .B(G128), .Z(new_n226));
  OAI211_X1 g040(.A(new_n200), .B(new_n226), .C1(new_n201), .C2(new_n203), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n192), .A2(KEYINPUT0), .A3(G128), .A4(new_n194), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n220), .A2(new_n222), .A3(new_n216), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G101), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT75), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT75), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(new_n235), .A3(G101), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n234), .A2(KEYINPUT4), .A3(new_n223), .A4(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n227), .A2(KEYINPUT66), .A3(new_n228), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT4), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n232), .A2(new_n239), .A3(G101), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n231), .A2(new_n237), .A3(new_n238), .A4(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT1), .B1(new_n193), .B2(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT77), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT77), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n244), .B(KEYINPUT1), .C1(new_n193), .C2(G146), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n243), .A2(G128), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n192), .A2(new_n194), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n197), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n224), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT10), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT11), .ZN(new_n253));
  INV_X1    g067(.A(G134), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n253), .B1(new_n254), .B2(G137), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(G137), .ZN(new_n256));
  INV_X1    g070(.A(G137), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT11), .A3(G134), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G131), .ZN(new_n260));
  INV_X1    g074(.A(G131), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n255), .A2(new_n258), .A3(new_n261), .A4(new_n256), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n260), .A2(KEYINPUT67), .A3(new_n262), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n225), .A2(new_n241), .A3(new_n252), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT78), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT10), .B1(new_n249), .B2(new_n224), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n227), .A2(KEYINPUT66), .A3(new_n228), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT66), .B1(new_n227), .B2(new_n228), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n240), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n232), .A2(new_n235), .A3(G101), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n223), .A2(KEYINPUT4), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n275), .B1(new_n278), .B2(new_n234), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n271), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT78), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n280), .A2(new_n281), .A3(new_n268), .A4(new_n225), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n270), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(G110), .B(G140), .ZN(new_n284));
  INV_X1    g098(.A(G953), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n285), .A2(G227), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n284), .B(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n280), .A2(new_n225), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n267), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n283), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n206), .A2(new_n224), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n212), .A2(new_n219), .A3(new_n223), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n293), .B1(new_n197), .B2(new_n248), .ZN(new_n294));
  OAI211_X1 g108(.A(KEYINPUT12), .B(new_n263), .C1(new_n292), .C2(new_n294), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n293), .B(new_n197), .C1(new_n204), .C2(new_n205), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n250), .A2(new_n296), .B1(new_n266), .B2(new_n265), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n297), .A2(KEYINPUT79), .A3(KEYINPUT12), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT79), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n267), .B1(new_n292), .B2(new_n294), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT12), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n295), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n288), .B1(new_n283), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n187), .B1(new_n291), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G469), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT80), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT80), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n305), .A2(new_n308), .A3(G469), .ZN(new_n309));
  XOR2_X1   g123(.A(KEYINPUT81), .B(G469), .Z(new_n310));
  NAND3_X1  g124(.A1(new_n283), .A2(new_n303), .A3(new_n288), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n288), .B1(new_n283), .B2(new_n290), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT82), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AOI211_X1 g128(.A(KEYINPUT82), .B(new_n288), .C1(new_n283), .C2(new_n290), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n187), .B(new_n310), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n307), .A2(new_n309), .A3(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(G214), .B1(G237), .B2(G902), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G140), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G125), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT16), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G140), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n321), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n324), .A2(KEYINPUT73), .A3(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n323), .B1(new_n329), .B2(new_n322), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G146), .ZN(new_n331));
  NOR2_X1   g145(.A1(G237), .A2(G953), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(G143), .A3(G214), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(G143), .B1(new_n332), .B2(G214), .ZN(new_n335));
  OAI21_X1  g149(.A(G131), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n335), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(new_n261), .A3(new_n333), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT17), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n189), .B(new_n323), .C1(new_n329), .C2(new_n322), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n337), .A2(new_n333), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(KEYINPUT17), .A3(G131), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n331), .A2(new_n340), .A3(new_n341), .A4(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(G113), .B(G122), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(new_n215), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(KEYINPUT18), .A3(G131), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n321), .A2(new_n325), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n198), .A2(new_n199), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(new_n329), .B2(new_n189), .ZN(new_n351));
  NAND2_X1  g165(.A1(KEYINPUT18), .A2(G131), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n337), .A2(new_n333), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n347), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n344), .A2(new_n346), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n336), .A2(new_n338), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT19), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n327), .B2(new_n328), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n348), .A2(KEYINPUT19), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n349), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n331), .A2(new_n356), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n346), .B1(new_n361), .B2(new_n354), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n355), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(G475), .A2(G902), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT20), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n344), .A2(new_n346), .A3(new_n354), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n361), .A2(new_n354), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n367), .B1(new_n368), .B2(new_n346), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT20), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(new_n364), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n346), .B1(new_n344), .B2(new_n354), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n187), .B1(new_n355), .B2(new_n372), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n366), .A2(new_n371), .B1(G475), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n285), .A2(G952), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n375), .B1(G234), .B2(G237), .ZN(new_n376));
  NAND2_X1  g190(.A1(G234), .A2(G237), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n377), .A2(G902), .A3(G953), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT21), .B(G898), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT72), .B(G217), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT9), .B(G234), .ZN(new_n383));
  NOR3_X1   g197(.A1(new_n382), .A2(new_n383), .A3(G953), .ZN(new_n384));
  INV_X1    g198(.A(G122), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G116), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n213), .B1(new_n386), .B2(KEYINPUT14), .ZN(new_n387));
  XNOR2_X1  g201(.A(G116), .B(G122), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n387), .B(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n193), .A2(G128), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n195), .A2(G143), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT88), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT88), .B1(new_n390), .B2(new_n391), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n393), .A2(new_n254), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n390), .A2(new_n391), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT88), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(G134), .B1(new_n398), .B2(new_n392), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n389), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT89), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n254), .B1(new_n393), .B2(new_n394), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n398), .A2(G134), .A3(new_n392), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(KEYINPUT89), .A3(new_n389), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G116), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G122), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n386), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT87), .B(G107), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n410), .B(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n193), .A2(G128), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n195), .A2(G143), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n413), .B1(KEYINPUT13), .B2(new_n414), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n414), .A2(KEYINPUT13), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n254), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR3_X1   g231(.A1(new_n412), .A2(new_n417), .A3(new_n399), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n384), .B1(new_n407), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n384), .ZN(new_n421));
  AOI211_X1 g235(.A(new_n421), .B(new_n418), .C1(new_n402), .C2(new_n406), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n187), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT15), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(G478), .ZN(new_n425));
  INV_X1    g239(.A(G478), .ZN(new_n426));
  OAI221_X1 g240(.A(new_n187), .B1(KEYINPUT15), .B2(new_n426), .C1(new_n420), .C2(new_n422), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n374), .A2(new_n381), .A3(new_n425), .A4(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G210), .B1(G237), .B2(G902), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT86), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n206), .A2(new_n324), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n227), .A2(G125), .A3(new_n228), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n285), .A2(G224), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(KEYINPUT85), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n435), .A2(new_n438), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G119), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G116), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n408), .A2(G119), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G113), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT2), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT2), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G113), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n447), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n449), .A2(new_n451), .ZN(new_n453));
  XNOR2_X1  g267(.A(G116), .B(G119), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n240), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n445), .A2(KEYINPUT5), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(new_n448), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n454), .A2(KEYINPUT5), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n460), .A2(new_n461), .B1(new_n454), .B2(new_n453), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n237), .A2(new_n458), .B1(new_n224), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G110), .B(G122), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n463), .A2(KEYINPUT6), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT83), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n463), .B2(new_n464), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n468), .B1(new_n463), .B2(new_n464), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n224), .A2(new_n462), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n235), .B1(new_n232), .B2(G101), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n276), .A2(new_n471), .A3(new_n277), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n470), .B1(new_n472), .B2(new_n457), .ZN(new_n473));
  INV_X1    g287(.A(new_n464), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(KEYINPUT83), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n467), .A2(new_n469), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT84), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT84), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n467), .A2(new_n469), .A3(new_n478), .A4(new_n475), .ZN(new_n479));
  AOI211_X1 g293(.A(new_n443), .B(new_n465), .C1(new_n477), .C2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT7), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n436), .B1(new_n481), .B2(new_n439), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n463), .A2(new_n464), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n462), .B(new_n293), .ZN(new_n484));
  XOR2_X1   g298(.A(new_n464), .B(KEYINPUT8), .Z(new_n485));
  OAI211_X1 g299(.A(new_n482), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n441), .A2(new_n481), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n187), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n432), .B1(new_n480), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n477), .A2(new_n479), .ZN(new_n490));
  INV_X1    g304(.A(new_n465), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n442), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n488), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n493), .A3(new_n431), .ZN(new_n494));
  AOI211_X1 g308(.A(new_n319), .B(new_n428), .C1(new_n489), .C2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(G221), .B1(new_n383), .B2(G902), .ZN(new_n496));
  XOR2_X1   g310(.A(new_n496), .B(KEYINPUT74), .Z(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n317), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT90), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n317), .A2(new_n495), .A3(KEYINPUT90), .A4(new_n498), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n382), .B1(G234), .B2(new_n187), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n331), .A2(new_n341), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT23), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n444), .B2(G128), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n195), .A2(KEYINPUT23), .A3(G119), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n508), .B(new_n509), .C1(G119), .C2(new_n195), .ZN(new_n510));
  XNOR2_X1  g324(.A(G119), .B(G128), .ZN(new_n511));
  XOR2_X1   g325(.A(KEYINPUT24), .B(G110), .Z(new_n512));
  AOI22_X1  g326(.A1(new_n510), .A2(G110), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  OAI22_X1  g328(.A1(new_n510), .A2(G110), .B1(new_n511), .B2(new_n512), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n331), .A2(new_n350), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT22), .B(G137), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n285), .A2(G221), .A3(G234), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n514), .A2(new_n516), .A3(new_n520), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(KEYINPUT25), .A3(new_n187), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(new_n187), .A3(new_n523), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT25), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n505), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n504), .A2(G902), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n332), .A2(G210), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(KEYINPUT27), .ZN(new_n536));
  XNOR2_X1  g350(.A(KEYINPUT26), .B(G101), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n267), .A2(new_n231), .A3(new_n238), .ZN(new_n540));
  INV_X1    g354(.A(new_n256), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n254), .A2(G137), .ZN(new_n542));
  OAI21_X1  g356(.A(G131), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n543), .A2(new_n262), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n207), .A2(new_n544), .A3(new_n209), .ZN(new_n545));
  INV_X1    g359(.A(new_n456), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n540), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT70), .B1(new_n547), .B2(KEYINPUT28), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n540), .A2(new_n545), .A3(new_n546), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT70), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT28), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n206), .A2(new_n544), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n229), .B1(new_n260), .B2(new_n262), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n456), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n551), .B1(new_n549), .B2(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n548), .B(new_n552), .C1(KEYINPUT69), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(KEYINPUT69), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n539), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n540), .A2(new_n545), .A3(KEYINPUT30), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT30), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(new_n553), .B2(new_n554), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(new_n456), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n564), .A2(new_n538), .A3(new_n549), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT31), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT31), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n564), .A2(new_n567), .A3(new_n538), .A4(new_n549), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n560), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(G472), .A2(G902), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT32), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT32), .ZN(new_n573));
  INV_X1    g387(.A(new_n571), .ZN(new_n574));
  AOI211_X1 g388(.A(new_n573), .B(new_n574), .C1(new_n560), .C2(new_n569), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n546), .B1(new_n540), .B2(new_n545), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT28), .B1(new_n547), .B2(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n538), .A2(KEYINPUT29), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n578), .A2(new_n548), .A3(new_n552), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT71), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n550), .B1(new_n549), .B2(new_n551), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT71), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n584), .A2(new_n585), .A3(new_n578), .A4(new_n579), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n549), .A2(new_n555), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT28), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT69), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n584), .A2(new_n591), .A3(new_n538), .A4(new_n558), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n564), .A2(new_n549), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT29), .B1(new_n593), .B2(new_n539), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n587), .A2(new_n595), .A3(new_n187), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G472), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n534), .B1(new_n576), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n503), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT91), .B(G101), .Z(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G3));
  INV_X1    g416(.A(KEYINPUT92), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n566), .A2(new_n568), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n584), .A2(new_n591), .A3(new_n558), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n604), .B1(new_n539), .B2(new_n605), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n603), .B(G472), .C1(new_n606), .C2(G902), .ZN(new_n607));
  INV_X1    g421(.A(G472), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n570), .B2(new_n187), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT92), .B1(new_n570), .B2(new_n571), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n607), .B(new_n533), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n305), .A2(new_n308), .A3(G469), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n308), .B1(new_n305), .B2(G469), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n497), .B1(new_n615), .B2(new_n316), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n612), .A2(KEYINPUT93), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT93), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n317), .A2(new_n498), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n618), .B1(new_n619), .B2(new_n611), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n429), .B1(new_n480), .B2(new_n488), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n492), .A2(new_n493), .A3(new_n430), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n622), .A2(new_n318), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n374), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT33), .B1(new_n420), .B2(new_n422), .ZN(new_n626));
  INV_X1    g440(.A(new_n406), .ZN(new_n627));
  AOI21_X1  g441(.A(KEYINPUT89), .B1(new_n405), .B2(new_n389), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n419), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n421), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT33), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n407), .A2(new_n419), .A3(new_n384), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n626), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT94), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n426), .A2(G902), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n634), .A2(new_n636), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n423), .ZN(new_n640));
  OAI21_X1  g454(.A(KEYINPUT94), .B1(new_n640), .B2(G478), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n625), .B(new_n637), .C1(new_n639), .C2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n624), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n380), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n621), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT95), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT34), .B(G104), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  NAND2_X1  g463(.A1(new_n492), .A2(new_n493), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n319), .B1(new_n650), .B2(new_n429), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n623), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n425), .A2(new_n427), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n374), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n652), .A2(new_n380), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n621), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT35), .B(G107), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G9));
  NOR2_X1   g472(.A1(new_n521), .A2(KEYINPUT36), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT96), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(new_n517), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n529), .B1(new_n530), .B2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n607), .B(new_n663), .C1(new_n609), .C2(new_n610), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n503), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT37), .B(G110), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  AOI21_X1  g481(.A(new_n662), .B1(new_n576), .B2(new_n597), .ZN(new_n668));
  INV_X1    g482(.A(new_n376), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT97), .B(G900), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n378), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n654), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n674), .A2(new_n318), .A3(new_n622), .A4(new_n623), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT98), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n651), .A2(KEYINPUT98), .A3(new_n623), .A4(new_n674), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n668), .A2(new_n616), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G128), .ZN(G30));
  XNOR2_X1  g495(.A(new_n672), .B(KEYINPUT39), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n616), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n683), .A2(KEYINPUT40), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(KEYINPUT40), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n547), .A2(new_n577), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n187), .B1(new_n686), .B2(new_n538), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n539), .B1(new_n564), .B2(new_n549), .ZN(new_n688));
  OAI21_X1  g502(.A(G472), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n663), .B1(new_n576), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n489), .A2(new_n494), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n489), .A2(new_n494), .A3(new_n692), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n374), .B1(new_n425), .B2(new_n427), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n696), .A2(new_n318), .A3(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n684), .A2(new_n685), .A3(new_n690), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G143), .ZN(G45));
  INV_X1    g514(.A(new_n644), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n668), .A2(new_n616), .A3(new_n701), .A4(new_n672), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT100), .B(G146), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G48));
  OAI21_X1  g518(.A(new_n187), .B1(new_n314), .B2(new_n315), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G469), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n496), .A3(new_n316), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT101), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT101), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n706), .A2(new_n709), .A3(new_n496), .A4(new_n316), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n598), .A2(new_n645), .A3(new_n708), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT41), .B(G113), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G15));
  NAND4_X1  g527(.A1(new_n598), .A2(new_n655), .A3(new_n708), .A4(new_n710), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  NAND4_X1  g529(.A1(new_n624), .A2(new_n496), .A3(new_n706), .A4(new_n316), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n428), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n668), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  OAI21_X1  g534(.A(G472), .B1(new_n606), .B2(G902), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n578), .A2(new_n548), .A3(new_n552), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT102), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n584), .A2(KEYINPUT102), .A3(new_n578), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n724), .A2(new_n725), .A3(new_n539), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n571), .B1(new_n726), .B2(new_n604), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n525), .A2(new_n528), .ZN(new_n728));
  OAI211_X1 g542(.A(KEYINPUT103), .B(new_n531), .C1(new_n728), .C2(new_n505), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n730), .B1(new_n529), .B2(new_n532), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n721), .A2(new_n727), .A3(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n651), .A2(new_n623), .A3(new_n697), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n380), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n708), .A2(new_n734), .A3(new_n736), .A4(new_n710), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NOR2_X1   g552(.A1(new_n642), .A2(new_n673), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n739), .A2(new_n721), .A3(new_n727), .A4(new_n663), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n716), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n324), .ZN(G27));
  INV_X1    g556(.A(new_n496), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n743), .B1(new_n316), .B2(new_n306), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n744), .A2(KEYINPUT104), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n489), .A2(new_n318), .A3(new_n494), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n746), .B1(new_n744), .B2(KEYINPUT104), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n598), .A2(new_n745), .A3(new_n739), .A4(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n574), .B1(new_n560), .B2(new_n569), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT32), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT105), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n572), .A2(KEYINPUT106), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT106), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n751), .A2(new_n755), .A3(KEYINPUT32), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n753), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT105), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n575), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n573), .B1(new_n606), .B2(new_n574), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n755), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n572), .A2(KEYINPUT106), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n759), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n757), .A2(new_n763), .A3(new_n597), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(KEYINPUT42), .A3(new_n732), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n744), .A2(KEYINPUT104), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT104), .ZN(new_n767));
  AOI211_X1 g581(.A(new_n767), .B(new_n743), .C1(new_n316), .C2(new_n306), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n766), .A2(new_n768), .A3(new_n746), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n739), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n750), .B1(new_n765), .B2(new_n770), .ZN(new_n771));
  XOR2_X1   g585(.A(KEYINPUT107), .B(G131), .Z(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(G33));
  NAND4_X1  g587(.A1(new_n598), .A2(new_n745), .A3(new_n674), .A4(new_n747), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT108), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n769), .A2(KEYINPUT108), .A3(new_n598), .A4(new_n674), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G134), .ZN(G36));
  OAI21_X1  g593(.A(new_n721), .B1(KEYINPUT92), .B2(new_n751), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n607), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n374), .B(new_n637), .C1(new_n639), .C2(new_n641), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT43), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n638), .B(KEYINPUT94), .C1(G478), .C2(new_n640), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT43), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(new_n785), .A3(new_n374), .A4(new_n637), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n783), .A2(new_n786), .A3(new_n663), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n781), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n746), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n781), .A2(new_n788), .A3(KEYINPUT44), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n797), .B1(new_n291), .B2(new_n304), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n283), .A2(new_n288), .A3(new_n290), .ZN(new_n799));
  OAI21_X1  g613(.A(KEYINPUT79), .B1(new_n297), .B2(KEYINPUT12), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n300), .A2(new_n299), .A3(new_n301), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n802), .A2(new_n295), .B1(new_n270), .B2(new_n282), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n799), .B(KEYINPUT45), .C1(new_n803), .C2(new_n288), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n798), .A2(G469), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(G469), .A2(G902), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT46), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n805), .A2(KEYINPUT46), .A3(new_n806), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n316), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n807), .B1(new_n809), .B2(KEYINPUT109), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT109), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n808), .A2(new_n811), .A3(new_n316), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n813), .A2(new_n496), .A3(new_n682), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n791), .A2(KEYINPUT110), .A3(new_n792), .A4(new_n793), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n796), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G137), .ZN(G39));
  NAND3_X1  g631(.A1(new_n813), .A2(KEYINPUT47), .A3(new_n496), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT47), .B1(new_n813), .B2(new_n496), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n792), .A2(new_n534), .A3(new_n739), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n597), .A2(new_n760), .A3(new_n752), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT111), .B1(new_n821), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n820), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n825), .B1(new_n827), .B2(new_n818), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT111), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G140), .ZN(G42));
  INV_X1    g646(.A(new_n741), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n735), .A2(new_n673), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n760), .A2(new_n752), .A3(new_n689), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n834), .A2(new_n662), .A3(new_n835), .A4(new_n744), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n702), .A2(new_n680), .A3(new_n833), .A4(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n823), .A2(new_n498), .A3(new_n317), .A4(new_n663), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n741), .B1(new_n840), .B2(new_n679), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(KEYINPUT115), .A3(new_n702), .A4(new_n836), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT52), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT52), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n839), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n691), .A2(new_n318), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n642), .A2(new_n654), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n848), .A2(new_n849), .A3(new_n380), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n617), .A2(new_n620), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n664), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n501), .B(new_n502), .C1(new_n598), .C2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n854), .B1(new_n851), .B2(new_n853), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n711), .A2(new_n714), .A3(new_n719), .A4(new_n737), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n746), .A2(new_n653), .A3(new_n625), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n668), .A2(new_n859), .A3(new_n616), .A4(new_n672), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n721), .A2(new_n727), .A3(new_n663), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n745), .A2(new_n747), .A3(new_n861), .A4(new_n739), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n771), .A2(new_n858), .A3(new_n778), .A4(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n857), .A2(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n847), .A2(new_n865), .A3(KEYINPUT53), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n846), .B1(new_n845), .B2(new_n837), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT53), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT54), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n855), .A2(new_n856), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n771), .A2(new_n858), .A3(new_n778), .A4(new_n863), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n839), .A2(new_n845), .A3(new_n842), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n845), .B1(new_n839), .B2(new_n842), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n870), .B(new_n871), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n865), .A2(KEYINPUT53), .A3(new_n867), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n835), .A2(new_n534), .A3(new_n669), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n707), .A2(new_n746), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(new_n643), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n375), .B(KEYINPUT118), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n783), .A2(new_n786), .A3(new_n376), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n733), .A2(new_n884), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n882), .B(new_n883), .C1(new_n716), .C2(new_n885), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n764), .A2(new_n732), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n707), .A2(new_n884), .A3(new_n746), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n889), .A2(KEYINPUT48), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(KEYINPUT48), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n886), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT50), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n318), .B1(new_n694), .B2(new_n695), .ZN(new_n894));
  INV_X1    g708(.A(new_n707), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n893), .B1(new_n896), .B2(new_n885), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n733), .A2(new_n884), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n898), .A2(KEYINPUT50), .A3(new_n895), .A4(new_n894), .ZN(new_n899));
  AOI22_X1  g713(.A1(new_n897), .A2(new_n899), .B1(new_n888), .B2(new_n861), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n625), .B1(new_n784), .B2(new_n637), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n880), .A2(new_n881), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT116), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n880), .A2(KEYINPUT116), .A3(new_n881), .A4(new_n901), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n900), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n706), .A2(new_n316), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT113), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n827), .B(new_n818), .C1(new_n498), .C2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n885), .A2(new_n746), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n892), .B1(new_n912), .B2(KEYINPUT51), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(KEYINPUT51), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT117), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n912), .A2(KEYINPUT117), .A3(KEYINPUT51), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n869), .A2(new_n879), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT119), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT119), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n869), .A2(new_n918), .A3(new_n921), .A4(new_n879), .ZN(new_n922));
  OR2_X1    g736(.A1(G952), .A2(G953), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n782), .A2(new_n497), .A3(new_n319), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n732), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT112), .Z(new_n927));
  NOR3_X1   g741(.A1(new_n927), .A2(new_n835), .A3(new_n696), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n909), .A2(KEYINPUT49), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n909), .A2(KEYINPUT49), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n924), .A2(new_n931), .ZN(G75));
  NAND2_X1  g746(.A1(new_n876), .A2(new_n878), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n933), .A2(G210), .A3(G902), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n465), .B1(new_n477), .B2(new_n479), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n935), .A2(new_n442), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(new_n480), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT55), .ZN(new_n938));
  XOR2_X1   g752(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n939));
  AND3_X1   g753(.A1(new_n934), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT56), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n938), .B1(new_n934), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n285), .A2(G952), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT121), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n940), .A2(new_n942), .A3(new_n945), .ZN(G51));
  XOR2_X1   g760(.A(new_n806), .B(KEYINPUT57), .Z(new_n947));
  AND3_X1   g761(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n877), .B1(new_n876), .B2(new_n878), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n315), .B2(new_n314), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n933), .A2(G902), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n952), .A2(new_n805), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n943), .B1(new_n951), .B2(new_n953), .ZN(G54));
  NAND2_X1  g768(.A1(KEYINPUT58), .A2(G475), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(new_n369), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n952), .A2(new_n363), .A3(new_n955), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n957), .A2(new_n943), .A3(new_n958), .ZN(G60));
  NAND2_X1  g773(.A1(G478), .A2(G902), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT59), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n634), .B(new_n961), .C1(new_n948), .C2(new_n949), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n944), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n869), .A2(new_n879), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n634), .B1(new_n964), .B2(new_n961), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n963), .A2(new_n965), .ZN(G63));
  XOR2_X1   g780(.A(new_n524), .B(KEYINPUT122), .Z(new_n967));
  AND2_X1   g781(.A1(new_n876), .A2(new_n878), .ZN(new_n968));
  NAND2_X1  g782(.A1(G217), .A2(G902), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT60), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n967), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n944), .B1(KEYINPUT123), .B2(KEYINPUT61), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n970), .B1(new_n876), .B2(new_n878), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n972), .B1(new_n973), .B2(new_n661), .ZN(new_n974));
  NAND2_X1  g788(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n971), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n975), .B1(new_n971), .B2(new_n974), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(G66));
  NAND2_X1  g792(.A1(G224), .A2(G953), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n379), .A2(new_n979), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n870), .A2(new_n858), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n980), .B1(new_n981), .B2(new_n285), .ZN(new_n982));
  INV_X1    g796(.A(new_n935), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(G898), .B2(new_n285), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n982), .B(new_n984), .ZN(G69));
  INV_X1    g799(.A(KEYINPUT126), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n814), .A2(new_n887), .A3(new_n624), .A4(new_n697), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n841), .A2(new_n702), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n816), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n771), .A2(new_n778), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(G953), .B1(new_n991), .B2(new_n831), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n285), .A2(G900), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n986), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n561), .A2(new_n563), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT124), .Z(new_n996));
  NOR2_X1   g810(.A1(new_n358), .A2(new_n359), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n996), .B(new_n997), .Z(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n826), .A2(new_n830), .ZN(new_n1000));
  INV_X1    g814(.A(new_n990), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n1001), .A2(new_n816), .A3(new_n988), .A4(new_n987), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n285), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n993), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1003), .A2(KEYINPUT126), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n994), .A2(new_n999), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT62), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n988), .A2(new_n699), .A3(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT125), .ZN(new_n1009));
  INV_X1    g823(.A(new_n816), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1007), .B1(new_n988), .B2(new_n699), .ZN(new_n1011));
  NOR4_X1   g825(.A1(new_n599), .A2(new_n683), .A3(new_n746), .A4(new_n849), .ZN(new_n1012));
  NOR3_X1   g826(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n1009), .A2(new_n831), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n998), .B1(new_n1014), .B2(G953), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1006), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n285), .B1(G227), .B2(G900), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1017), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1006), .A2(new_n1019), .A3(new_n1015), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1018), .A2(new_n1020), .ZN(G72));
  INV_X1    g835(.A(new_n688), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1014), .A2(new_n981), .ZN(new_n1023));
  XNOR2_X1  g837(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n608), .A2(new_n187), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1022), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n866), .A2(new_n868), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n564), .A2(new_n539), .A3(new_n549), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1022), .A2(new_n1029), .A3(new_n1026), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n991), .A2(new_n981), .A3(new_n831), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1029), .B1(new_n1032), .B2(new_n1026), .ZN(new_n1033));
  NOR4_X1   g847(.A1(new_n1027), .A2(new_n1031), .A3(new_n943), .A4(new_n1033), .ZN(G57));
endmodule


