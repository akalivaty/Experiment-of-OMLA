//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n559, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n581, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1208, new_n1209;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  NAND2_X1  g033(.A1(G101), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT66), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n470), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n471));
  OR2_X1    g046(.A1(new_n471), .A2(new_n467), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n466), .A2(new_n473), .A3(new_n467), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n469), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n470), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n464), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n467), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(KEYINPUT68), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n470), .A2(KEYINPUT67), .A3(G138), .A4(new_n467), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n488), .A2(KEYINPUT4), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n486), .B(new_n491), .C1(new_n487), .C2(KEYINPUT68), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n461), .A2(new_n463), .A3(G126), .ZN(new_n493));
  NAND2_X1  g068(.A1(G114), .A2(G2104), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n460), .A2(G2105), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n495), .A2(G2105), .B1(G102), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n490), .A2(new_n492), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G62), .ZN(new_n506));
  NAND2_X1  g081(.A1(G75), .A2(G543), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n500), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(G50), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OAI211_X1 g088(.A(new_n502), .B(new_n504), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n510), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT69), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n510), .B(new_n518), .C1(new_n514), .C2(new_n515), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n508), .B1(new_n517), .B2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT70), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT7), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n522), .B(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n513), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n501), .B1(new_n525), .B2(new_n511), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n509), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n502), .A2(new_n504), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT71), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g108(.A(KEYINPUT71), .B1(new_n524), .B2(new_n530), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(G168));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n529), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G651), .ZN(new_n539));
  XOR2_X1   g114(.A(new_n539), .B(KEYINPUT72), .Z(new_n540));
  NAND2_X1  g115(.A1(new_n509), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n541), .A2(new_n542), .B1(new_n514), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n540), .A2(new_n545), .ZN(G171));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n529), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n541), .A2(new_n552), .B1(new_n514), .B2(new_n553), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT73), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n526), .A2(new_n564), .A3(new_n565), .A4(G53), .ZN(new_n566));
  OAI211_X1 g141(.A(G53), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT9), .B1(new_n567), .B2(KEYINPUT74), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n514), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G91), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT75), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT76), .ZN(new_n574));
  AOI21_X1  g149(.A(KEYINPUT76), .B1(new_n502), .B2(new_n504), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n573), .B1(new_n576), .B2(G65), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n569), .B(new_n571), .C1(new_n577), .C2(new_n500), .ZN(G299));
  NAND2_X1  g153(.A1(new_n540), .A2(new_n545), .ZN(G301));
  INV_X1    g154(.A(G168), .ZN(G286));
  INV_X1    g155(.A(new_n508), .ZN(new_n581));
  INV_X1    g156(.A(new_n519), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n505), .A2(G88), .A3(new_n509), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n518), .B1(new_n583), .B2(new_n510), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n581), .B1(new_n582), .B2(new_n584), .ZN(G303));
  NAND2_X1  g160(.A1(new_n570), .A2(G87), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n526), .A2(G49), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(new_n505), .A2(G61), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G651), .ZN(new_n593));
  INV_X1    g168(.A(G48), .ZN(new_n594));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n541), .A2(new_n594), .B1(new_n514), .B2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(G305));
  INV_X1    g173(.A(G47), .ZN(new_n599));
  INV_X1    g174(.A(G85), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n541), .A2(new_n599), .B1(new_n514), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(G72), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G60), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n529), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G651), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n602), .A2(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n576), .A2(G66), .ZN(new_n609));
  INV_X1    g184(.A(G79), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n501), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n526), .B(KEYINPUT77), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n611), .A2(G651), .B1(G54), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n570), .A2(G92), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT10), .Z(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n608), .B1(new_n617), .B2(G868), .ZN(G284));
  XNOR2_X1  g193(.A(G284), .B(KEYINPUT78), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  INV_X1    g195(.A(G299), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(G868), .B2(new_n621), .ZN(G297));
  OAI21_X1  g197(.A(new_n620), .B1(G868), .B2(new_n621), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(new_n624), .B2(G860), .ZN(G148));
  NOR2_X1   g200(.A1(new_n616), .A2(G559), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT79), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n470), .A2(new_n496), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT12), .Z(new_n632));
  XOR2_X1   g207(.A(KEYINPUT13), .B(G2100), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n478), .A2(G123), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n480), .A2(G135), .ZN(new_n636));
  NOR2_X1   g211(.A1(G99), .A2(G2105), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(new_n467), .B2(G111), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT80), .Z(new_n640));
  AND2_X1   g215(.A1(new_n640), .A2(G2096), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n640), .A2(G2096), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n634), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT81), .Z(G156));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2435), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2438), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT14), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G1341), .B(G1348), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT82), .Z(new_n657));
  OR2_X1    g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n658), .A2(G14), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT83), .Z(G401));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2067), .B(G2678), .Z(new_n664));
  XNOR2_X1  g239(.A(G2072), .B(G2078), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n663), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT84), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT18), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n665), .B(KEYINPUT17), .Z(new_n670));
  NAND3_X1  g245(.A1(new_n670), .A2(new_n664), .A3(new_n662), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT85), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n666), .A2(new_n664), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n663), .B(new_n673), .C1(new_n670), .C2(new_n664), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n669), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(G2096), .Z(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(G2100), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT86), .ZN(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1971), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n680), .A2(new_n681), .ZN(new_n687));
  AOI22_X1  g262(.A1(new_n685), .A2(new_n686), .B1(new_n684), .B2(new_n687), .ZN(new_n688));
  OR3_X1    g263(.A1(new_n682), .A2(new_n687), .A3(new_n684), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n688), .B(new_n689), .C1(new_n686), .C2(new_n685), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(G1986), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT22), .B(G1981), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n694), .B(new_n695), .Z(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  NAND2_X1  g272(.A1(new_n475), .A2(G29), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  INV_X1    g274(.A(G34), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n700), .A2(KEYINPUT24), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(KEYINPUT24), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n704), .A2(G2084), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT96), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n480), .A2(G139), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT94), .ZN(new_n708));
  AOI22_X1  g283(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n709), .A2(new_n467), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n496), .A2(G103), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT25), .Z(new_n712));
  NAND3_X1  g287(.A1(new_n708), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n713), .A2(new_n699), .ZN(new_n714));
  INV_X1    g289(.A(G33), .ZN(new_n715));
  AOI21_X1  g290(.A(KEYINPUT93), .B1(new_n699), .B2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT93), .ZN(new_n717));
  NOR3_X1   g292(.A1(new_n717), .A2(G29), .A3(G33), .ZN(new_n718));
  NOR3_X1   g293(.A1(new_n714), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(G2072), .ZN(new_n720));
  OR2_X1    g295(.A1(G29), .A2(G32), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n478), .A2(G129), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n496), .A2(G105), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n480), .A2(G141), .ZN(new_n724));
  NAND3_X1  g299(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT26), .Z(new_n726));
  NAND4_X1  g301(.A1(new_n722), .A2(new_n723), .A3(new_n724), .A4(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n721), .B1(new_n727), .B2(new_n699), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT27), .B(G1996), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT30), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(G28), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(G28), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n732), .A2(new_n733), .A3(new_n699), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n706), .A2(new_n720), .A3(new_n730), .A4(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(G16), .A2(G19), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n556), .B2(G16), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1341), .ZN(new_n738));
  NOR2_X1   g313(.A1(G29), .A2(G35), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G162), .B2(G29), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT29), .B(G2090), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n728), .A2(new_n729), .ZN(new_n743));
  INV_X1    g318(.A(new_n640), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT95), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n744), .A2(new_n745), .A3(new_n699), .ZN(new_n746));
  AOI21_X1  g321(.A(KEYINPUT95), .B1(new_n640), .B2(G29), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n743), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR4_X1   g323(.A1(new_n735), .A2(new_n738), .A3(new_n742), .A4(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G16), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n750), .A2(KEYINPUT23), .A3(G20), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT23), .ZN(new_n752));
  INV_X1    g327(.A(G20), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(G16), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n751), .B(new_n754), .C1(new_n621), .C2(new_n750), .ZN(new_n755));
  INV_X1    g330(.A(G1956), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G4), .B2(G16), .ZN(new_n759));
  OR3_X1    g334(.A1(new_n758), .A2(G4), .A3(G16), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n759), .B(new_n760), .C1(new_n616), .C2(new_n750), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT90), .B(G1348), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n699), .A2(G27), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G164), .B2(new_n699), .ZN(new_n765));
  MUX2_X1   g340(.A(new_n764), .B(new_n765), .S(KEYINPUT97), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT98), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n757), .B(new_n763), .C1(new_n767), .C2(G2078), .ZN(new_n768));
  INV_X1    g343(.A(G11), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n719), .A2(G2072), .B1(KEYINPUT31), .B2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT28), .ZN(new_n771));
  INV_X1    g346(.A(G26), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G29), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n772), .A2(G29), .ZN(new_n774));
  INV_X1    g349(.A(G116), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n460), .B1(new_n775), .B2(G2105), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT91), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G104), .B2(G2105), .ZN(new_n778));
  INV_X1    g353(.A(G104), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n779), .A2(new_n467), .A3(KEYINPUT91), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n776), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT92), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n478), .A2(G128), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n480), .A2(G140), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n774), .B1(new_n785), .B2(G29), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n773), .B1(new_n786), .B2(new_n771), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G2067), .ZN(new_n788));
  NAND2_X1  g363(.A1(G168), .A2(G16), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G16), .B2(G21), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n790), .A2(G1966), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n790), .A2(G1966), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n770), .B(new_n788), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n768), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n704), .A2(G2084), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n767), .A2(G2078), .ZN(new_n796));
  AND4_X1   g371(.A1(new_n749), .A2(new_n794), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(G290), .A2(G16), .ZN(new_n798));
  INV_X1    g373(.A(G24), .ZN(new_n799));
  OAI21_X1  g374(.A(KEYINPUT87), .B1(new_n799), .B2(G16), .ZN(new_n800));
  OR3_X1    g375(.A1(new_n799), .A2(KEYINPUT87), .A3(G16), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n798), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1986), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n699), .A2(G25), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n478), .A2(G119), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n480), .A2(G131), .ZN(new_n806));
  OR2_X1    g381(.A1(G95), .A2(G2105), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n807), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n805), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n804), .B1(new_n810), .B2(new_n699), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT35), .B(G1991), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n803), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT34), .ZN(new_n817));
  NAND2_X1  g392(.A1(G305), .A2(G16), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n750), .A2(G6), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT32), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT32), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n818), .A2(new_n822), .A3(new_n819), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT88), .B(G1981), .Z(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n824), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n750), .A2(G22), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G166), .B2(new_n750), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(G1971), .Z(new_n830));
  NOR2_X1   g405(.A1(G16), .A2(G23), .ZN(new_n831));
  INV_X1    g406(.A(G288), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n831), .B1(new_n832), .B2(G16), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT33), .B(G1976), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n830), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n817), .B1(new_n827), .B2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  NOR3_X1   g413(.A1(new_n827), .A2(new_n836), .A3(new_n817), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n816), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT36), .ZN(new_n841));
  OR3_X1    g416(.A1(new_n827), .A2(new_n836), .A3(new_n817), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(new_n837), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT36), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n843), .A2(new_n844), .A3(new_n816), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(G171), .A2(new_n750), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(G5), .B2(new_n750), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(G1961), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n797), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT99), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n787), .A2(G2067), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n769), .A2(KEYINPUT31), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n850), .A2(new_n851), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n797), .A2(new_n846), .A3(new_n854), .A4(new_n849), .ZN(new_n856));
  OAI21_X1  g431(.A(KEYINPUT99), .B1(new_n856), .B2(new_n852), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(G311));
  NAND4_X1  g433(.A1(new_n850), .A2(KEYINPUT100), .A3(new_n853), .A4(new_n854), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n856), .B2(new_n852), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(G150));
  AOI22_X1  g437(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(new_n500), .ZN(new_n864));
  INV_X1    g439(.A(G55), .ZN(new_n865));
  INV_X1    g440(.A(G93), .ZN(new_n866));
  OAI22_X1  g441(.A1(new_n541), .A2(new_n865), .B1(new_n514), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(G860), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT37), .Z(new_n869));
  NOR2_X1   g444(.A1(new_n616), .A2(new_n624), .ZN(new_n870));
  XNOR2_X1  g445(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT39), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n870), .B(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n864), .A2(new_n867), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n555), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n873), .B(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n869), .B1(new_n877), .B2(G860), .ZN(G145));
  NAND2_X1  g453(.A1(new_n478), .A2(G130), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n480), .A2(G142), .ZN(new_n880));
  OR2_X1    g455(.A1(G106), .A2(G2105), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n881), .B(G2104), .C1(G118), .C2(new_n467), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n632), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n809), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT102), .Z(new_n886));
  XNOR2_X1  g461(.A(new_n785), .B(new_n498), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n727), .ZN(new_n888));
  INV_X1    g463(.A(new_n713), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n888), .B(new_n713), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n885), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n475), .B(new_n484), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n640), .B(new_n894), .Z(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n891), .A2(new_n893), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n891), .A2(new_n893), .A3(KEYINPUT104), .A4(new_n896), .ZN(new_n900));
  AOI21_X1  g475(.A(G37), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n886), .A2(new_n890), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(KEYINPUT103), .A3(new_n891), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n886), .A2(new_n904), .A3(new_n890), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n905), .A3(new_n895), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n901), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g483(.A1(new_n627), .A2(new_n875), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n616), .A2(G299), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n621), .A2(new_n613), .A3(new_n615), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n627), .A2(new_n875), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n909), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n909), .A2(new_n913), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n910), .A2(new_n916), .A3(new_n911), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n916), .B1(new_n910), .B2(new_n911), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n914), .B1(new_n915), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT42), .ZN(new_n922));
  XNOR2_X1  g497(.A(G305), .B(KEYINPUT105), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(G303), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n832), .B(G290), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT106), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n925), .A2(KEYINPUT106), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n924), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n914), .B(new_n933), .C1(new_n915), .C2(new_n920), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n922), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n932), .B1(new_n922), .B2(new_n934), .ZN(new_n936));
  OAI21_X1  g511(.A(G868), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(G868), .B2(new_n874), .ZN(G295));
  OAI21_X1  g513(.A(new_n937), .B1(G868), .B2(new_n874), .ZN(G331));
  INV_X1    g514(.A(new_n912), .ZN(new_n940));
  NOR2_X1   g515(.A1(G171), .A2(G168), .ZN(new_n941));
  AOI21_X1  g516(.A(G301), .B1(new_n534), .B2(new_n533), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n941), .A2(new_n942), .A3(new_n875), .ZN(new_n943));
  NAND2_X1  g518(.A1(G286), .A2(G301), .ZN(new_n944));
  NAND2_X1  g519(.A1(G171), .A2(G168), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n876), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n940), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n875), .B1(new_n941), .B2(new_n942), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n944), .A2(new_n876), .A3(new_n945), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n948), .B(new_n949), .C1(new_n917), .C2(new_n918), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT107), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n947), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(new_n932), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n951), .ZN(new_n956));
  AOI21_X1  g531(.A(G37), .B1(new_n956), .B2(new_n931), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  OR3_X1    g533(.A1(new_n958), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n919), .A2(KEYINPUT109), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n943), .A2(new_n946), .ZN(new_n962));
  OR3_X1    g537(.A1(new_n912), .A2(KEYINPUT109), .A3(KEYINPUT41), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(KEYINPUT110), .A3(new_n947), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n961), .A2(new_n966), .A3(new_n962), .A4(new_n963), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n932), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n957), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n960), .B1(new_n969), .B2(KEYINPUT43), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT111), .B1(new_n958), .B2(KEYINPUT43), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n959), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n947), .A2(new_n950), .A3(new_n953), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n953), .B1(new_n947), .B2(new_n950), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n974), .A2(new_n975), .A3(new_n931), .ZN(new_n976));
  INV_X1    g551(.A(G37), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n932), .B2(new_n951), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n973), .B(KEYINPUT43), .C1(new_n976), .C2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT43), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n968), .A2(new_n980), .A3(new_n957), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n973), .B1(new_n958), .B2(KEYINPUT43), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n960), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n972), .A2(new_n984), .ZN(G397));
  INV_X1    g560(.A(G1384), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n488), .A2(KEYINPUT4), .A3(new_n489), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n495), .A2(G2105), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n496), .A2(G102), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n492), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n986), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n469), .A2(new_n472), .A3(G40), .A4(new_n474), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G2067), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n785), .B(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n809), .A2(new_n812), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n809), .A2(new_n812), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n727), .B(G1996), .ZN(new_n1001));
  NOR4_X1   g576(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(G290), .A2(G1986), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(G290), .A2(G1986), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n995), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G8), .ZN(new_n1007));
  NOR2_X1   g582(.A1(G168), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT51), .B1(new_n1008), .B2(KEYINPUT125), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n994), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n986), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n993), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1966), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT117), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n991), .A2(KEYINPUT50), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1019), .B(new_n986), .C1(new_n987), .C2(new_n990), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1018), .A2(new_n1012), .A3(new_n1020), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n1021), .A2(G2084), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1014), .A2(new_n1023), .A3(new_n1015), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1017), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1009), .B(new_n1011), .C1(new_n1025), .C2(new_n1007), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1017), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1027));
  OAI211_X1 g602(.A(G8), .B(new_n1010), .C1(new_n1027), .C2(G286), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT124), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n1029), .A3(new_n1008), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1029), .B1(new_n1027), .B2(new_n1008), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1026), .B(new_n1028), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT62), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1032), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n1030), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT62), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1036), .A2(new_n1037), .A3(new_n1028), .A4(new_n1026), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT126), .ZN(new_n1039));
  INV_X1    g614(.A(G2078), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n993), .A2(new_n1040), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n994), .B1(new_n991), .B2(KEYINPUT50), .ZN(new_n1044));
  AOI21_X1  g619(.A(G1961), .B1(new_n1044), .B2(new_n1020), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1039), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1047));
  INV_X1    g622(.A(G1961), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1021), .A2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1049), .B(KEYINPUT126), .C1(new_n1042), .C2(new_n1041), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1046), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(G171), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT112), .B(G1971), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1014), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G2090), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1044), .A2(new_n1057), .A3(new_n1020), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  XOR2_X1   g634(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(G166), .B2(new_n1007), .ZN(new_n1061));
  NOR2_X1   g636(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1062));
  NAND3_X1  g637(.A1(G303), .A2(G8), .A3(new_n1062), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1061), .A2(new_n1063), .A3(KEYINPUT114), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT114), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1059), .A2(new_n1066), .A3(G8), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n991), .A2(new_n994), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n500), .B1(new_n590), .B2(new_n591), .ZN(new_n1070));
  OR3_X1    g645(.A1(new_n1070), .A2(new_n596), .A3(G1981), .ZN(new_n1071));
  OAI21_X1  g646(.A(G1981), .B1(new_n1070), .B2(new_n596), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT49), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1071), .A2(KEYINPUT49), .A3(new_n1072), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1069), .A2(new_n1075), .A3(G8), .A4(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n832), .A2(G1976), .ZN(new_n1078));
  INV_X1    g653(.A(G1976), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT52), .B1(G288), .B2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1069), .A2(G8), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1078), .B(G8), .C1(new_n991), .C2(new_n994), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT52), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1077), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1067), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1020), .A2(KEYINPUT115), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n498), .A2(new_n1088), .A3(new_n1019), .A4(new_n986), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1044), .A2(new_n1087), .A3(new_n1057), .A4(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1056), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT116), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT116), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1056), .A2(new_n1093), .A3(new_n1090), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(G8), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1085), .B1(new_n1086), .B2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1034), .A2(new_n1038), .A3(new_n1053), .A4(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1044), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n756), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1013), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT45), .B1(new_n498), .B2(new_n986), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT56), .B(G2072), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n1012), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1099), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(G299), .A2(KEYINPUT119), .ZN(new_n1106));
  INV_X1    g681(.A(G65), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n574), .A2(new_n575), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(G651), .B1(new_n1108), .B2(new_n573), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1109), .A2(new_n1110), .A3(new_n569), .A4(new_n571), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1106), .A2(KEYINPUT57), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT57), .B1(new_n1106), .B2(new_n1111), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1105), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(G1348), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1021), .A2(new_n1117), .B1(new_n996), .B2(new_n1068), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1116), .B1(new_n616), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1114), .A2(new_n1099), .A3(new_n1104), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1114), .A2(new_n1099), .A3(new_n1104), .A4(new_n1122), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1119), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1121), .A2(new_n1116), .A3(new_n1123), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n1127));
  AND3_X1   g702(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1126), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1116), .A2(KEYINPUT61), .A3(new_n1120), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT58), .B(G1341), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1014), .A2(G1996), .B1(new_n1068), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n556), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1134), .A2(KEYINPUT59), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1134), .A2(KEYINPUT59), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1131), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n617), .B1(new_n1118), .B2(KEYINPUT60), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g715(.A(KEYINPUT123), .B(new_n617), .C1(new_n1118), .C2(KEYINPUT60), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1142), .A2(KEYINPUT60), .A3(new_n1118), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1118), .A2(KEYINPUT60), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1140), .A2(new_n1144), .A3(new_n1141), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1137), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1124), .B1(new_n1130), .B2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1102), .A2(KEYINPUT53), .A3(new_n1040), .A4(new_n1012), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1148), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(G171), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1150), .B(KEYINPUT54), .C1(new_n1051), .C2(G171), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1096), .A2(new_n1151), .ZN(new_n1152));
  AND4_X1   g727(.A1(G301), .A2(new_n1148), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1052), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n1156));
  AOI21_X1  g731(.A(KEYINPUT127), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1153), .B1(new_n1051), .B2(G171), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1158), .A2(new_n1159), .A3(KEYINPUT54), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1033), .B(new_n1152), .C1(new_n1157), .C2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1097), .B1(new_n1147), .B2(new_n1161), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1025), .A2(new_n1007), .A3(G286), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1085), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1095), .A2(new_n1086), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT63), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1007), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1086), .ZN(new_n1169));
  OAI21_X1  g744(.A(KEYINPUT63), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1085), .A2(new_n1170), .ZN(new_n1171));
  AOI22_X1  g746(.A1(new_n1166), .A2(new_n1167), .B1(new_n1163), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1067), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1077), .A2(new_n1079), .A3(new_n832), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(new_n1071), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1068), .A2(new_n1007), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1173), .A2(new_n1084), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT118), .B1(new_n1172), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT118), .ZN(new_n1180));
  AOI21_X1  g755(.A(KEYINPUT63), .B1(new_n1096), .B2(new_n1163), .ZN(new_n1181));
  AND2_X1   g756(.A1(new_n1171), .A2(new_n1163), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1180), .B(new_n1177), .C1(new_n1181), .C2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1179), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1006), .B1(new_n1162), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n995), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n998), .A2(new_n1001), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(new_n1000), .ZN(new_n1188));
  OR2_X1    g763(.A1(new_n785), .A2(G2067), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1186), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT46), .ZN(new_n1191));
  OR3_X1    g766(.A1(new_n1186), .A2(new_n1191), .A3(G1996), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n995), .B1(new_n998), .B2(new_n727), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1191), .B1(new_n1186), .B2(G1996), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  XOR2_X1   g770(.A(new_n1195), .B(KEYINPUT47), .Z(new_n1196));
  OR2_X1    g771(.A1(new_n1002), .A2(new_n1186), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n995), .A2(new_n1005), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1198), .B(KEYINPUT48), .ZN(new_n1199));
  AOI211_X1 g774(.A(new_n1190), .B(new_n1196), .C1(new_n1197), .C2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1185), .A2(new_n1200), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g776(.A(G319), .B(new_n696), .C1(new_n982), .C2(new_n983), .ZN(new_n1203));
  NAND2_X1  g777(.A1(new_n660), .A2(new_n677), .ZN(new_n1204));
  AOI21_X1  g778(.A(new_n1204), .B1(new_n901), .B2(new_n906), .ZN(new_n1205));
  INV_X1    g779(.A(new_n1205), .ZN(new_n1206));
  NOR2_X1   g780(.A1(new_n1203), .A2(new_n1206), .ZN(G308));
  INV_X1    g781(.A(new_n983), .ZN(new_n1208));
  NAND3_X1  g782(.A1(new_n1208), .A2(new_n981), .A3(new_n979), .ZN(new_n1209));
  NAND4_X1  g783(.A1(new_n1209), .A2(G319), .A3(new_n696), .A4(new_n1205), .ZN(G225));
endmodule


