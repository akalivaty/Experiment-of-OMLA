//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT66), .A2(G128), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT66), .A2(G128), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n196), .B1(G143), .B2(new_n188), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n192), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G125), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n200), .B1(new_n190), .B2(G146), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n188), .A2(KEYINPUT64), .A3(G143), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G128), .A4(new_n191), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n198), .B(new_n199), .C1(KEYINPUT1), .C2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT80), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n201), .A2(new_n191), .A3(new_n202), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(new_n196), .A3(G128), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n208), .A2(KEYINPUT80), .A3(new_n199), .A4(new_n198), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT0), .A2(G128), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT0), .ZN(new_n212));
  INV_X1    g026(.A(G128), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n192), .A2(new_n211), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(new_n212), .B2(new_n203), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G125), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT81), .B(G224), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(G953), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n219), .B(KEYINPUT82), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n210), .A2(new_n217), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n220), .B1(new_n210), .B2(new_n217), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G119), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G116), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n226));
  INV_X1    g040(.A(G116), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n226), .B1(new_n227), .B2(G119), .ZN(new_n228));
  NOR3_X1   g042(.A1(new_n224), .A2(KEYINPUT67), .A3(G116), .ZN(new_n229));
  OAI211_X1 g043(.A(KEYINPUT5), .B(new_n225), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(G113), .B1(new_n225), .B2(KEYINPUT5), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n227), .A2(G119), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT67), .B1(new_n224), .B2(G116), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n226), .A2(new_n227), .A3(G119), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  XOR2_X1   g050(.A(KEYINPUT2), .B(G113), .Z(new_n237));
  AOI22_X1  g051(.A1(new_n230), .A2(new_n232), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G104), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT3), .B1(new_n239), .B2(G107), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n241));
  INV_X1    g055(.A(G107), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n242), .A3(G104), .ZN(new_n243));
  INV_X1    g057(.A(G101), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n239), .A2(G107), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n240), .A2(new_n243), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n239), .A2(G107), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n242), .A2(G104), .ZN(new_n248));
  OAI21_X1  g062(.A(G101), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT78), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT78), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n246), .A2(new_n249), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n238), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n240), .A2(new_n243), .A3(new_n245), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT76), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n255), .A2(new_n256), .A3(G101), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n256), .B1(new_n255), .B2(G101), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n246), .A2(KEYINPUT4), .ZN(new_n259));
  NOR3_X1   g073(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n255), .A2(new_n261), .A3(G101), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n236), .A2(new_n237), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n236), .A2(new_n237), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n254), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G110), .B(G122), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n254), .B(new_n267), .C1(new_n260), .C2(new_n265), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(KEYINPUT6), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n266), .A2(new_n272), .A3(new_n268), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n223), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT83), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT83), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n223), .A2(new_n271), .A3(new_n276), .A4(new_n273), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n250), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n231), .B1(new_n236), .B2(KEYINPUT5), .ZN(new_n280));
  OAI221_X1 g094(.A(new_n279), .B1(new_n252), .B2(KEYINPUT84), .C1(new_n263), .C2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n267), .B(KEYINPUT8), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n251), .A2(KEYINPUT84), .A3(new_n253), .ZN(new_n283));
  INV_X1    g097(.A(new_n238), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n281), .B(new_n282), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT7), .B1(new_n218), .B2(G953), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n210), .A2(new_n217), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n285), .A2(new_n288), .A3(new_n270), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT85), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n210), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n206), .A2(KEYINPUT85), .A3(new_n209), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n217), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n286), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n289), .B1(new_n294), .B2(KEYINPUT86), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT86), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n293), .A2(new_n296), .A3(new_n286), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G210), .B1(G237), .B2(G902), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n278), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n299), .B1(new_n278), .B2(new_n298), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n187), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G902), .ZN(new_n303));
  XNOR2_X1  g117(.A(G113), .B(G122), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n304), .B(new_n239), .ZN(new_n305));
  INV_X1    g119(.A(G237), .ZN(new_n306));
  INV_X1    g120(.A(G953), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n307), .A3(G214), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT87), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(new_n190), .ZN(new_n310));
  NOR2_X1   g124(.A1(KEYINPUT87), .A2(G143), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n308), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n311), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n313), .A2(G214), .A3(new_n306), .A4(new_n307), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(KEYINPUT18), .A3(G131), .ZN(new_n316));
  NAND2_X1  g130(.A1(KEYINPUT18), .A2(G131), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n312), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(new_n188), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n316), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n315), .A2(KEYINPUT17), .A3(G131), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT89), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT89), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n315), .A2(new_n324), .A3(KEYINPUT17), .A4(G131), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G140), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G125), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n199), .A2(G140), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(KEYINPUT16), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT16), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n327), .A3(G125), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT71), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n331), .A2(new_n327), .A3(KEYINPUT71), .A4(G125), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n330), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n188), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n330), .A2(new_n334), .A3(G146), .A4(new_n335), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n315), .A2(G131), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT17), .ZN(new_n342));
  INV_X1    g156(.A(G131), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n312), .A2(new_n314), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n305), .B(new_n321), .C1(new_n326), .C2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n323), .A2(new_n325), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n340), .A3(new_n345), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n305), .B1(new_n350), .B2(new_n321), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n303), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G475), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n307), .A2(G952), .ZN(new_n354));
  INV_X1    g168(.A(G234), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n354), .B1(new_n355), .B2(new_n306), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AOI211_X1 g171(.A(new_n303), .B(new_n307), .C1(G234), .C2(G237), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT21), .B(G898), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n321), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n341), .A2(new_n344), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT88), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n319), .A2(KEYINPUT19), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n319), .A2(KEYINPUT19), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n188), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n364), .B1(new_n367), .B2(new_n338), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n364), .A3(new_n338), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n362), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n347), .B1(new_n371), .B2(new_n305), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT20), .ZN(new_n373));
  NOR2_X1   g187(.A1(G475), .A2(G902), .ZN(new_n374));
  XOR2_X1   g188(.A(new_n374), .B(KEYINPUT90), .Z(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n372), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n373), .B1(new_n372), .B2(new_n376), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n353), .B(new_n361), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(G110), .B(G140), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n307), .A2(G227), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n381), .B(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT11), .ZN(new_n384));
  INV_X1    g198(.A(G134), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n384), .B1(new_n385), .B2(G137), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(G137), .ZN(new_n387));
  INV_X1    g201(.A(G137), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(KEYINPUT11), .A3(G134), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G131), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n386), .A2(new_n389), .A3(new_n343), .A4(new_n387), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  OR3_X1    g208(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n207), .A2(KEYINPUT0), .A3(G128), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n215), .A3(new_n262), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n253), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n252), .B1(new_n246), .B2(new_n249), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT10), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n402), .B1(new_n208), .B2(new_n198), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n395), .A2(new_n398), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT77), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n207), .A2(new_n405), .A3(new_n196), .A4(G128), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n201), .A2(new_n191), .A3(new_n202), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n407), .B1(new_n213), .B2(new_n197), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT77), .B1(new_n203), .B2(KEYINPUT1), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n406), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT10), .B1(new_n410), .B2(new_n279), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n394), .B1(new_n404), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n198), .B1(KEYINPUT1), .B2(new_n203), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n251), .A2(new_n414), .A3(KEYINPUT10), .A4(new_n253), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n260), .B2(new_n397), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n416), .A2(new_n411), .A3(new_n393), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n383), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n404), .A2(new_n412), .A3(new_n394), .ZN(new_n419));
  INV_X1    g233(.A(new_n383), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n410), .A2(new_n279), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n198), .B(new_n208), .C1(new_n399), .C2(new_n400), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT12), .B1(new_n423), .B2(new_n393), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT12), .ZN(new_n425));
  AOI211_X1 g239(.A(new_n425), .B(new_n394), .C1(new_n421), .C2(new_n422), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n419), .B(new_n420), .C1(new_n424), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n418), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G469), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n429), .A3(new_n303), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT79), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n417), .B2(new_n383), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n419), .A2(KEYINPUT79), .A3(new_n420), .ZN(new_n433));
  INV_X1    g247(.A(new_n413), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n419), .B1(new_n424), .B2(new_n426), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n383), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(new_n437), .A3(G469), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n429), .A2(new_n303), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n430), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G478), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(KEYINPUT15), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G122), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G116), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n227), .A2(G122), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(new_n242), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT91), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n449), .B1(new_n213), .B2(G143), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n190), .A2(KEYINPUT91), .A3(G128), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OR2_X1    g266(.A1(KEYINPUT66), .A2(G128), .ZN(new_n453));
  NAND2_X1  g267(.A1(KEYINPUT66), .A2(G128), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(G143), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n452), .A2(new_n455), .A3(new_n385), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n385), .B1(new_n452), .B2(new_n455), .ZN(new_n458));
  OR2_X1    g272(.A1(new_n447), .A2(KEYINPUT14), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT94), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(new_n446), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n461), .B1(KEYINPUT14), .B2(new_n447), .ZN(new_n462));
  OAI21_X1  g276(.A(G107), .B1(new_n459), .B2(new_n460), .ZN(new_n463));
  OAI221_X1 g277(.A(new_n448), .B1(new_n457), .B2(new_n458), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT13), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n190), .A2(KEYINPUT91), .A3(G128), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT91), .B1(new_n190), .B2(G128), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT92), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n469), .A3(new_n455), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT13), .B1(new_n450), .B2(new_n451), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n193), .A2(new_n194), .A3(new_n190), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT92), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n450), .A2(KEYINPUT13), .A3(new_n451), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G134), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n446), .A2(new_n447), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G107), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n448), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n456), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(KEYINPUT93), .B1(new_n476), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT93), .ZN(new_n483));
  AOI211_X1 g297(.A(new_n483), .B(new_n480), .C1(new_n475), .C2(G134), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n464), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT9), .B(G234), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(G217), .A3(new_n307), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n488), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n464), .B(new_n490), .C1(new_n482), .C2(new_n484), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n444), .B1(new_n492), .B2(new_n303), .ZN(new_n493));
  AOI211_X1 g307(.A(G902), .B(new_n443), .C1(new_n489), .C2(new_n491), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G221), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n496), .B1(new_n487), .B2(new_n303), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n497), .B(KEYINPUT75), .Z(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n380), .A2(new_n441), .A3(new_n495), .A4(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n302), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT31), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT28), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n263), .A2(new_n264), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n216), .B1(new_n392), .B2(new_n391), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n388), .A2(KEYINPUT65), .A3(G134), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT65), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n508), .B1(new_n388), .B2(G134), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n385), .A2(G137), .ZN(new_n510));
  OAI211_X1 g324(.A(G131), .B(new_n507), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n392), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(new_n208), .B2(new_n198), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n505), .B1(new_n506), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n393), .A2(new_n396), .A3(new_n215), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n511), .A2(new_n392), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n414), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n517), .A3(new_n504), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n503), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n503), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n306), .A2(new_n307), .A3(G210), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT27), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT26), .B(G101), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n519), .A2(new_n521), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n525), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n515), .A2(new_n517), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n528), .B1(new_n515), .B2(new_n517), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n505), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n527), .B1(new_n532), .B2(new_n518), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n502), .B1(new_n526), .B2(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n532), .A2(KEYINPUT31), .A3(new_n518), .A4(new_n525), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n535), .A2(new_n303), .ZN(new_n536));
  INV_X1    g350(.A(G472), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n534), .A2(new_n536), .A3(KEYINPUT32), .A4(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n525), .B1(new_n519), .B2(new_n521), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n532), .A2(new_n518), .A3(new_n527), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT29), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n515), .A2(new_n517), .A3(new_n504), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n504), .B1(new_n515), .B2(new_n517), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT28), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n544), .A2(KEYINPUT29), .A3(new_n525), .A4(new_n520), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n303), .ZN(new_n546));
  OAI21_X1  g360(.A(G472), .B1(new_n541), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT30), .B1(new_n506), .B2(new_n513), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n504), .B1(new_n548), .B2(new_n529), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n525), .B1(new_n549), .B2(new_n542), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n544), .A2(new_n527), .A3(new_n520), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT31), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n535), .A2(new_n303), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n552), .A2(new_n553), .A3(G472), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT68), .B(KEYINPUT32), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n538), .B(new_n547), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(G217), .B1(new_n355), .B2(G902), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n328), .A2(new_n329), .ZN(new_n558));
  INV_X1    g372(.A(G110), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT24), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT24), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G110), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT69), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n563), .B1(new_n560), .B2(new_n562), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n213), .A2(G119), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n567), .B1(new_n195), .B2(G119), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT23), .B1(new_n213), .B2(G119), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT70), .B1(new_n224), .B2(G128), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT70), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(new_n213), .A3(G119), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n453), .A2(KEYINPUT23), .A3(G119), .A4(new_n454), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n576), .A2(G110), .ZN(new_n577));
  OAI221_X1 g391(.A(new_n338), .B1(G146), .B2(new_n558), .C1(new_n569), .C2(new_n577), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n566), .A2(new_n568), .B1(new_n576), .B2(G110), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT72), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n579), .A2(new_n339), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n580), .B1(new_n579), .B2(new_n339), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n578), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT22), .B(G137), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n496), .A2(new_n355), .A3(G953), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n584), .B(new_n585), .Z(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n578), .B(new_n586), .C1(new_n581), .C2(new_n582), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n303), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT73), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT25), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n557), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n590), .A2(new_n591), .A3(KEYINPUT25), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n557), .A2(new_n303), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT74), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n588), .A2(new_n589), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n594), .A2(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n556), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n501), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT95), .B(G101), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G3));
  NAND2_X1  g418(.A1(new_n278), .A2(new_n298), .ZN(new_n605));
  INV_X1    g419(.A(new_n299), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT96), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n278), .A2(new_n298), .A3(new_n299), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n278), .A2(new_n298), .A3(KEYINPUT96), .A4(new_n299), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n611), .A2(new_n187), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n368), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n341), .A2(new_n344), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n614), .A2(new_n615), .A3(new_n370), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n305), .B1(new_n616), .B2(new_n321), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n376), .B1(new_n348), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(KEYINPUT20), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n372), .A2(new_n373), .A3(new_n376), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n619), .A2(new_n620), .B1(G475), .B2(new_n352), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n442), .A2(G902), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n489), .A2(new_n623), .A3(new_n491), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n623), .B1(new_n489), .B2(new_n491), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT97), .B(G478), .Z(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n492), .B2(new_n303), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n621), .B1(new_n626), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n360), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n613), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(G902), .B1(new_n418), .B2(new_n427), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n439), .B1(new_n635), .B2(new_n429), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n498), .B1(new_n636), .B2(new_n438), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n599), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n640));
  OAI21_X1  g454(.A(G472), .B1(new_n552), .B2(new_n553), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n638), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n634), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT34), .B(G104), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  OAI21_X1  g461(.A(new_n353), .B1(new_n377), .B2(new_n378), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n495), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n361), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n613), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n644), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT35), .B(G107), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  AND3_X1   g469(.A1(new_n590), .A2(new_n591), .A3(KEYINPUT25), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT25), .B1(new_n590), .B2(new_n591), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n656), .A2(new_n657), .A3(new_n557), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n587), .A2(KEYINPUT36), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n583), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n583), .A2(new_n660), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n597), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(KEYINPUT98), .B1(new_n658), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n642), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n594), .A2(new_n595), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT98), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n668), .A2(new_n669), .A3(new_n664), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n666), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT99), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n666), .A2(new_n670), .A3(KEYINPUT99), .A4(new_n667), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n673), .A2(new_n501), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  AND4_X1   g491(.A1(new_n556), .A2(new_n666), .A3(new_n637), .A4(new_n670), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n678), .A2(new_n613), .ZN(new_n679));
  INV_X1    g493(.A(new_n358), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n356), .B1(new_n680), .B2(G900), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n649), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G128), .ZN(G30));
  NOR2_X1   g499(.A1(new_n658), .A2(new_n665), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n514), .A2(new_n518), .A3(new_n527), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n303), .ZN(new_n688));
  OAI21_X1  g502(.A(G472), .B1(new_n533), .B2(new_n688), .ZN(new_n689));
  OAI211_X1 g503(.A(new_n538), .B(new_n689), .C1(new_n554), .C2(new_n555), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n495), .A2(new_n621), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n686), .A2(new_n690), .A3(new_n691), .A4(new_n187), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n681), .B(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n638), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n692), .B1(new_n696), .B2(KEYINPUT40), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n300), .A2(new_n301), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n697), .B(new_n701), .C1(KEYINPUT40), .C2(new_n696), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  INV_X1    g517(.A(new_n622), .ZN(new_n704));
  INV_X1    g518(.A(new_n474), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n468), .A2(new_n455), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n705), .B1(new_n706), .B2(KEYINPUT92), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n385), .B1(new_n707), .B2(new_n470), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n483), .B1(new_n708), .B2(new_n480), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n476), .A2(KEYINPUT93), .A3(new_n481), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n490), .B1(new_n711), .B2(new_n464), .ZN(new_n712));
  INV_X1    g526(.A(new_n491), .ZN(new_n713));
  OAI21_X1  g527(.A(KEYINPUT33), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n489), .A2(new_n623), .A3(new_n491), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n704), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n648), .B(new_n681), .C1(new_n716), .C2(new_n629), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT102), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n626), .A2(new_n630), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(new_n720), .A3(new_n648), .A4(new_n681), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n679), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G146), .ZN(G48));
  NAND2_X1  g538(.A1(new_n428), .A2(new_n303), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(G469), .ZN(new_n726));
  INV_X1    g540(.A(new_n497), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n430), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n600), .A2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n634), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g545(.A(KEYINPUT41), .B(G113), .Z(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G15));
  NOR2_X1   g547(.A1(new_n652), .A2(new_n730), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n227), .ZN(G18));
  NOR3_X1   g549(.A1(new_n379), .A2(new_n493), .A3(new_n494), .ZN(new_n736));
  AND4_X1   g550(.A1(new_n556), .A2(new_n666), .A3(new_n736), .A4(new_n670), .ZN(new_n737));
  INV_X1    g551(.A(new_n728), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n610), .A2(new_n612), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G119), .ZN(G21));
  AND3_X1   g555(.A1(new_n610), .A2(new_n612), .A3(new_n691), .ZN(new_n742));
  NOR4_X1   g556(.A1(new_n639), .A2(new_n728), .A3(new_n360), .A4(new_n642), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G122), .ZN(G24));
  AOI21_X1  g559(.A(new_n642), .B1(new_n668), .B2(new_n664), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n718), .A2(new_n746), .A3(new_n721), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(new_n739), .A3(KEYINPUT103), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT103), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n718), .A2(new_n746), .A3(new_n721), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n610), .A2(new_n612), .A3(new_n738), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G125), .ZN(G27));
  NAND2_X1  g568(.A1(new_n698), .A2(new_n187), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n441), .A2(new_n727), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n755), .A2(new_n600), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT42), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n758), .A3(new_n722), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n607), .A2(new_n187), .A3(new_n609), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n554), .A2(KEYINPUT32), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n538), .A3(new_n547), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n497), .B1(new_n636), .B2(new_n438), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n760), .A2(new_n762), .A3(new_n599), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n718), .A2(new_n721), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT42), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n759), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G131), .ZN(G33));
  NAND2_X1  g582(.A1(new_n757), .A2(new_n683), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  NOR2_X1   g584(.A1(new_n716), .A2(new_n629), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n648), .ZN(new_n772));
  XOR2_X1   g586(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT43), .ZN(new_n775));
  OAI22_X1  g589(.A1(new_n771), .A2(new_n648), .B1(KEYINPUT106), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n777), .B(new_n642), .C1(new_n658), .C2(new_n665), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT44), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  OR3_X1    g595(.A1(new_n780), .A2(new_n781), .A3(new_n755), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT45), .B1(new_n435), .B2(new_n437), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n429), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n435), .A2(new_n437), .A3(KEYINPUT45), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n439), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n786), .A2(KEYINPUT46), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n430), .B1(new_n786), .B2(KEYINPUT46), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n727), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n694), .ZN(new_n791));
  XNOR2_X1  g605(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n792), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(new_n789), .B2(new_n694), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n782), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(new_n388), .ZN(G39));
  XNOR2_X1  g612(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n790), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n790), .A2(new_n799), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n755), .A2(new_n599), .A3(new_n556), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n722), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G140), .ZN(G42));
  NAND3_X1  g619(.A1(new_n599), .A2(new_n187), .A3(new_n499), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n806), .B(KEYINPUT108), .Z(new_n807));
  INV_X1    g621(.A(KEYINPUT49), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n726), .A2(new_n430), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT109), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n807), .B(new_n772), .C1(new_n808), .C2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(KEYINPUT110), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n690), .B1(new_n810), .B2(new_n808), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n812), .A2(new_n700), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT103), .B1(new_n747), .B2(new_n739), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n750), .A2(new_n751), .A3(new_n749), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n678), .B(new_n613), .C1(new_n722), .C2(new_n683), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT111), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n668), .A2(new_n664), .A3(new_n681), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n820), .B1(new_n821), .B2(new_n756), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n686), .A2(new_n763), .A3(KEYINPUT111), .A4(new_n681), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n742), .A3(new_n690), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n819), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n815), .B1(new_n818), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n753), .A2(KEYINPUT52), .A3(new_n819), .A4(new_n825), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n666), .A2(new_n670), .A3(new_n556), .A4(new_n637), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n495), .A2(new_n621), .A3(new_n681), .ZN(new_n831));
  OAI22_X1  g645(.A1(new_n750), .A2(new_n756), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n760), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(new_n766), .A3(new_n759), .A4(new_n769), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n737), .A2(new_n739), .B1(new_n742), .B2(new_n743), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n361), .B1(new_n631), .B2(new_n649), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(new_n302), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n837), .A2(new_n643), .B1(new_n601), .B2(new_n501), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n613), .B(new_n729), .C1(new_n633), .C2(new_n651), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n835), .A2(new_n838), .A3(new_n675), .A4(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n834), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT53), .B1(new_n829), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT112), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n829), .A2(KEYINPUT53), .A3(new_n841), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT113), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT54), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n819), .A2(new_n825), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT52), .B1(new_n848), .B2(new_n753), .ZN(new_n849));
  AND4_X1   g663(.A1(KEYINPUT52), .A2(new_n753), .A3(new_n819), .A4(new_n825), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n841), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n853), .A2(new_n854), .A3(new_n844), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n847), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n701), .A2(new_n187), .A3(new_n728), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n639), .A2(new_n642), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n777), .A2(new_n357), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT114), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT114), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n857), .A2(new_n863), .A3(new_n860), .ZN(new_n864));
  XOR2_X1   g678(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n865));
  NAND3_X1  g679(.A1(new_n862), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT116), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n862), .A2(new_n868), .A3(new_n864), .A4(new_n865), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n857), .A2(KEYINPUT50), .A3(new_n860), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT117), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n870), .A2(new_n871), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n867), .A2(new_n869), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n859), .A2(new_n755), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n810), .A2(new_n498), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n876), .B1(new_n802), .B2(new_n877), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n755), .A2(new_n356), .A3(new_n728), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n639), .A2(new_n690), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n881), .A2(new_n648), .A3(new_n719), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n879), .A2(new_n777), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n746), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n884), .A2(KEYINPUT118), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(KEYINPUT118), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n882), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n878), .A2(new_n887), .ZN(new_n888));
  OR3_X1    g702(.A1(new_n874), .A2(new_n875), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n875), .B1(new_n874), .B2(new_n888), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n883), .A2(new_n599), .A3(new_n762), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT48), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(KEYINPUT119), .A3(new_n892), .ZN(new_n893));
  XOR2_X1   g707(.A(KEYINPUT119), .B(KEYINPUT48), .Z(new_n894));
  OAI21_X1  g708(.A(new_n893), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  OAI221_X1 g709(.A(new_n354), .B1(new_n859), .B2(new_n751), .C1(new_n881), .C2(new_n632), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n889), .A2(new_n890), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT120), .B1(new_n856), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n899), .B1(G952), .B2(G953), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n856), .A2(new_n898), .A3(KEYINPUT120), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n814), .B1(new_n900), .B2(new_n901), .ZN(G75));
  NOR2_X1   g716(.A1(new_n307), .A2(G952), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n303), .B1(new_n853), .B2(new_n844), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT56), .B1(new_n905), .B2(G210), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n271), .A2(new_n273), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT121), .Z(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT55), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(new_n223), .Z(new_n910));
  OAI21_X1  g724(.A(new_n904), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(new_n906), .B2(new_n910), .ZN(G51));
  AND3_X1   g726(.A1(new_n905), .A2(new_n785), .A3(new_n784), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n829), .A2(KEYINPUT53), .A3(new_n841), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT54), .B1(new_n914), .B2(new_n842), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT122), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n855), .A3(new_n916), .ZN(new_n917));
  OAI211_X1 g731(.A(KEYINPUT122), .B(KEYINPUT54), .C1(new_n914), .C2(new_n842), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n439), .B(KEYINPUT57), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(KEYINPUT123), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n917), .A2(new_n922), .A3(new_n918), .A4(new_n919), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n428), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n913), .B1(new_n925), .B2(KEYINPUT124), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT124), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n924), .A2(new_n927), .A3(new_n428), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n903), .B1(new_n926), .B2(new_n928), .ZN(G54));
  NAND3_X1  g743(.A1(new_n905), .A2(KEYINPUT58), .A3(G475), .ZN(new_n930));
  INV_X1    g744(.A(new_n372), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n932), .A2(new_n933), .A3(new_n903), .ZN(G60));
  NAND2_X1  g748(.A1(new_n714), .A2(new_n715), .ZN(new_n935));
  XOR2_X1   g749(.A(KEYINPUT125), .B(KEYINPUT59), .Z(new_n936));
  NOR2_X1   g750(.A1(new_n442), .A2(new_n303), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n935), .B1(new_n856), .B2(new_n939), .ZN(new_n940));
  AND4_X1   g754(.A1(new_n935), .A2(new_n917), .A3(new_n918), .A4(new_n939), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n940), .A2(new_n903), .A3(new_n941), .ZN(G63));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT60), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n853), .B2(new_n844), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n663), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n946), .B(new_n904), .C1(new_n598), .C2(new_n945), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g762(.A(G953), .B1(new_n218), .B2(new_n359), .ZN(new_n949));
  INV_X1    g763(.A(new_n840), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n949), .B1(new_n950), .B2(G953), .ZN(new_n951));
  INV_X1    g765(.A(new_n908), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(G898), .B2(new_n307), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n951), .B(new_n953), .ZN(G69));
  AND2_X1   g768(.A1(new_n767), .A2(new_n769), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n804), .A2(new_n753), .A3(new_n819), .A4(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n742), .A2(new_n599), .A3(new_n762), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n793), .B2(new_n795), .ZN(new_n958));
  NOR4_X1   g772(.A1(new_n956), .A2(G953), .A3(new_n797), .A4(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n548), .A2(new_n529), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n365), .A2(new_n366), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT126), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n960), .B(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(G900), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n963), .B1(new_n964), .B2(new_n307), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n959), .A2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n967));
  AND2_X1   g781(.A1(G227), .A2(G900), .ZN(new_n968));
  OAI22_X1  g782(.A1(new_n966), .A2(new_n967), .B1(new_n307), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n702), .A2(new_n753), .A3(new_n819), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT62), .Z(new_n971));
  INV_X1    g785(.A(new_n797), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n631), .A2(new_n649), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n695), .A2(new_n973), .A3(new_n601), .A4(new_n760), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n971), .A2(new_n972), .A3(new_n804), .A4(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n963), .B1(new_n975), .B2(new_n307), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n966), .A2(new_n976), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n969), .B(new_n977), .Z(G72));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n975), .B2(new_n840), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n533), .ZN(new_n982));
  INV_X1    g796(.A(new_n540), .ZN(new_n983));
  NOR4_X1   g797(.A1(new_n956), .A2(new_n797), .A3(new_n840), .A4(new_n958), .ZN(new_n984));
  INV_X1    g798(.A(new_n980), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n982), .A2(new_n986), .A3(new_n904), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n983), .A2(new_n533), .A3(new_n985), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n987), .B1(new_n846), .B2(new_n988), .ZN(G57));
endmodule


