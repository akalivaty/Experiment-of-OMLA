//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n536, new_n537, new_n538, new_n539, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n550, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1111, new_n1112,
    new_n1113;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT66), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  OR4_X1    g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT67), .Z(new_n459));
  NAND2_X1  g034(.A1(new_n455), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND3_X1   g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n468));
  INV_X1    g043(.A(G113), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n469), .B2(new_n463), .ZN(new_n470));
  NAND3_X1  g045(.A1(KEYINPUT68), .A2(G113), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g047(.A(G2105), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(G101), .A3(G2104), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n476), .B(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  XNOR2_X1  g054(.A(KEYINPUT3), .B(G2104), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n480), .A2(G137), .A3(new_n475), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NOR3_X1   g057(.A1(new_n474), .A2(new_n479), .A3(new_n482), .ZN(G160));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n463), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI221_X1 g061(.A(new_n486), .B1(new_n485), .B2(new_n484), .C1(G112), .C2(new_n475), .ZN(new_n487));
  XOR2_X1   g062(.A(new_n487), .B(KEYINPUT71), .Z(new_n488));
  NAND2_X1  g063(.A1(new_n464), .A2(new_n466), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  AND3_X1   g066(.A1(new_n464), .A2(new_n466), .A3(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n488), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  XNOR2_X1  g069(.A(new_n494), .B(KEYINPUT72), .ZN(G162));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT73), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G114), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n497), .A2(new_n499), .A3(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n464), .A2(new_n466), .A3(G126), .A4(G2105), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n475), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n480), .A2(new_n508), .A3(G138), .A4(new_n475), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n505), .B1(new_n507), .B2(new_n509), .ZN(G164));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(KEYINPUT6), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT74), .A3(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(KEYINPUT6), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(G543), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G50), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT5), .B(G543), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n516), .A2(new_n517), .A3(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G88), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n525), .A2(new_n512), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n520), .A2(new_n524), .A3(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND2_X1  g103(.A1(new_n519), .A2(G51), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n523), .A2(G89), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n529), .A2(new_n530), .A3(new_n532), .A4(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  NAND2_X1  g110(.A1(new_n523), .A2(G90), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n519), .A2(G52), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(new_n512), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT5), .B(G543), .Z(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n519), .A2(G43), .B1(new_n545), .B2(G651), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n523), .A2(G81), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  NAND3_X1  g129(.A1(new_n519), .A2(KEYINPUT9), .A3(G53), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n523), .A2(G91), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n521), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n512), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n518), .B2(new_n560), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n555), .A2(new_n556), .A3(new_n558), .A4(new_n561), .ZN(G299));
  NAND2_X1  g137(.A1(new_n519), .A2(G49), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n523), .A2(G87), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(G288));
  AOI22_X1  g141(.A1(new_n521), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n512), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n516), .A2(G86), .A3(new_n517), .A4(new_n521), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n516), .A2(G48), .A3(G543), .A4(new_n517), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G305));
  XOR2_X1   g146(.A(KEYINPUT75), .B(G85), .Z(new_n572));
  AOI22_X1  g147(.A1(G47), .A2(new_n519), .B1(new_n523), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT76), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n575), .A2(new_n512), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(G290));
  NAND2_X1  g152(.A1(G301), .A2(G868), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n523), .A2(KEYINPUT10), .A3(G92), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT10), .ZN(new_n580));
  INV_X1    g155(.A(G92), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n522), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(G79), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G66), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n543), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n579), .A2(new_n582), .B1(G651), .B2(new_n585), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n518), .A2(KEYINPUT77), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n518), .A2(KEYINPUT77), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n587), .A2(G54), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(KEYINPUT78), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n586), .B2(new_n589), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n578), .B1(new_n594), .B2(G868), .ZN(G284));
  OAI21_X1  g170(.A(new_n578), .B1(new_n594), .B2(G868), .ZN(G321));
  INV_X1    g171(.A(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(G299), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(G168), .B2(new_n597), .ZN(G297));
  OAI21_X1  g174(.A(new_n598), .B1(G168), .B2(new_n597), .ZN(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n594), .B1(new_n601), .B2(G860), .ZN(G148));
  INV_X1    g177(.A(new_n548), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(new_n597), .ZN(new_n604));
  INV_X1    g179(.A(new_n594), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n604), .B1(new_n606), .B2(new_n597), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT79), .Z(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g184(.A1(new_n475), .A2(G2104), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n489), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT13), .Z(new_n613));
  INV_X1    g188(.A(G2100), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n490), .A2(G135), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n492), .A2(G123), .ZN(new_n617));
  NOR2_X1   g192(.A1(G99), .A2(G2105), .ZN(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(new_n475), .B2(G111), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n616), .B(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(G2096), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n613), .A2(new_n614), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n615), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT80), .Z(G156));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2430), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2435), .ZN(new_n627));
  XOR2_X1   g202(.A(G2427), .B(G2438), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2451), .B(G2454), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2443), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(G2446), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n632), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT82), .Z(new_n639));
  OAI211_X1 g214(.A(new_n639), .B(G14), .C1(new_n637), .C2(new_n636), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(G401));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT17), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2067), .B(G2678), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT83), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  AOI211_X1 g222(.A(new_n642), .B(new_n647), .C1(new_n643), .C2(new_n646), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT84), .ZN(new_n649));
  INV_X1    g224(.A(new_n643), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n650), .A2(new_n642), .A3(new_n645), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT18), .Z(new_n652));
  NAND3_X1  g227(.A1(new_n644), .A2(new_n642), .A3(new_n646), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n649), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(new_n621), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(new_n614), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G227));
  XNOR2_X1  g232(.A(G1971), .B(G1976), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  XOR2_X1   g234(.A(G1956), .B(G2474), .Z(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n659), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  AOI22_X1  g240(.A1(new_n663), .A2(KEYINPUT20), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n667), .A2(new_n659), .A3(new_n662), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n666), .B(new_n668), .C1(KEYINPUT20), .C2(new_n663), .ZN(new_n669));
  XOR2_X1   g244(.A(G1991), .B(G1996), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G229));
  MUX2_X1   g250(.A(G6), .B(G305), .S(G16), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT32), .ZN(new_n677));
  INV_X1    g252(.A(G1981), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(G16), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G23), .ZN(new_n681));
  INV_X1    g256(.A(G288), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n681), .B1(new_n682), .B2(new_n680), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT33), .Z(new_n684));
  OR2_X1    g259(.A1(new_n684), .A2(G1976), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n680), .A2(G22), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(G166), .B2(new_n680), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT86), .B(G1971), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n684), .A2(G1976), .ZN(new_n690));
  NAND4_X1  g265(.A1(new_n679), .A2(new_n685), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT34), .Z(new_n692));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G25), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n490), .A2(G131), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n492), .A2(G119), .ZN(new_n696));
  OR2_X1    g271(.A1(G95), .A2(G2105), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n697), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n694), .B1(new_n700), .B2(new_n693), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT35), .B(G1991), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n701), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G290), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(KEYINPUT85), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(KEYINPUT85), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n680), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G24), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n708), .B1(new_n680), .B2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G1986), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n692), .A2(new_n704), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT36), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n693), .A2(G32), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n490), .A2(G141), .B1(new_n492), .B2(G129), .ZN(new_n716));
  NAND3_X1  g291(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT26), .Z(new_n718));
  INV_X1    g293(.A(G105), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n716), .B(new_n718), .C1(new_n719), .C2(new_n610), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT91), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n715), .B1(new_n721), .B2(new_n693), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT92), .Z(new_n723));
  XOR2_X1   g298(.A(KEYINPUT27), .B(G1996), .Z(new_n724));
  INV_X1    g299(.A(G2084), .ZN(new_n725));
  AND2_X1   g300(.A1(KEYINPUT24), .A2(G34), .ZN(new_n726));
  NOR2_X1   g301(.A1(KEYINPUT24), .A2(G34), .ZN(new_n727));
  NOR3_X1   g302(.A1(new_n726), .A2(new_n727), .A3(G29), .ZN(new_n728));
  INV_X1    g303(.A(G160), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(G29), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n723), .A2(new_n724), .B1(new_n725), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n680), .A2(G5), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G171), .B2(new_n680), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT94), .Z(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n731), .B1(G1961), .B2(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT95), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n693), .A2(G26), .ZN(new_n738));
  OAI21_X1  g313(.A(G2104), .B1(new_n475), .B2(G116), .ZN(new_n739));
  INV_X1    g314(.A(G104), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(new_n475), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT87), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n490), .A2(G140), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n492), .A2(G128), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n738), .B1(new_n746), .B2(new_n693), .ZN(new_n747));
  MUX2_X1   g322(.A(new_n738), .B(new_n747), .S(KEYINPUT28), .Z(new_n748));
  XOR2_X1   g323(.A(KEYINPUT88), .B(G2067), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n680), .A2(G19), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n548), .B2(new_n680), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(G1341), .Z(new_n753));
  INV_X1    g328(.A(G28), .ZN(new_n754));
  AOI21_X1  g329(.A(G29), .B1(new_n754), .B2(KEYINPUT30), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(KEYINPUT30), .B2(new_n754), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n620), .B2(new_n693), .ZN(new_n757));
  NOR2_X1   g332(.A1(G164), .A2(new_n693), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G27), .B2(new_n693), .ZN(new_n759));
  INV_X1    g334(.A(G2078), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n757), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n750), .A2(new_n753), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT93), .B(G11), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT31), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n730), .A2(new_n725), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(KEYINPUT90), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(KEYINPUT90), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n766), .B(new_n767), .C1(new_n760), .C2(new_n759), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n762), .A2(new_n764), .A3(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(G29), .A2(G33), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n490), .A2(G139), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT25), .Z(new_n773));
  AOI22_X1  g348(.A1(new_n480), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT89), .Z(new_n775));
  OAI211_X1 g350(.A(new_n771), .B(new_n773), .C1(new_n775), .C2(new_n475), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n770), .B1(new_n776), .B2(new_n693), .ZN(new_n777));
  INV_X1    g352(.A(G2072), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(G168), .A2(G16), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G16), .B2(G21), .ZN(new_n781));
  INV_X1    g356(.A(G1966), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n783), .B(new_n784), .C1(new_n777), .C2(new_n778), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT96), .B(G1956), .Z(new_n786));
  AND2_X1   g361(.A1(new_n680), .A2(G20), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G299), .B2(G16), .ZN(new_n788));
  MUX2_X1   g363(.A(new_n787), .B(new_n788), .S(KEYINPUT23), .Z(new_n789));
  AOI21_X1  g364(.A(new_n785), .B1(new_n786), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n693), .A2(G35), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G162), .B2(new_n693), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT29), .B(G2090), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n769), .A2(new_n779), .A3(new_n790), .A4(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n594), .A2(new_n680), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G4), .B2(new_n680), .ZN(new_n797));
  INV_X1    g372(.A(G1348), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  OAI221_X1 g375(.A(new_n800), .B1(new_n786), .B2(new_n789), .C1(new_n723), .C2(new_n724), .ZN(new_n801));
  NOR4_X1   g376(.A1(new_n737), .A2(new_n795), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G1961), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n734), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n714), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(G311));
  XNOR2_X1  g381(.A(new_n805), .B(KEYINPUT97), .ZN(G150));
  NAND2_X1  g382(.A1(new_n519), .A2(G55), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT98), .B(G93), .Z(new_n810));
  OAI221_X1 g385(.A(new_n808), .B1(new_n512), .B2(new_n809), .C1(new_n522), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G860), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT37), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n594), .A2(G559), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT38), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n811), .B(new_n548), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT39), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n815), .B(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n813), .B1(new_n818), .B2(G860), .ZN(G145));
  NAND2_X1  g394(.A1(new_n490), .A2(G142), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n820), .A2(KEYINPUT99), .B1(G130), .B2(new_n492), .ZN(new_n821));
  NOR2_X1   g396(.A1(G106), .A2(G2105), .ZN(new_n822));
  OAI21_X1  g397(.A(G2104), .B1(new_n475), .B2(G118), .ZN(new_n823));
  OAI221_X1 g398(.A(new_n821), .B1(KEYINPUT99), .B2(new_n820), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(new_n700), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(new_n776), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n729), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n745), .B(KEYINPUT100), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n612), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n721), .B(G164), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n827), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(G162), .B(new_n620), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT101), .B(G37), .Z(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g412(.A1(new_n811), .A2(new_n597), .ZN(new_n838));
  XNOR2_X1  g413(.A(G303), .B(G288), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G305), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n705), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(KEYINPUT102), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT42), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n606), .B(new_n816), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n590), .B(G299), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT41), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n846), .B2(new_n845), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n844), .B(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n838), .B1(new_n850), .B2(new_n597), .ZN(G295));
  OAI21_X1  g426(.A(new_n838), .B1(new_n850), .B2(new_n597), .ZN(G331));
  INV_X1    g427(.A(KEYINPUT44), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n816), .B(G301), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G286), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n846), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n847), .B2(new_n855), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(new_n841), .ZN(new_n858));
  INV_X1    g433(.A(G37), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n856), .B(new_n842), .C1(new_n847), .C2(new_n855), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT43), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n858), .A2(KEYINPUT43), .A3(new_n835), .A4(new_n860), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n853), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n861), .A2(KEYINPUT43), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n858), .A2(new_n862), .A3(new_n835), .A4(new_n860), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT44), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n865), .A2(new_n868), .A3(KEYINPUT103), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(G397));
  NAND2_X1  g448(.A1(new_n705), .A2(new_n711), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT104), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT45), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(G164), .B2(G1384), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n473), .A2(G40), .A3(new_n478), .A4(new_n481), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT48), .ZN(new_n881));
  INV_X1    g456(.A(new_n879), .ZN(new_n882));
  INV_X1    g457(.A(G1996), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n721), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n721), .A2(new_n883), .ZN(new_n885));
  INV_X1    g460(.A(G2067), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n745), .B(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n700), .A2(new_n703), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n699), .A2(new_n702), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n881), .B1(new_n882), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n882), .B1(new_n887), .B2(new_n721), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n879), .A2(KEYINPUT46), .A3(new_n883), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT46), .B1(new_n879), .B2(new_n883), .ZN(new_n895));
  NOR3_X1   g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n896), .B(KEYINPUT47), .Z(new_n897));
  INV_X1    g472(.A(new_n890), .ZN(new_n898));
  OAI22_X1  g473(.A1(new_n888), .A2(new_n898), .B1(G2067), .B2(new_n745), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n879), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n892), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n507), .A2(new_n509), .ZN(new_n902));
  AOI22_X1  g477(.A1(new_n492), .A2(G126), .B1(new_n500), .B2(new_n502), .ZN(new_n903));
  AOI21_X1  g478(.A(G1384), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI211_X1 g481(.A(KEYINPUT105), .B(G1384), .C1(new_n902), .C2(new_n903), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n876), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n878), .B1(new_n904), .B2(KEYINPUT45), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT50), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(new_n906), .B2(new_n907), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n902), .A2(new_n903), .ZN(new_n914));
  INV_X1    g489(.A(G1384), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n878), .B1(new_n916), .B2(KEYINPUT50), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  OAI22_X1  g493(.A1(new_n911), .A2(G1966), .B1(G2084), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(G8), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n920), .A2(G286), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n569), .A2(new_n570), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT108), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n568), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(KEYINPUT109), .A3(G1981), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT111), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT49), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT108), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT108), .B1(new_n569), .B2(new_n570), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n678), .B1(new_n933), .B2(new_n568), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n568), .A2(new_n678), .A3(new_n569), .A4(new_n570), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n935), .A2(KEYINPUT109), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n927), .B(new_n930), .C1(new_n934), .C2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n928), .B1(KEYINPUT110), .B2(new_n929), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n927), .B(new_n938), .C1(new_n934), .C2(new_n936), .ZN(new_n941));
  INV_X1    g516(.A(new_n878), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(new_n906), .B2(new_n907), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(G8), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n940), .A2(new_n941), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G1976), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT52), .B1(G288), .B2(new_n947), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n945), .B(new_n948), .C1(new_n947), .C2(G288), .ZN(new_n949));
  NOR2_X1   g524(.A1(G288), .A2(new_n947), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT52), .B1(new_n944), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n946), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n946), .A2(new_n949), .A3(KEYINPUT112), .A4(new_n951), .ZN(new_n955));
  INV_X1    g530(.A(G8), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n910), .A2(new_n877), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n957), .A2(G1971), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G2090), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n913), .A2(new_n960), .A3(new_n917), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n956), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(G303), .A2(G8), .ZN(new_n963));
  XOR2_X1   g538(.A(KEYINPUT106), .B(KEYINPUT55), .Z(new_n964));
  XNOR2_X1  g539(.A(new_n963), .B(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  OR2_X1    g541(.A1(new_n962), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n921), .A2(new_n954), .A3(new_n955), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT63), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n970), .B1(new_n962), .B2(new_n966), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n962), .A2(new_n970), .A3(new_n966), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n952), .A2(KEYINPUT116), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT116), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n946), .A2(new_n949), .A3(new_n976), .A4(new_n951), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n920), .A2(KEYINPUT63), .A3(G286), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n906), .A2(new_n907), .A3(new_n912), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n878), .B1(new_n904), .B2(new_n912), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n980), .A2(G2090), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(G8), .B1(new_n983), .B2(new_n958), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n965), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n974), .A2(new_n978), .A3(new_n979), .A4(new_n985), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n954), .A2(new_n955), .ZN(new_n987));
  INV_X1    g562(.A(new_n973), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(new_n971), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n682), .A2(new_n947), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT114), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n946), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n935), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT115), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n944), .A2(KEYINPUT113), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n993), .A2(new_n997), .A3(new_n935), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n944), .A2(KEYINPUT113), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n995), .A2(new_n996), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n969), .A2(new_n986), .A3(new_n990), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT117), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI22_X1  g578(.A1(KEYINPUT63), .A2(new_n968), .B1(new_n987), .B2(new_n989), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1004), .A2(KEYINPUT117), .A3(new_n986), .A4(new_n1000), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(G168), .A2(new_n956), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n919), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1007), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n920), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1009), .B1(new_n920), .B2(new_n1010), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1008), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT123), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1008), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n920), .A2(new_n1010), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT51), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1016), .B1(new_n1018), .B2(new_n1011), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT123), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n911), .A2(KEYINPUT53), .A3(new_n760), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n957), .A2(new_n760), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n1023), .A2(new_n1024), .B1(new_n918), .B2(new_n803), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(G171), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1015), .A2(new_n1021), .A3(KEYINPUT62), .A4(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1027), .A2(KEYINPUT62), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1348), .B1(new_n913), .B2(new_n917), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n886), .B(new_n942), .C1(new_n906), .C2(new_n907), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n594), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(G299), .B(KEYINPUT57), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1036), .B(new_n778), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n910), .A2(new_n877), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT119), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n910), .A2(new_n877), .A3(new_n1040), .A4(new_n1037), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n916), .A2(KEYINPUT105), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n904), .A2(new_n905), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(KEYINPUT50), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(G1956), .B1(new_n1045), .B2(new_n981), .ZN(new_n1046));
  OAI211_X1 g621(.A(KEYINPUT120), .B(new_n1035), .C1(new_n1042), .C2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1956), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(new_n980), .B2(new_n982), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1050), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT120), .B1(new_n1051), .B2(new_n1035), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1034), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1035), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1050), .A2(new_n1054), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT60), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT122), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT50), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1059));
  INV_X1    g634(.A(new_n917), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n798), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1057), .B1(new_n1061), .B2(new_n1032), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1058), .B(new_n1034), .C1(new_n1062), .C2(new_n594), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT60), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n605), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1058), .B1(new_n1066), .B2(new_n1034), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1057), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1034), .B1(new_n1062), .B2(new_n594), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT122), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1070), .A2(KEYINPUT60), .A3(new_n1063), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1055), .A2(KEYINPUT61), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT58), .B(G1341), .Z(new_n1075));
  AOI22_X1  g650(.A1(new_n957), .A2(new_n883), .B1(new_n943), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(new_n603), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1077), .B(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1035), .B1(new_n1042), .B2(new_n1046), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n1055), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT61), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1080), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI211_X1 g659(.A(KEYINPUT121), .B(KEYINPUT61), .C1(new_n1081), .C2(new_n1055), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1074), .B(new_n1079), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1056), .B1(new_n1072), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1025), .B1(new_n1024), .B2(new_n1023), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1088), .A2(G171), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT54), .B1(new_n1089), .B2(new_n1027), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1088), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT125), .B1(new_n1088), .B2(G171), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1022), .A2(G301), .A3(new_n1025), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1090), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1030), .B1(new_n1087), .B2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1019), .B(KEYINPUT123), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1029), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n978), .A2(new_n974), .A3(new_n985), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1100), .B(KEYINPUT124), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1006), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n875), .B1(G1986), .B2(G290), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n882), .B1(new_n1103), .B2(new_n891), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n901), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT126), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT126), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1107), .B(new_n901), .C1(new_n1102), .C2(new_n1104), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1108), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g684(.A1(new_n866), .A2(new_n867), .ZN(new_n1111));
  NOR2_X1   g685(.A1(G229), .A2(new_n461), .ZN(new_n1112));
  NOR2_X1   g686(.A1(G401), .A2(G227), .ZN(new_n1113));
  NAND4_X1  g687(.A1(new_n1111), .A2(new_n836), .A3(new_n1112), .A4(new_n1113), .ZN(G225));
  XNOR2_X1  g688(.A(G225), .B(KEYINPUT127), .ZN(G308));
endmodule


