//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT83), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G122), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT3), .B1(new_n192), .B2(G107), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n194));
  INV_X1    g008(.A(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G104), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n192), .A2(G107), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n193), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT77), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n199), .A3(G101), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n193), .A2(new_n196), .A3(new_n201), .A4(new_n197), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT4), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n198), .A2(new_n199), .A3(KEYINPUT4), .A4(G101), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT2), .A2(G113), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT65), .B1(KEYINPUT2), .B2(G113), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NOR3_X1   g023(.A1(KEYINPUT65), .A2(KEYINPUT2), .A3(G113), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n207), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G119), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G116), .ZN(new_n213));
  INV_X1    g027(.A(G116), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G119), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n211), .B(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n206), .A2(new_n217), .ZN(new_n218));
  OR2_X1    g032(.A1(new_n213), .A2(KEYINPUT5), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT5), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(G113), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT81), .ZN(new_n222));
  OR2_X1    g036(.A1(new_n211), .A2(new_n216), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n195), .A2(G104), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n192), .A2(G107), .ZN(new_n225));
  OAI21_X1  g039(.A(G101), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n202), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT81), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n219), .A2(new_n228), .A3(new_n220), .A4(G113), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n222), .A2(new_n223), .A3(new_n227), .A4(new_n229), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n218), .A2(KEYINPUT82), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT82), .B1(new_n218), .B2(new_n230), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n189), .B(new_n191), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT6), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n218), .A2(new_n230), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n218), .A2(KEYINPUT82), .A3(new_n230), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n240), .A2(new_n189), .A3(KEYINPUT6), .A4(new_n191), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n218), .A2(new_n190), .A3(new_n230), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n235), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G146), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G143), .ZN(new_n245));
  INV_X1    g059(.A(G143), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G146), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n245), .A2(new_n247), .A3(new_n249), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G125), .ZN(new_n255));
  INV_X1    g069(.A(G128), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(KEYINPUT1), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(new_n245), .A3(new_n247), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n244), .A3(G143), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n246), .B(G146), .C1(new_n256), .C2(KEYINPUT1), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n255), .B1(G125), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G953), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G224), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n265), .B(KEYINPUT84), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n263), .B(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n243), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G902), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT7), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n263), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT85), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n223), .A2(new_n221), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n227), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n190), .B(KEYINPUT8), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n222), .A2(new_n223), .A3(new_n229), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n277), .B(new_n278), .C1(new_n279), .C2(new_n227), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n263), .A2(KEYINPUT85), .A3(new_n272), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n275), .A2(new_n280), .A3(new_n242), .A4(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n263), .A2(new_n272), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n270), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n269), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(G210), .B1(G237), .B2(G902), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n269), .A2(new_n287), .A3(new_n285), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n188), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OR2_X1    g105(.A1(KEYINPUT64), .A2(G134), .ZN(new_n292));
  NAND2_X1  g106(.A1(KEYINPUT64), .A2(G134), .ZN(new_n293));
  INV_X1    g107(.A(G137), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n292), .A2(new_n293), .B1(KEYINPUT11), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(KEYINPUT11), .A3(G134), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT11), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G137), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n295), .A2(new_n299), .A3(G131), .ZN(new_n300));
  INV_X1    g114(.A(G131), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n296), .A2(new_n298), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n294), .A2(KEYINPUT11), .ZN(new_n303));
  AND2_X1   g117(.A1(KEYINPUT64), .A2(G134), .ZN(new_n304));
  NOR2_X1   g118(.A1(KEYINPUT64), .A2(G134), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n301), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n300), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n206), .A2(new_n254), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n261), .A2(new_n226), .A3(new_n202), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT10), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT10), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n227), .A2(new_n313), .A3(new_n261), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT79), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n310), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n316), .B1(new_n310), .B2(new_n315), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n309), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT80), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n310), .A2(new_n315), .A3(new_n308), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT80), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n322), .B(new_n309), .C1(new_n317), .C2(new_n318), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n320), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(G110), .B(G140), .ZN(new_n325));
  INV_X1    g139(.A(G227), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n326), .A2(G953), .ZN(new_n327));
  XOR2_X1   g141(.A(new_n325), .B(new_n327), .Z(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n311), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n202), .A2(new_n226), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n262), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n262), .A2(new_n333), .A3(new_n331), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n309), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT12), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT12), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n340), .A3(new_n309), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n321), .A3(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n342), .A2(new_n329), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(G902), .B1(new_n330), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G469), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n346), .A2(new_n270), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n320), .A2(new_n328), .A3(new_n321), .A4(new_n323), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n342), .A2(new_n329), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(G469), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n347), .A2(new_n349), .A3(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT91), .B1(new_n256), .B2(G143), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT91), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(new_n246), .A3(G128), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT13), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n354), .A2(new_n356), .A3(KEYINPUT13), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n256), .A2(G143), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G134), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n357), .B(new_n361), .C1(new_n305), .C2(new_n304), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT89), .ZN(new_n365));
  INV_X1    g179(.A(G122), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(KEYINPUT89), .A2(G122), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n214), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n366), .A2(G116), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT90), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n368), .ZN(new_n372));
  NOR2_X1   g186(.A1(KEYINPUT89), .A2(G122), .ZN(new_n373));
  OAI21_X1  g187(.A(G116), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT90), .ZN(new_n375));
  INV_X1    g189(.A(new_n370), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n371), .A2(new_n195), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n195), .B1(new_n371), .B2(new_n377), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n363), .B(new_n364), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  XOR2_X1   g194(.A(new_n370), .B(KEYINPUT14), .Z(new_n381));
  OAI21_X1  g195(.A(G107), .B1(new_n381), .B2(new_n369), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n357), .A2(new_n361), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n292), .A3(new_n293), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n364), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n371), .A2(new_n195), .A3(new_n377), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n380), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT9), .B(G234), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(KEYINPUT76), .ZN(new_n390));
  XOR2_X1   g204(.A(KEYINPUT70), .B(G217), .Z(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n390), .A2(G953), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n388), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n380), .A2(new_n387), .A3(new_n393), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(KEYINPUT92), .A3(new_n396), .ZN(new_n397));
  OR3_X1    g211(.A1(new_n388), .A2(KEYINPUT92), .A3(new_n394), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(new_n270), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT93), .ZN(new_n400));
  INV_X1    g214(.A(G478), .ZN(new_n401));
  OR2_X1    g215(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n402));
  NAND2_X1  g216(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT93), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n397), .A2(new_n398), .A3(new_n405), .A4(new_n270), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n400), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  OR2_X1    g221(.A1(new_n399), .A2(new_n404), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n264), .A2(G952), .ZN(new_n410));
  INV_X1    g224(.A(G234), .ZN(new_n411));
  INV_X1    g225(.A(G237), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT21), .B(G898), .ZN(new_n415));
  XOR2_X1   g229(.A(new_n415), .B(KEYINPUT95), .Z(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  AOI211_X1 g231(.A(new_n270), .B(new_n264), .C1(G234), .C2(G237), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n414), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G475), .ZN(new_n420));
  INV_X1    g234(.A(G125), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n421), .A2(KEYINPUT16), .A3(G140), .ZN(new_n422));
  XNOR2_X1  g236(.A(G125), .B(G140), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n422), .B1(new_n423), .B2(KEYINPUT16), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(G146), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(KEYINPUT86), .A2(G143), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n412), .A2(new_n264), .A3(G214), .ZN(new_n429));
  NAND2_X1  g243(.A1(KEYINPUT86), .A2(G143), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n427), .A2(G214), .A3(new_n412), .A4(new_n264), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n431), .A2(KEYINPUT17), .A3(G131), .A4(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n432), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(G131), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n426), .B(new_n433), .C1(new_n436), .C2(KEYINPUT17), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n423), .A2(new_n244), .ZN(new_n438));
  OR2_X1    g252(.A1(G125), .A2(G140), .ZN(new_n439));
  NAND2_X1  g253(.A1(G125), .A2(G140), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(G146), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(KEYINPUT87), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT18), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n434), .B1(new_n444), .B2(new_n301), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n438), .A2(KEYINPUT87), .A3(new_n441), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n431), .A2(KEYINPUT18), .A3(G131), .A4(new_n432), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n443), .A2(new_n445), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT88), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n446), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n451), .A2(new_n442), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n452), .A2(KEYINPUT88), .A3(new_n445), .A4(new_n447), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G113), .B(G122), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(new_n192), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n437), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n424), .A2(G146), .ZN(new_n458));
  XOR2_X1   g272(.A(new_n423), .B(KEYINPUT19), .Z(new_n459));
  OAI21_X1  g273(.A(new_n458), .B1(new_n459), .B2(G146), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(new_n435), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n456), .B1(new_n454), .B2(new_n462), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n420), .B(new_n270), .C1(new_n457), .C2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT20), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n456), .B1(new_n437), .B2(new_n454), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n270), .B1(new_n457), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G475), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n437), .A2(new_n454), .A3(new_n456), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n461), .B1(new_n450), .B2(new_n453), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n470), .B1(new_n456), .B2(new_n471), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n472), .A2(KEYINPUT20), .A3(new_n420), .A4(new_n270), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n466), .A2(new_n469), .A3(new_n473), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n409), .A2(new_n419), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(G221), .B1(new_n390), .B2(G902), .ZN(new_n476));
  AND4_X1   g290(.A1(new_n291), .A2(new_n353), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT32), .ZN(new_n478));
  OAI21_X1  g292(.A(G131), .B1(new_n295), .B2(new_n299), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n306), .A2(new_n301), .A3(new_n296), .A4(new_n298), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n479), .A2(new_n480), .B1(new_n252), .B2(new_n253), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n294), .B1(new_n304), .B2(new_n305), .ZN(new_n482));
  NAND2_X1  g296(.A1(G134), .A2(G137), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(G131), .A3(new_n483), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n480), .A2(new_n261), .A3(new_n484), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n481), .A2(new_n485), .A3(KEYINPUT30), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT30), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n254), .B1(new_n300), .B2(new_n307), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n480), .A2(new_n261), .A3(new_n484), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n217), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n216), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n211), .B(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n488), .A2(new_n493), .A3(new_n489), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(G101), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n412), .A2(new_n264), .A3(G210), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n496), .B(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(KEYINPUT66), .A2(KEYINPUT31), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n491), .A2(new_n494), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(KEYINPUT66), .A2(KEYINPUT31), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n494), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT30), .B1(new_n481), .B2(new_n485), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n488), .A2(new_n487), .A3(new_n489), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n503), .B1(new_n506), .B2(new_n217), .ZN(new_n507));
  INV_X1    g321(.A(new_n501), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n507), .A2(new_n498), .A3(new_n508), .A4(new_n499), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT28), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n494), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n217), .B1(new_n481), .B2(new_n485), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT67), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT67), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n514), .B(new_n217), .C1(new_n481), .C2(new_n485), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n503), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n511), .B1(new_n516), .B2(new_n510), .ZN(new_n517));
  INV_X1    g331(.A(new_n498), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n502), .A2(new_n509), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(G472), .A2(G902), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n478), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n517), .A2(new_n498), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n507), .A2(new_n518), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT29), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT68), .ZN(new_n527));
  INV_X1    g341(.A(new_n511), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n510), .B1(new_n512), .B2(new_n494), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n498), .A2(KEYINPUT29), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n527), .B(new_n270), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n528), .A2(new_n529), .A3(new_n531), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT68), .B1(new_n533), .B2(G902), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(G472), .B1(new_n526), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT69), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n502), .A2(new_n509), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n517), .A2(new_n518), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n521), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n537), .B1(new_n540), .B2(KEYINPUT32), .ZN(new_n541));
  NOR4_X1   g355(.A1(new_n519), .A2(KEYINPUT69), .A3(new_n478), .A4(new_n521), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n522), .B(new_n536), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  OR3_X1    g357(.A1(new_n256), .A2(KEYINPUT71), .A3(G119), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT71), .B1(new_n256), .B2(G119), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n544), .A2(new_n545), .B1(G119), .B2(new_n256), .ZN(new_n546));
  XOR2_X1   g360(.A(KEYINPUT24), .B(G110), .Z(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT72), .B1(new_n212), .B2(G128), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT23), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT23), .ZN(new_n551));
  OAI211_X1 g365(.A(KEYINPUT72), .B(new_n551), .C1(new_n212), .C2(G128), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n550), .B(new_n552), .C1(G119), .C2(new_n256), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G110), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n425), .A2(new_n548), .A3(new_n554), .ZN(new_n555));
  OAI22_X1  g369(.A1(new_n553), .A2(G110), .B1(new_n546), .B2(new_n547), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(new_n438), .A3(new_n458), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n264), .A2(G221), .A3(G234), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT22), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(G137), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n555), .A2(new_n557), .A3(new_n561), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n270), .A3(new_n564), .ZN(new_n565));
  OR2_X1    g379(.A1(new_n565), .A2(KEYINPUT25), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(KEYINPUT25), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n392), .B1(G234), .B2(new_n270), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT74), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n563), .A2(new_n564), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n568), .A2(G902), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n572), .B(KEYINPUT73), .Z(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n569), .A2(new_n570), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n570), .B1(new_n569), .B2(new_n574), .ZN(new_n576));
  OR2_X1    g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n543), .A2(KEYINPUT75), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT75), .B1(new_n543), .B2(new_n577), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n477), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(G101), .ZN(G3));
  INV_X1    g395(.A(new_n419), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n466), .A2(new_n469), .A3(new_n473), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n400), .A2(new_n401), .A3(new_n406), .ZN(new_n584));
  XOR2_X1   g398(.A(KEYINPUT96), .B(KEYINPUT33), .Z(new_n585));
  NAND3_X1  g399(.A1(new_n397), .A2(new_n398), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n395), .A2(KEYINPUT33), .A3(new_n396), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(G478), .A3(new_n270), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n583), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n291), .A2(KEYINPUT97), .A3(new_n582), .A4(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT97), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n287), .B1(new_n269), .B2(new_n285), .ZN(new_n593));
  AOI211_X1 g407(.A(new_n288), .B(new_n284), .C1(new_n243), .C2(new_n268), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n187), .B(new_n582), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n589), .A2(new_n584), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n474), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n592), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n591), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n538), .A2(new_n539), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n270), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n540), .B1(new_n601), .B2(G472), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n353), .A2(new_n476), .A3(new_n577), .A4(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT34), .B(G104), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G6));
  NAND2_X1  g420(.A1(new_n409), .A2(new_n583), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n607), .A2(KEYINPUT98), .A3(new_n419), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n289), .A2(new_n290), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n187), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n474), .B1(new_n408), .B2(new_n407), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n611), .B1(new_n612), .B2(new_n582), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n608), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n353), .A2(new_n476), .A3(new_n577), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n614), .A2(new_n602), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT35), .B(G107), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G9));
  NOR2_X1   g432(.A1(new_n562), .A2(KEYINPUT36), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(new_n558), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n573), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n569), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n477), .A2(new_n602), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n623), .B(KEYINPUT37), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G110), .ZN(G12));
  INV_X1    g439(.A(new_n622), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n600), .A2(KEYINPUT32), .A3(new_n520), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT69), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n540), .A2(new_n537), .A3(KEYINPUT32), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n524), .B1(new_n517), .B2(new_n498), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n534), .B(new_n532), .C1(new_n631), .C2(KEYINPUT29), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n600), .A2(new_n520), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n632), .A2(G472), .B1(new_n633), .B2(new_n478), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n626), .B1(new_n630), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n476), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n348), .B1(new_n345), .B2(new_n346), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n636), .B1(new_n637), .B2(new_n352), .ZN(new_n638));
  INV_X1    g452(.A(G900), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n418), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n413), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n607), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n635), .A2(new_n638), .A3(new_n291), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G128), .ZN(G30));
  NAND3_X1  g459(.A1(new_n409), .A2(new_n187), .A3(new_n474), .ZN(new_n646));
  INV_X1    g460(.A(new_n512), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n503), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n270), .B1(new_n649), .B2(new_n498), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n507), .A2(new_n518), .ZN(new_n651));
  OAI21_X1  g465(.A(G472), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n630), .A2(new_n522), .A3(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n641), .B(KEYINPUT39), .Z(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n638), .A2(new_n656), .ZN(new_n657));
  AOI211_X1 g471(.A(new_n646), .B(new_n654), .C1(KEYINPUT40), .C2(new_n657), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n657), .A2(KEYINPUT40), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n609), .B(KEYINPUT38), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n658), .A2(new_n626), .A3(new_n659), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G143), .ZN(G45));
  AND3_X1   g476(.A1(new_n596), .A2(new_n474), .A3(new_n641), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n635), .A2(new_n638), .A3(new_n291), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G146), .ZN(G48));
  NOR2_X1   g479(.A1(new_n575), .A2(new_n576), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n630), .B2(new_n634), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n343), .B1(new_n324), .B2(new_n329), .ZN(new_n668));
  OAI21_X1  g482(.A(G469), .B1(new_n668), .B2(G902), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n347), .A2(new_n669), .A3(new_n476), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n591), .A2(new_n598), .A3(new_n667), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT99), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT41), .B(G113), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G15));
  NOR2_X1   g489(.A1(new_n608), .A2(new_n613), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n676), .A2(new_n291), .A3(new_n667), .A4(new_n671), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G116), .ZN(G18));
  NOR2_X1   g492(.A1(new_n610), .A2(new_n670), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n475), .A3(new_n635), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G119), .ZN(G21));
  NAND2_X1  g495(.A1(new_n601), .A2(G472), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n569), .A2(new_n574), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n530), .A2(new_n518), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n538), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n520), .B(KEYINPUT100), .Z(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n682), .A2(new_n683), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n670), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n595), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n689), .A2(new_n409), .A3(new_n474), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G122), .ZN(G24));
  AND3_X1   g506(.A1(new_n682), .A2(new_n622), .A3(new_n687), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n671), .A2(new_n663), .A3(new_n291), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G125), .ZN(G27));
  INV_X1    g509(.A(KEYINPUT42), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n351), .A2(KEYINPUT101), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n342), .A2(new_n698), .A3(new_n329), .ZN(new_n699));
  AND4_X1   g513(.A1(G469), .A2(new_n697), .A3(new_n350), .A4(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n637), .A2(new_n701), .ZN(new_n702));
  NOR4_X1   g516(.A1(new_n593), .A2(new_n594), .A3(new_n188), .A4(new_n636), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n667), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n596), .A2(new_n474), .A3(new_n641), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n696), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n536), .A2(new_n522), .A3(new_n627), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n683), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT102), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT102), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n707), .A2(new_n710), .A3(new_n683), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n668), .A2(G469), .A3(G902), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n713), .A2(new_n700), .A3(new_n348), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n289), .A2(new_n187), .A3(new_n290), .A4(new_n476), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n714), .A2(new_n715), .A3(new_n705), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n712), .A2(new_n716), .A3(KEYINPUT42), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n706), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G131), .ZN(G33));
  NAND4_X1  g533(.A1(new_n667), .A2(new_n643), .A3(new_n702), .A4(new_n703), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G134), .ZN(G36));
  NOR2_X1   g535(.A1(new_n593), .A2(new_n594), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n187), .ZN(new_n723));
  AOI211_X1 g537(.A(KEYINPUT43), .B(new_n474), .C1(new_n589), .C2(new_n584), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n474), .B(KEYINPUT104), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n596), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n724), .B1(new_n726), .B2(KEYINPUT43), .ZN(new_n727));
  INV_X1    g541(.A(new_n602), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n727), .A2(new_n728), .A3(new_n622), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n723), .B1(new_n729), .B2(KEYINPUT44), .ZN(new_n730));
  XOR2_X1   g544(.A(new_n730), .B(KEYINPUT105), .Z(new_n731));
  AND3_X1   g545(.A1(new_n697), .A2(new_n350), .A3(new_n699), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n732), .A2(KEYINPUT103), .A3(KEYINPUT45), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT103), .B1(new_n732), .B2(KEYINPUT45), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT45), .B1(new_n350), .B2(new_n351), .ZN(new_n735));
  OR4_X1    g549(.A1(new_n346), .A2(new_n733), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n349), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT46), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n736), .A2(KEYINPUT46), .A3(new_n349), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n347), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n476), .A3(new_n656), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n743));
  INV_X1    g557(.A(new_n729), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n731), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G137), .ZN(G39));
  NAND2_X1  g561(.A1(new_n741), .A2(new_n476), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT47), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n741), .A2(KEYINPUT47), .A3(new_n476), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR4_X1   g566(.A1(new_n723), .A2(new_n543), .A3(new_n705), .A4(new_n577), .ZN(new_n753));
  XOR2_X1   g567(.A(new_n753), .B(KEYINPUT106), .Z(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G140), .ZN(G42));
  INV_X1    g570(.A(KEYINPUT54), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n644), .A2(new_n694), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT108), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n653), .A2(new_n626), .A3(new_n702), .ZN(new_n761));
  NOR4_X1   g575(.A1(new_n722), .A2(new_n646), .A3(new_n636), .A4(new_n642), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n644), .A2(new_n764), .A3(new_n694), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n759), .A2(new_n664), .A3(new_n763), .A4(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n664), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n758), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n761), .A2(new_n762), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n760), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n769), .B1(new_n758), .B2(KEYINPUT108), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(KEYINPUT109), .A3(new_n763), .A4(new_n765), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n768), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT107), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n590), .A2(new_n612), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n603), .A2(new_n595), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n667), .B(KEYINPUT75), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n779), .B1(new_n780), .B2(new_n477), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n667), .A2(new_n671), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n671), .A2(new_n291), .A3(new_n475), .ZN(new_n783));
  AOI22_X1  g597(.A1(new_n614), .A2(new_n782), .B1(new_n783), .B2(new_n635), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n672), .A2(new_n691), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n781), .A2(new_n623), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n682), .A2(new_n687), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n703), .A2(new_n663), .A3(new_n787), .A4(new_n702), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n703), .A2(new_n353), .A3(new_n543), .A4(new_n641), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n583), .A2(new_n408), .A3(new_n407), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n622), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n718), .A2(new_n792), .A3(new_n720), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n777), .B1(new_n786), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n677), .A2(new_n672), .A3(new_n680), .A4(new_n691), .ZN(new_n795));
  INV_X1    g609(.A(new_n778), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n615), .A2(new_n796), .A3(new_n690), .A4(new_n602), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n580), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n623), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n795), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n718), .A2(new_n720), .A3(new_n792), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(new_n801), .A3(KEYINPUT107), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n776), .A2(new_n794), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n803), .A2(KEYINPUT110), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT110), .B1(new_n803), .B2(new_n804), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n800), .A2(new_n801), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n772), .A2(new_n760), .B1(new_n770), .B2(new_n763), .ZN(new_n809));
  OR3_X1    g623(.A1(new_n808), .A2(new_n809), .A3(new_n804), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n757), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n776), .A2(KEYINPUT53), .A3(new_n801), .A4(new_n800), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n804), .B1(new_n808), .B2(new_n809), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n812), .A2(new_n757), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT111), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n814), .B(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT112), .B1(new_n811), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n723), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n727), .A2(new_n414), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n688), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n347), .A2(new_n669), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n476), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n818), .B(new_n820), .C1(new_n752), .C2(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n653), .A2(new_n723), .A3(new_n670), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n414), .A3(new_n577), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n825), .A2(new_n474), .A3(new_n596), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n826), .A2(KEYINPUT113), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n819), .A2(new_n670), .A3(new_n723), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n828), .A2(new_n693), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n826), .A2(KEYINPUT113), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n827), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n689), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n819), .A2(new_n187), .A3(new_n660), .A4(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT50), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n823), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n825), .A2(new_n597), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n831), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n836), .B1(new_n831), .B2(new_n839), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n823), .A3(new_n841), .A4(new_n834), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n410), .A2(new_n837), .A3(new_n838), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n803), .A2(new_n804), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT110), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n803), .A2(KEYINPUT110), .A3(new_n804), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n810), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT54), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n814), .B(KEYINPUT111), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT112), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n820), .A2(new_n679), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n817), .A2(new_n843), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n828), .A2(new_n712), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(KEYINPUT48), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n855), .B(new_n857), .Z(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n856), .B2(KEYINPUT48), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(G952), .A2(G953), .ZN(new_n861));
  INV_X1    g675(.A(new_n660), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n862), .B(new_n683), .C1(KEYINPUT49), .C2(new_n821), .ZN(new_n863));
  AOI211_X1 g677(.A(new_n653), .B(new_n863), .C1(KEYINPUT49), .C2(new_n821), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n187), .A3(new_n476), .ZN(new_n865));
  OAI22_X1  g679(.A1(new_n860), .A2(new_n861), .B1(new_n726), .B2(new_n865), .ZN(G75));
  AOI21_X1  g680(.A(new_n270), .B1(new_n812), .B2(new_n813), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT56), .B1(new_n867), .B2(G210), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n243), .B(new_n268), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT55), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n868), .B(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n264), .A2(G952), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(KEYINPUT116), .Z(G51));
  INV_X1    g689(.A(KEYINPUT117), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n814), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n814), .A2(new_n876), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n812), .A2(new_n813), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n879), .B1(new_n880), .B2(KEYINPUT54), .ZN(new_n881));
  AOI211_X1 g695(.A(KEYINPUT118), .B(new_n757), .C1(new_n812), .C2(new_n813), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n877), .B(new_n878), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n348), .B(KEYINPUT57), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n668), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT119), .ZN(new_n886));
  INV_X1    g700(.A(new_n867), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n887), .A2(new_n736), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n872), .B1(new_n886), .B2(new_n888), .ZN(G54));
  NAND3_X1  g703(.A1(new_n867), .A2(KEYINPUT58), .A3(G475), .ZN(new_n890));
  INV_X1    g704(.A(new_n472), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT120), .Z(new_n893));
  OAI21_X1  g707(.A(new_n873), .B1(new_n890), .B2(new_n891), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(G60));
  NAND2_X1  g709(.A1(G478), .A2(G902), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT59), .Z(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n588), .B(KEYINPUT121), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n883), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n873), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n897), .B1(new_n817), .B2(new_n852), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n903), .B1(new_n904), .B2(new_n900), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n849), .A2(new_n851), .A3(new_n850), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n851), .B1(new_n849), .B2(new_n850), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n898), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(KEYINPUT122), .A3(new_n899), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n902), .B1(new_n905), .B2(new_n909), .ZN(G63));
  NAND2_X1  g724(.A1(G217), .A2(G902), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT60), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n812), .B2(new_n813), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n873), .B1(new_n913), .B2(new_n571), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n620), .B2(new_n913), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(new_n914), .B2(KEYINPUT123), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n915), .B(new_n917), .ZN(G66));
  AOI21_X1  g732(.A(new_n264), .B1(new_n416), .B2(G224), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n786), .B2(new_n264), .ZN(new_n920));
  INV_X1    g734(.A(G898), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n243), .B1(new_n921), .B2(G953), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT124), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n920), .B(new_n923), .ZN(G69));
  OAI21_X1  g738(.A(G953), .B1(new_n326), .B2(new_n639), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n506), .B(new_n459), .Z(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n746), .A2(new_n755), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n774), .A2(new_n765), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n928), .A2(new_n718), .A3(new_n720), .A4(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n712), .ZN(new_n932));
  NOR4_X1   g746(.A1(new_n742), .A2(new_n722), .A3(new_n646), .A4(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n264), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n639), .A2(G953), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT126), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n927), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n925), .B1(new_n937), .B2(KEYINPUT125), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n930), .A2(new_n661), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n939), .A2(KEYINPUT62), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(KEYINPUT62), .ZN(new_n941));
  INV_X1    g755(.A(new_n657), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n780), .A2(new_n942), .A3(new_n818), .A4(new_n796), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n928), .A2(new_n940), .A3(new_n941), .A4(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n926), .B1(new_n944), .B2(new_n264), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n937), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n938), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n934), .A2(new_n936), .ZN(new_n948));
  AOI221_X4 g762(.A(new_n945), .B1(KEYINPUT125), .B2(new_n925), .C1(new_n948), .C2(new_n926), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n947), .A2(new_n949), .ZN(G72));
  NAND2_X1  g764(.A1(G472), .A2(G902), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT63), .Z(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(new_n944), .B2(new_n786), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n872), .B1(new_n953), .B2(new_n651), .ZN(new_n954));
  INV_X1    g768(.A(new_n952), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n931), .A2(new_n933), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n955), .B1(new_n956), .B2(new_n800), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n954), .B1(new_n957), .B2(new_n525), .ZN(new_n958));
  INV_X1    g772(.A(new_n651), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n848), .A2(new_n525), .A3(new_n959), .A4(new_n952), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT127), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n958), .A2(new_n961), .ZN(G57));
endmodule


