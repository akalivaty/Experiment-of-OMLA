

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U554 ( .A1(n585), .A2(n584), .ZN(G164) );
  NOR2_X4 U555 ( .A1(G2104), .A2(n525), .ZN(n881) );
  NOR2_X1 U556 ( .A1(n795), .A2(n794), .ZN(n797) );
  BUF_X1 U557 ( .A(n578), .Z(n558) );
  NAND2_X2 U558 ( .A1(n690), .A2(G8), .ZN(n771) );
  NOR2_X1 U559 ( .A1(n956), .A2(n706), .ZN(n705) );
  INV_X1 U560 ( .A(KEYINPUT95), .ZN(n692) );
  NAND2_X1 U561 ( .A1(n722), .A2(n721), .ZN(n724) );
  OR2_X1 U562 ( .A1(n523), .A2(G2105), .ZN(n524) );
  XNOR2_X2 U563 ( .A(n687), .B(KEYINPUT64), .ZN(n690) );
  NOR2_X1 U564 ( .A1(n771), .A2(n758), .ZN(n521) );
  OR2_X1 U565 ( .A1(n820), .A2(n1017), .ZN(n522) );
  XNOR2_X1 U566 ( .A(n701), .B(KEYINPUT93), .ZN(n704) );
  INV_X1 U567 ( .A(KEYINPUT29), .ZN(n723) );
  XNOR2_X1 U568 ( .A(n724), .B(n723), .ZN(n727) );
  OR2_X1 U569 ( .A1(n690), .A2(G2084), .ZN(n691) );
  NOR2_X1 U570 ( .A1(G1384), .A2(G164), .ZN(n685) );
  INV_X1 U571 ( .A(G2105), .ZN(n525) );
  INV_X1 U572 ( .A(KEYINPUT99), .ZN(n796) );
  AND2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n883) );
  NOR2_X1 U574 ( .A1(n533), .A2(n532), .ZN(G160) );
  NAND2_X1 U575 ( .A1(G2104), .A2(G101), .ZN(n523) );
  XOR2_X1 U576 ( .A(n524), .B(KEYINPUT23), .Z(n527) );
  NAND2_X1 U577 ( .A1(n881), .A2(G125), .ZN(n526) );
  NAND2_X1 U578 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U579 ( .A(n528), .B(KEYINPUT66), .ZN(n533) );
  NOR2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  XOR2_X1 U581 ( .A(KEYINPUT17), .B(n529), .Z(n578) );
  NAND2_X1 U582 ( .A1(n578), .A2(G137), .ZN(n531) );
  NAND2_X1 U583 ( .A1(n883), .A2(G113), .ZN(n530) );
  NAND2_X1 U584 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U585 ( .A1(G651), .A2(G543), .ZN(n648) );
  NAND2_X1 U586 ( .A1(G85), .A2(n648), .ZN(n535) );
  XOR2_X1 U587 ( .A(KEYINPUT0), .B(G543), .Z(n641) );
  INV_X1 U588 ( .A(G651), .ZN(n536) );
  NOR2_X1 U589 ( .A1(n641), .A2(n536), .ZN(n644) );
  NAND2_X1 U590 ( .A1(G72), .A2(n644), .ZN(n534) );
  NAND2_X1 U591 ( .A1(n535), .A2(n534), .ZN(n541) );
  NOR2_X1 U592 ( .A1(G543), .A2(n536), .ZN(n537) );
  XOR2_X1 U593 ( .A(KEYINPUT1), .B(n537), .Z(n647) );
  NAND2_X1 U594 ( .A1(G60), .A2(n647), .ZN(n539) );
  NOR2_X1 U595 ( .A1(G651), .A2(n641), .ZN(n654) );
  NAND2_X1 U596 ( .A1(G47), .A2(n654), .ZN(n538) );
  NAND2_X1 U597 ( .A1(n539), .A2(n538), .ZN(n540) );
  OR2_X1 U598 ( .A1(n541), .A2(n540), .ZN(G290) );
  NAND2_X1 U599 ( .A1(n647), .A2(G62), .ZN(n548) );
  NAND2_X1 U600 ( .A1(G75), .A2(n644), .ZN(n543) );
  NAND2_X1 U601 ( .A1(G50), .A2(n654), .ZN(n542) );
  NAND2_X1 U602 ( .A1(n543), .A2(n542), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n648), .A2(G88), .ZN(n544) );
  XOR2_X1 U604 ( .A(KEYINPUT80), .B(n544), .Z(n545) );
  NOR2_X1 U605 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U607 ( .A(KEYINPUT81), .B(n549), .Z(G303) );
  INV_X1 U608 ( .A(G303), .ZN(G166) );
  NAND2_X1 U609 ( .A1(G64), .A2(n647), .ZN(n550) );
  XNOR2_X1 U610 ( .A(n550), .B(KEYINPUT67), .ZN(n557) );
  NAND2_X1 U611 ( .A1(G90), .A2(n648), .ZN(n552) );
  NAND2_X1 U612 ( .A1(G77), .A2(n644), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U614 ( .A(n553), .B(KEYINPUT9), .ZN(n555) );
  NAND2_X1 U615 ( .A1(G52), .A2(n654), .ZN(n554) );
  NAND2_X1 U616 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U617 ( .A1(n557), .A2(n556), .ZN(G171) );
  AND2_X1 U618 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U619 ( .A1(G111), .A2(n883), .ZN(n560) );
  NAND2_X1 U620 ( .A1(G135), .A2(n558), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n560), .A2(n559), .ZN(n563) );
  NAND2_X1 U622 ( .A1(n881), .A2(G123), .ZN(n561) );
  XOR2_X1 U623 ( .A(KEYINPUT18), .B(n561), .Z(n562) );
  NOR2_X1 U624 ( .A1(n563), .A2(n562), .ZN(n565) );
  AND2_X1 U625 ( .A1(n525), .A2(G2104), .ZN(n889) );
  NAND2_X1 U626 ( .A1(n889), .A2(G99), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n565), .A2(n564), .ZN(n1008) );
  XNOR2_X1 U628 ( .A(G2096), .B(n1008), .ZN(n566) );
  OR2_X1 U629 ( .A1(G2100), .A2(n566), .ZN(G156) );
  INV_X1 U630 ( .A(G860), .ZN(n621) );
  NAND2_X1 U631 ( .A1(G81), .A2(n648), .ZN(n567) );
  XOR2_X1 U632 ( .A(KEYINPUT71), .B(n567), .Z(n568) );
  XNOR2_X1 U633 ( .A(n568), .B(KEYINPUT12), .ZN(n570) );
  NAND2_X1 U634 ( .A1(G68), .A2(n644), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(KEYINPUT13), .ZN(n573) );
  NAND2_X1 U637 ( .A1(G43), .A2(n654), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U639 ( .A1(n647), .A2(G56), .ZN(n574) );
  XOR2_X1 U640 ( .A(KEYINPUT14), .B(n574), .Z(n575) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U642 ( .A(KEYINPUT72), .B(n577), .Z(n953) );
  OR2_X1 U643 ( .A1(n621), .A2(n953), .ZN(G153) );
  INV_X1 U644 ( .A(G132), .ZN(G219) );
  INV_X1 U645 ( .A(G82), .ZN(G220) );
  INV_X1 U646 ( .A(G57), .ZN(G237) );
  NAND2_X1 U647 ( .A1(n578), .A2(G138), .ZN(n581) );
  NAND2_X1 U648 ( .A1(G126), .A2(n881), .ZN(n579) );
  XOR2_X1 U649 ( .A(KEYINPUT85), .B(n579), .Z(n580) );
  NAND2_X1 U650 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U651 ( .A1(G102), .A2(n889), .ZN(n583) );
  NAND2_X1 U652 ( .A1(G114), .A2(n883), .ZN(n582) );
  NAND2_X1 U653 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n648), .A2(G89), .ZN(n586) );
  XNOR2_X1 U655 ( .A(n586), .B(KEYINPUT4), .ZN(n588) );
  NAND2_X1 U656 ( .A1(G76), .A2(n644), .ZN(n587) );
  NAND2_X1 U657 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U658 ( .A(KEYINPUT5), .B(n589), .ZN(n595) );
  NAND2_X1 U659 ( .A1(G63), .A2(n647), .ZN(n591) );
  NAND2_X1 U660 ( .A1(G51), .A2(n654), .ZN(n590) );
  NAND2_X1 U661 ( .A1(n591), .A2(n590), .ZN(n593) );
  XOR2_X1 U662 ( .A(KEYINPUT6), .B(KEYINPUT74), .Z(n592) );
  XNOR2_X1 U663 ( .A(n593), .B(n592), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U665 ( .A(KEYINPUT7), .B(n596), .ZN(G168) );
  XOR2_X1 U666 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U667 ( .A1(G7), .A2(G661), .ZN(n597) );
  XNOR2_X1 U668 ( .A(n597), .B(KEYINPUT10), .ZN(n598) );
  XNOR2_X1 U669 ( .A(KEYINPUT70), .B(n598), .ZN(G223) );
  INV_X1 U670 ( .A(G223), .ZN(n826) );
  NAND2_X1 U671 ( .A1(n826), .A2(G567), .ZN(n599) );
  XOR2_X1 U672 ( .A(KEYINPUT11), .B(n599), .Z(G234) );
  INV_X1 U673 ( .A(G171), .ZN(G301) );
  NAND2_X1 U674 ( .A1(G868), .A2(G301), .ZN(n609) );
  NAND2_X1 U675 ( .A1(n647), .A2(G66), .ZN(n606) );
  NAND2_X1 U676 ( .A1(G79), .A2(n644), .ZN(n601) );
  NAND2_X1 U677 ( .A1(G54), .A2(n654), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U679 ( .A1(G92), .A2(n648), .ZN(n602) );
  XNOR2_X1 U680 ( .A(KEYINPUT73), .B(n602), .ZN(n603) );
  NOR2_X1 U681 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U682 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U683 ( .A(KEYINPUT15), .B(n607), .Z(n948) );
  INV_X1 U684 ( .A(G868), .ZN(n666) );
  NAND2_X1 U685 ( .A1(n948), .A2(n666), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n609), .A2(n608), .ZN(G284) );
  NAND2_X1 U687 ( .A1(G91), .A2(n648), .ZN(n611) );
  NAND2_X1 U688 ( .A1(G78), .A2(n644), .ZN(n610) );
  NAND2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U690 ( .A(KEYINPUT68), .B(n612), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G53), .A2(n654), .ZN(n613) );
  XNOR2_X1 U692 ( .A(KEYINPUT69), .B(n613), .ZN(n614) );
  NOR2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U694 ( .A1(n647), .A2(G65), .ZN(n616) );
  NAND2_X1 U695 ( .A1(n617), .A2(n616), .ZN(G299) );
  NOR2_X1 U696 ( .A1(G286), .A2(n666), .ZN(n619) );
  NOR2_X1 U697 ( .A1(G868), .A2(G299), .ZN(n618) );
  NOR2_X1 U698 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U699 ( .A(KEYINPUT75), .B(n620), .Z(G297) );
  NAND2_X1 U700 ( .A1(n621), .A2(G559), .ZN(n622) );
  INV_X1 U701 ( .A(n948), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n622), .A2(n627), .ZN(n623) );
  XNOR2_X1 U703 ( .A(n623), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U704 ( .A1(n953), .A2(G868), .ZN(n626) );
  NAND2_X1 U705 ( .A1(G868), .A2(n627), .ZN(n624) );
  NOR2_X1 U706 ( .A1(G559), .A2(n624), .ZN(n625) );
  NOR2_X1 U707 ( .A1(n626), .A2(n625), .ZN(G282) );
  NAND2_X1 U708 ( .A1(G559), .A2(n627), .ZN(n628) );
  XNOR2_X1 U709 ( .A(n628), .B(n953), .ZN(n663) );
  XNOR2_X1 U710 ( .A(KEYINPUT76), .B(n663), .ZN(n629) );
  NOR2_X1 U711 ( .A1(G860), .A2(n629), .ZN(n637) );
  NAND2_X1 U712 ( .A1(G80), .A2(n644), .ZN(n631) );
  NAND2_X1 U713 ( .A1(G55), .A2(n654), .ZN(n630) );
  NAND2_X1 U714 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U715 ( .A1(G93), .A2(n648), .ZN(n632) );
  XNOR2_X1 U716 ( .A(KEYINPUT77), .B(n632), .ZN(n633) );
  NOR2_X1 U717 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U718 ( .A1(n647), .A2(G67), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n636), .A2(n635), .ZN(n665) );
  XOR2_X1 U720 ( .A(n637), .B(n665), .Z(G145) );
  NAND2_X1 U721 ( .A1(G49), .A2(n654), .ZN(n639) );
  NAND2_X1 U722 ( .A1(G74), .A2(G651), .ZN(n638) );
  NAND2_X1 U723 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U724 ( .A1(n647), .A2(n640), .ZN(n643) );
  NAND2_X1 U725 ( .A1(n641), .A2(G87), .ZN(n642) );
  NAND2_X1 U726 ( .A1(n643), .A2(n642), .ZN(G288) );
  XOR2_X1 U727 ( .A(KEYINPUT78), .B(KEYINPUT2), .Z(n646) );
  NAND2_X1 U728 ( .A1(G73), .A2(n644), .ZN(n645) );
  XNOR2_X1 U729 ( .A(n646), .B(n645), .ZN(n652) );
  NAND2_X1 U730 ( .A1(n647), .A2(G61), .ZN(n650) );
  NAND2_X1 U731 ( .A1(n648), .A2(G86), .ZN(n649) );
  NAND2_X1 U732 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U733 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U734 ( .A(KEYINPUT79), .B(n653), .Z(n656) );
  NAND2_X1 U735 ( .A1(n654), .A2(G48), .ZN(n655) );
  NAND2_X1 U736 ( .A1(n656), .A2(n655), .ZN(G305) );
  XOR2_X1 U737 ( .A(KEYINPUT19), .B(KEYINPUT82), .Z(n657) );
  XNOR2_X1 U738 ( .A(G290), .B(n657), .ZN(n660) );
  INV_X1 U739 ( .A(G299), .ZN(n956) );
  XNOR2_X1 U740 ( .A(n956), .B(G288), .ZN(n658) );
  XNOR2_X1 U741 ( .A(n658), .B(n665), .ZN(n659) );
  XNOR2_X1 U742 ( .A(n660), .B(n659), .ZN(n662) );
  XNOR2_X1 U743 ( .A(G305), .B(G166), .ZN(n661) );
  XNOR2_X1 U744 ( .A(n662), .B(n661), .ZN(n901) );
  XNOR2_X1 U745 ( .A(n663), .B(n901), .ZN(n664) );
  NAND2_X1 U746 ( .A1(n664), .A2(G868), .ZN(n668) );
  NAND2_X1 U747 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U748 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XNOR2_X1 U750 ( .A(n669), .B(KEYINPUT20), .ZN(n670) );
  XNOR2_X1 U751 ( .A(n670), .B(KEYINPUT83), .ZN(n671) );
  NAND2_X1 U752 ( .A1(n671), .A2(G2090), .ZN(n672) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U754 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U756 ( .A1(G69), .A2(G120), .ZN(n674) );
  NOR2_X1 U757 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U758 ( .A1(G108), .A2(n675), .ZN(n831) );
  NAND2_X1 U759 ( .A1(n831), .A2(G567), .ZN(n681) );
  NOR2_X1 U760 ( .A1(G220), .A2(G219), .ZN(n676) );
  XOR2_X1 U761 ( .A(KEYINPUT22), .B(n676), .Z(n677) );
  NOR2_X1 U762 ( .A1(G218), .A2(n677), .ZN(n678) );
  NAND2_X1 U763 ( .A1(G96), .A2(n678), .ZN(n830) );
  NAND2_X1 U764 ( .A1(G2106), .A2(n830), .ZN(n679) );
  XNOR2_X1 U765 ( .A(KEYINPUT84), .B(n679), .ZN(n680) );
  NAND2_X1 U766 ( .A1(n681), .A2(n680), .ZN(n832) );
  NAND2_X1 U767 ( .A1(G483), .A2(G661), .ZN(n682) );
  NOR2_X1 U768 ( .A1(n832), .A2(n682), .ZN(n829) );
  NAND2_X1 U769 ( .A1(n829), .A2(G36), .ZN(G176) );
  NAND2_X1 U770 ( .A1(G40), .A2(G160), .ZN(n683) );
  XOR2_X1 U771 ( .A(KEYINPUT86), .B(n683), .Z(n775) );
  XNOR2_X1 U772 ( .A(n685), .B(KEYINPUT65), .ZN(n774) );
  INV_X1 U773 ( .A(n774), .ZN(n686) );
  NAND2_X1 U774 ( .A1(n775), .A2(n686), .ZN(n687) );
  INV_X1 U775 ( .A(n690), .ZN(n711) );
  XNOR2_X1 U776 ( .A(KEYINPUT25), .B(G2078), .ZN(n926) );
  NAND2_X1 U777 ( .A1(n711), .A2(n926), .ZN(n689) );
  XOR2_X1 U778 ( .A(G1961), .B(KEYINPUT92), .Z(n991) );
  NAND2_X1 U779 ( .A1(n690), .A2(n991), .ZN(n688) );
  NAND2_X1 U780 ( .A1(n689), .A2(n688), .ZN(n725) );
  NOR2_X1 U781 ( .A1(G171), .A2(n725), .ZN(n698) );
  NOR2_X1 U782 ( .A1(G1966), .A2(n771), .ZN(n742) );
  XNOR2_X1 U783 ( .A(KEYINPUT91), .B(n691), .ZN(n739) );
  NOR2_X1 U784 ( .A1(n742), .A2(n739), .ZN(n693) );
  XNOR2_X1 U785 ( .A(n693), .B(n692), .ZN(n694) );
  NAND2_X1 U786 ( .A1(n694), .A2(G8), .ZN(n695) );
  XNOR2_X1 U787 ( .A(KEYINPUT30), .B(n695), .ZN(n696) );
  NOR2_X1 U788 ( .A1(G168), .A2(n696), .ZN(n697) );
  NOR2_X1 U789 ( .A1(n698), .A2(n697), .ZN(n700) );
  INV_X1 U790 ( .A(KEYINPUT31), .ZN(n699) );
  XNOR2_X1 U791 ( .A(n700), .B(n699), .ZN(n741) );
  NAND2_X1 U792 ( .A1(n690), .A2(G1956), .ZN(n701) );
  NAND2_X1 U793 ( .A1(G2072), .A2(n711), .ZN(n702) );
  XNOR2_X1 U794 ( .A(KEYINPUT27), .B(n702), .ZN(n703) );
  NOR2_X1 U795 ( .A1(n704), .A2(n703), .ZN(n706) );
  XOR2_X1 U796 ( .A(n705), .B(KEYINPUT28), .Z(n722) );
  NAND2_X1 U797 ( .A1(n956), .A2(n706), .ZN(n720) );
  XOR2_X1 U798 ( .A(KEYINPUT94), .B(G1996), .Z(n925) );
  NOR2_X1 U799 ( .A1(n690), .A2(n925), .ZN(n707) );
  XOR2_X1 U800 ( .A(n707), .B(KEYINPUT26), .Z(n709) );
  NAND2_X1 U801 ( .A1(n690), .A2(G1341), .ZN(n708) );
  NAND2_X1 U802 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U803 ( .A1(n953), .A2(n710), .ZN(n715) );
  NAND2_X1 U804 ( .A1(G2067), .A2(n711), .ZN(n713) );
  NAND2_X1 U805 ( .A1(n690), .A2(G1348), .ZN(n712) );
  NAND2_X1 U806 ( .A1(n713), .A2(n712), .ZN(n716) );
  NOR2_X1 U807 ( .A1(n948), .A2(n716), .ZN(n714) );
  OR2_X1 U808 ( .A1(n715), .A2(n714), .ZN(n718) );
  NAND2_X1 U809 ( .A1(n948), .A2(n716), .ZN(n717) );
  NAND2_X1 U810 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U811 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U812 ( .A1(G171), .A2(n725), .ZN(n726) );
  NAND2_X1 U813 ( .A1(n727), .A2(n726), .ZN(n740) );
  INV_X1 U814 ( .A(G8), .ZN(n732) );
  NOR2_X1 U815 ( .A1(G1971), .A2(n771), .ZN(n729) );
  NOR2_X1 U816 ( .A1(n690), .A2(G2090), .ZN(n728) );
  NOR2_X1 U817 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U818 ( .A1(n730), .A2(G303), .ZN(n731) );
  OR2_X1 U819 ( .A1(n732), .A2(n731), .ZN(n734) );
  AND2_X1 U820 ( .A1(n740), .A2(n734), .ZN(n733) );
  NAND2_X1 U821 ( .A1(n741), .A2(n733), .ZN(n737) );
  INV_X1 U822 ( .A(n734), .ZN(n735) );
  OR2_X1 U823 ( .A1(n735), .A2(G286), .ZN(n736) );
  NAND2_X1 U824 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U825 ( .A(n738), .B(KEYINPUT32), .ZN(n747) );
  NAND2_X1 U826 ( .A1(G8), .A2(n739), .ZN(n745) );
  AND2_X1 U827 ( .A1(n741), .A2(n740), .ZN(n743) );
  NOR2_X1 U828 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U829 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U830 ( .A1(n747), .A2(n746), .ZN(n757) );
  NAND2_X1 U831 ( .A1(G8), .A2(G166), .ZN(n748) );
  NOR2_X1 U832 ( .A1(G2090), .A2(n748), .ZN(n749) );
  XNOR2_X1 U833 ( .A(n749), .B(KEYINPUT97), .ZN(n750) );
  NAND2_X1 U834 ( .A1(n757), .A2(n750), .ZN(n751) );
  NAND2_X1 U835 ( .A1(n751), .A2(n771), .ZN(n766) );
  NOR2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n945) );
  NOR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n752) );
  XNOR2_X1 U838 ( .A(KEYINPUT96), .B(n752), .ZN(n753) );
  NOR2_X1 U839 ( .A1(n945), .A2(n753), .ZN(n755) );
  INV_X1 U840 ( .A(KEYINPUT33), .ZN(n754) );
  AND2_X1 U841 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U842 ( .A1(n757), .A2(n756), .ZN(n764) );
  NAND2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n946) );
  INV_X1 U844 ( .A(n946), .ZN(n758) );
  NOR2_X1 U845 ( .A1(KEYINPUT33), .A2(n521), .ZN(n761) );
  NAND2_X1 U846 ( .A1(n945), .A2(KEYINPUT33), .ZN(n759) );
  NOR2_X1 U847 ( .A1(n759), .A2(n771), .ZN(n760) );
  NOR2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U849 ( .A(G1981), .B(G305), .Z(n959) );
  AND2_X1 U850 ( .A1(n762), .A2(n959), .ZN(n763) );
  NAND2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U852 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U853 ( .A(n767), .B(KEYINPUT98), .ZN(n773) );
  NOR2_X1 U854 ( .A1(G1981), .A2(G305), .ZN(n768) );
  XOR2_X1 U855 ( .A(n768), .B(KEYINPUT24), .Z(n769) );
  XNOR2_X1 U856 ( .A(KEYINPUT90), .B(n769), .ZN(n770) );
  NOR2_X1 U857 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U858 ( .A1(n773), .A2(n772), .ZN(n795) );
  NAND2_X1 U859 ( .A1(n775), .A2(n774), .ZN(n820) );
  NAND2_X1 U860 ( .A1(G107), .A2(n883), .ZN(n777) );
  NAND2_X1 U861 ( .A1(G131), .A2(n558), .ZN(n776) );
  NAND2_X1 U862 ( .A1(n777), .A2(n776), .ZN(n781) );
  NAND2_X1 U863 ( .A1(G95), .A2(n889), .ZN(n779) );
  NAND2_X1 U864 ( .A1(G119), .A2(n881), .ZN(n778) );
  NAND2_X1 U865 ( .A1(n779), .A2(n778), .ZN(n780) );
  OR2_X1 U866 ( .A1(n781), .A2(n780), .ZN(n864) );
  NAND2_X1 U867 ( .A1(G1991), .A2(n864), .ZN(n792) );
  NAND2_X1 U868 ( .A1(G117), .A2(n883), .ZN(n783) );
  NAND2_X1 U869 ( .A1(G141), .A2(n558), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n788) );
  XOR2_X1 U871 ( .A(KEYINPUT38), .B(KEYINPUT89), .Z(n785) );
  NAND2_X1 U872 ( .A1(G105), .A2(n889), .ZN(n784) );
  XNOR2_X1 U873 ( .A(n785), .B(n784), .ZN(n786) );
  XOR2_X1 U874 ( .A(KEYINPUT88), .B(n786), .Z(n787) );
  NOR2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n790) );
  NAND2_X1 U876 ( .A1(n881), .A2(G129), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n877) );
  NAND2_X1 U878 ( .A1(G1996), .A2(n877), .ZN(n791) );
  NAND2_X1 U879 ( .A1(n792), .A2(n791), .ZN(n1006) );
  XNOR2_X1 U880 ( .A(G1986), .B(G290), .ZN(n944) );
  NOR2_X1 U881 ( .A1(n1006), .A2(n944), .ZN(n793) );
  NOR2_X1 U882 ( .A1(n820), .A2(n793), .ZN(n794) );
  XNOR2_X1 U883 ( .A(n797), .B(n796), .ZN(n808) );
  XOR2_X1 U884 ( .A(G2067), .B(KEYINPUT37), .Z(n809) );
  NAND2_X1 U885 ( .A1(G104), .A2(n889), .ZN(n799) );
  NAND2_X1 U886 ( .A1(G140), .A2(n558), .ZN(n798) );
  NAND2_X1 U887 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U888 ( .A(KEYINPUT34), .B(n800), .ZN(n806) );
  NAND2_X1 U889 ( .A1(G128), .A2(n881), .ZN(n802) );
  NAND2_X1 U890 ( .A1(G116), .A2(n883), .ZN(n801) );
  NAND2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U892 ( .A(KEYINPUT87), .B(n803), .ZN(n804) );
  XNOR2_X1 U893 ( .A(KEYINPUT35), .B(n804), .ZN(n805) );
  NOR2_X1 U894 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U895 ( .A(KEYINPUT36), .B(n807), .Z(n898) );
  NAND2_X1 U896 ( .A1(n809), .A2(n898), .ZN(n1017) );
  NAND2_X1 U897 ( .A1(n808), .A2(n522), .ZN(n824) );
  INV_X1 U898 ( .A(n1017), .ZN(n816) );
  NAND2_X1 U899 ( .A1(n816), .A2(KEYINPUT99), .ZN(n819) );
  NOR2_X1 U900 ( .A1(n809), .A2(n898), .ZN(n1023) );
  NOR2_X1 U901 ( .A1(G1996), .A2(n877), .ZN(n1011) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n810) );
  NOR2_X1 U903 ( .A1(G1991), .A2(n864), .ZN(n1007) );
  NOR2_X1 U904 ( .A1(n810), .A2(n1007), .ZN(n811) );
  XNOR2_X1 U905 ( .A(n811), .B(KEYINPUT100), .ZN(n812) );
  NOR2_X1 U906 ( .A1(n1006), .A2(n812), .ZN(n813) );
  NOR2_X1 U907 ( .A1(n1011), .A2(n813), .ZN(n814) );
  XOR2_X1 U908 ( .A(KEYINPUT39), .B(n814), .Z(n815) );
  NOR2_X1 U909 ( .A1(n816), .A2(n815), .ZN(n817) );
  NOR2_X1 U910 ( .A1(n1023), .A2(n817), .ZN(n818) );
  NAND2_X1 U911 ( .A1(n819), .A2(n818), .ZN(n822) );
  INV_X1 U912 ( .A(n820), .ZN(n821) );
  NAND2_X1 U913 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U914 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U915 ( .A(n825), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n826), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U918 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U920 ( .A1(n829), .A2(n828), .ZN(G188) );
  INV_X1 U922 ( .A(G120), .ZN(G236) );
  INV_X1 U923 ( .A(G96), .ZN(G221) );
  INV_X1 U924 ( .A(G69), .ZN(G235) );
  NOR2_X1 U925 ( .A1(n831), .A2(n830), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  INV_X1 U927 ( .A(n832), .ZN(G319) );
  XNOR2_X1 U928 ( .A(G1971), .B(KEYINPUT41), .ZN(n842) );
  XOR2_X1 U929 ( .A(G1986), .B(G1976), .Z(n834) );
  XNOR2_X1 U930 ( .A(G1961), .B(G1956), .ZN(n833) );
  XNOR2_X1 U931 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U932 ( .A(G1991), .B(G1996), .Z(n836) );
  XNOR2_X1 U933 ( .A(G1981), .B(G1966), .ZN(n835) );
  XNOR2_X1 U934 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U935 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U936 ( .A(KEYINPUT104), .B(G2474), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(G229) );
  XOR2_X1 U939 ( .A(KEYINPUT43), .B(G2678), .Z(n844) );
  XNOR2_X1 U940 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U942 ( .A(KEYINPUT42), .B(G2090), .Z(n846) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2072), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U945 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U946 ( .A(G2096), .B(G2100), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(n852) );
  XOR2_X1 U948 ( .A(G2078), .B(G2084), .Z(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(G227) );
  NAND2_X1 U950 ( .A1(n889), .A2(G100), .ZN(n853) );
  XOR2_X1 U951 ( .A(KEYINPUT107), .B(n853), .Z(n855) );
  NAND2_X1 U952 ( .A1(n883), .A2(G112), .ZN(n854) );
  NAND2_X1 U953 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U954 ( .A(KEYINPUT108), .B(n856), .ZN(n863) );
  NAND2_X1 U955 ( .A1(G136), .A2(n558), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n857), .B(KEYINPUT106), .ZN(n861) );
  XOR2_X1 U957 ( .A(KEYINPUT105), .B(KEYINPUT44), .Z(n859) );
  NAND2_X1 U958 ( .A1(G124), .A2(n881), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(n860) );
  NAND2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U961 ( .A1(n863), .A2(n862), .ZN(G162) );
  XNOR2_X1 U962 ( .A(G160), .B(G162), .ZN(n897) );
  XNOR2_X1 U963 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n866) );
  XNOR2_X1 U964 ( .A(n864), .B(KEYINPUT114), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n867) );
  XNOR2_X1 U966 ( .A(KEYINPUT110), .B(n867), .ZN(n879) );
  NAND2_X1 U967 ( .A1(G130), .A2(n881), .ZN(n869) );
  NAND2_X1 U968 ( .A1(G118), .A2(n883), .ZN(n868) );
  NAND2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n875) );
  NAND2_X1 U970 ( .A1(G106), .A2(n889), .ZN(n871) );
  NAND2_X1 U971 ( .A1(G142), .A2(n558), .ZN(n870) );
  NAND2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U973 ( .A(KEYINPUT109), .B(n872), .ZN(n873) );
  XNOR2_X1 U974 ( .A(KEYINPUT45), .B(n873), .ZN(n874) );
  NOR2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U976 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U977 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U978 ( .A(n1008), .B(n880), .ZN(n895) );
  NAND2_X1 U979 ( .A1(n881), .A2(G127), .ZN(n882) );
  XNOR2_X1 U980 ( .A(n882), .B(KEYINPUT112), .ZN(n885) );
  NAND2_X1 U981 ( .A1(G115), .A2(n883), .ZN(n884) );
  NAND2_X1 U982 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U983 ( .A(n886), .B(KEYINPUT47), .ZN(n888) );
  NAND2_X1 U984 ( .A1(G139), .A2(n558), .ZN(n887) );
  NAND2_X1 U985 ( .A1(n888), .A2(n887), .ZN(n892) );
  NAND2_X1 U986 ( .A1(G103), .A2(n889), .ZN(n890) );
  XNOR2_X1 U987 ( .A(KEYINPUT111), .B(n890), .ZN(n891) );
  NOR2_X1 U988 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U989 ( .A(KEYINPUT113), .B(n893), .Z(n1001) );
  XNOR2_X1 U990 ( .A(G164), .B(n1001), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n897), .B(n896), .ZN(n899) );
  XNOR2_X1 U993 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U994 ( .A1(G37), .A2(n900), .ZN(G395) );
  XNOR2_X1 U995 ( .A(n948), .B(n901), .ZN(n903) );
  XNOR2_X1 U996 ( .A(G171), .B(n953), .ZN(n902) );
  XNOR2_X1 U997 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U998 ( .A(n904), .B(G286), .ZN(n905) );
  NOR2_X1 U999 ( .A1(G37), .A2(n905), .ZN(G397) );
  XOR2_X1 U1000 ( .A(G2430), .B(G2451), .Z(n907) );
  XNOR2_X1 U1001 ( .A(G2446), .B(G2427), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n914) );
  XOR2_X1 U1003 ( .A(G2438), .B(KEYINPUT101), .Z(n909) );
  XNOR2_X1 U1004 ( .A(G2443), .B(G2454), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1006 ( .A(n910), .B(G2435), .Z(n912) );
  XNOR2_X1 U1007 ( .A(G1341), .B(G1348), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(n914), .B(n913), .ZN(n915) );
  NAND2_X1 U1010 ( .A1(n915), .A2(G14), .ZN(n921) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n921), .ZN(n918) );
  NOR2_X1 U1012 ( .A1(G229), .A2(G227), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1016 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(G108), .ZN(G238) );
  INV_X1 U1019 ( .A(n921), .ZN(G401) );
  XOR2_X1 U1020 ( .A(G29), .B(KEYINPUT120), .Z(n942) );
  XOR2_X1 U1021 ( .A(G1991), .B(G25), .Z(n922) );
  NAND2_X1 U1022 ( .A1(n922), .A2(G28), .ZN(n932) );
  XNOR2_X1 U1023 ( .A(G2067), .B(G26), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(G33), .B(G2072), .ZN(n923) );
  NOR2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n930) );
  XOR2_X1 U1026 ( .A(n925), .B(G32), .Z(n928) );
  XOR2_X1 U1027 ( .A(n926), .B(G27), .Z(n927) );
  NOR2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1031 ( .A(KEYINPUT53), .B(n933), .Z(n937) );
  XNOR2_X1 U1032 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(n934), .B(G34), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(G2084), .B(n935), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(G35), .B(G2090), .ZN(n938) );
  NOR2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1038 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n1025) );
  XOR2_X1 U1039 ( .A(n940), .B(n1025), .Z(n941) );
  NAND2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1041 ( .A1(G11), .A2(n943), .ZN(n1000) );
  XNOR2_X1 U1042 ( .A(G16), .B(KEYINPUT56), .ZN(n968) );
  XNOR2_X1 U1043 ( .A(G166), .B(G1971), .ZN(n952) );
  NOR2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n947) );
  NAND2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(G1348), .B(n948), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(G1341), .B(n953), .ZN(n954) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n966) );
  XNOR2_X1 U1051 ( .A(n956), .B(G1956), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(G171), .B(G1961), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n964) );
  XNOR2_X1 U1054 ( .A(G1966), .B(G168), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(n961), .B(KEYINPUT121), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(n962), .B(KEYINPUT57), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n998) );
  INV_X1 U1061 ( .A(G16), .ZN(n996) );
  XOR2_X1 U1062 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n978) );
  XNOR2_X1 U1063 ( .A(G1981), .B(G6), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(G1341), .B(G19), .ZN(n969) );
  NOR2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n976) );
  XOR2_X1 U1066 ( .A(KEYINPUT122), .B(G4), .Z(n972) );
  XNOR2_X1 U1067 ( .A(G1348), .B(KEYINPUT59), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(n972), .B(n971), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(G1956), .B(G20), .ZN(n973) );
  NOR2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(n978), .B(n977), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(G21), .B(G1966), .ZN(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(KEYINPUT124), .B(n981), .ZN(n990) );
  XOR2_X1 U1076 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n988) );
  XNOR2_X1 U1077 ( .A(G1971), .B(G22), .ZN(n983) );
  XNOR2_X1 U1078 ( .A(G1986), .B(G24), .ZN(n982) );
  NOR2_X1 U1079 ( .A1(n983), .A2(n982), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(G1976), .B(KEYINPUT125), .ZN(n984) );
  XNOR2_X1 U1081 ( .A(n984), .B(G23), .ZN(n985) );
  NAND2_X1 U1082 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1083 ( .A(n988), .B(n987), .ZN(n989) );
  NAND2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n993) );
  XOR2_X1 U1085 ( .A(n991), .B(G5), .Z(n992) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1087 ( .A(KEYINPUT61), .B(n994), .ZN(n995) );
  NAND2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1030) );
  XOR2_X1 U1091 ( .A(G2072), .B(n1001), .Z(n1003) );
  XOR2_X1 U1092 ( .A(G164), .B(G2078), .Z(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(KEYINPUT50), .B(n1004), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(n1005), .B(KEYINPUT116), .ZN(n1021) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1016) );
  XNOR2_X1 U1098 ( .A(G160), .B(G2084), .ZN(n1014) );
  XOR2_X1 U1099 ( .A(G2090), .B(G162), .Z(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1101 ( .A(KEYINPUT51), .B(n1012), .Z(n1013) );
  NAND2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(KEYINPUT115), .B(n1019), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1108 ( .A(KEYINPUT52), .B(n1024), .ZN(n1026) );
  NAND2_X1 U1109 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1110 ( .A1(n1027), .A2(G29), .ZN(n1028) );
  XNOR2_X1 U1111 ( .A(KEYINPUT118), .B(n1028), .ZN(n1029) );
  NAND2_X1 U1112 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1113 ( .A(n1031), .B(KEYINPUT127), .ZN(n1032) );
  XNOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1032), .ZN(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

