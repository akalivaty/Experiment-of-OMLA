//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n844, new_n845, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961;
  AOI21_X1  g000(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT90), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT91), .ZN(new_n205));
  XNOR2_X1  g004(.A(G71gat), .B(G78gat), .ZN(new_n206));
  INV_X1    g005(.A(G64gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G57gat), .ZN(new_n208));
  INV_X1    g007(.A(G57gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G64gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND4_X1  g010(.A1(new_n204), .A2(new_n205), .A3(new_n206), .A4(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G71gat), .A2(G78gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT9), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(new_n203), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n202), .A2(KEYINPUT90), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n216), .A2(new_n211), .A3(new_n206), .A4(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT91), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n216), .A2(new_n211), .A3(new_n217), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT89), .ZN(new_n221));
  OR3_X1    g020(.A1(new_n221), .A2(G71gat), .A3(G78gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n221), .B1(G71gat), .B2(G78gat), .ZN(new_n223));
  AND3_X1   g022(.A1(new_n222), .A2(new_n223), .A3(new_n213), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n212), .A2(new_n219), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OR3_X1    g024(.A1(new_n225), .A2(KEYINPUT93), .A3(KEYINPUT21), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT93), .B1(new_n225), .B2(KEYINPUT21), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G211gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT16), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(G1gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(G1gat), .B2(new_n231), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G8gat), .ZN(new_n235));
  INV_X1    g034(.A(G8gat), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n233), .B(new_n236), .C1(G1gat), .C2(new_n231), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n224), .A2(new_n220), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n218), .A2(KEYINPUT91), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n218), .A2(KEYINPUT91), .ZN(new_n242));
  OAI211_X1 g041(.A(KEYINPUT21), .B(new_n240), .C1(new_n241), .C2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G183gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n239), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n244), .B1(new_n239), .B2(new_n243), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT20), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n247), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT20), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n250), .A3(new_n245), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n252));
  AND3_X1   g051(.A1(new_n248), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n252), .B1(new_n248), .B2(new_n251), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n230), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(G127gat), .B(G155gat), .Z(new_n256));
  NAND2_X1  g055(.A1(G231gat), .A2(G233gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n252), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n250), .B1(new_n249), .B2(new_n245), .ZN(new_n260));
  NOR3_X1   g059(.A1(new_n246), .A2(KEYINPUT20), .A3(new_n247), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n228), .B(G211gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n248), .A2(new_n251), .A3(new_n252), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  AND3_X1   g064(.A1(new_n255), .A2(new_n258), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n258), .B1(new_n255), .B2(new_n265), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(G134gat), .B(G162gat), .Z(new_n269));
  AOI21_X1  g068(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n271), .B(KEYINPUT98), .Z(new_n272));
  NAND3_X1  g071(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(G99gat), .A2(G106gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT94), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT94), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n276), .A2(G99gat), .A3(G106gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n275), .A2(new_n277), .A3(KEYINPUT8), .ZN(new_n278));
  NAND2_X1  g077(.A1(G85gat), .A2(G92gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT7), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT7), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n281), .A2(G85gat), .A3(G92gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  OR2_X1    g082(.A1(G85gat), .A2(G92gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n278), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(G99gat), .B(G106gat), .Z(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n285), .B(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT84), .ZN(new_n289));
  INV_X1    g088(.A(G50gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n289), .B1(new_n290), .B2(G43gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT15), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G29gat), .A2(G36gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT14), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(G29gat), .B2(G36gat), .ZN(new_n296));
  INV_X1    g095(.A(G29gat), .ZN(new_n297));
  INV_X1    g096(.A(G36gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT14), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n293), .A2(new_n294), .A3(new_n296), .A4(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G43gat), .B(G50gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n296), .A3(new_n294), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n292), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n300), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G43gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G50gat), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT15), .B1(new_n306), .B2(new_n289), .ZN(new_n307));
  OR3_X1    g106(.A1(new_n302), .A2(new_n307), .A3(new_n301), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT97), .ZN(new_n310));
  XNOR2_X1  g109(.A(G190gat), .B(G218gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n311), .B(KEYINPUT96), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n288), .A2(new_n309), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT85), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT17), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(KEYINPUT85), .A2(KEYINPUT17), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n309), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n304), .A2(new_n308), .A3(new_n314), .A4(new_n315), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n285), .B(new_n286), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n322), .A2(KEYINPUT95), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT95), .B1(new_n322), .B2(new_n323), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n273), .B(new_n313), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n312), .A2(new_n310), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n326), .A2(new_n327), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n272), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n330), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n271), .A2(KEYINPUT98), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n333), .A3(new_n328), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT99), .B1(new_n268), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT99), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n335), .B(new_n338), .C1(new_n266), .C2(new_n267), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G230gat), .A2(G233gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT100), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n285), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n240), .B(new_n343), .C1(new_n241), .C2(new_n242), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n288), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n225), .A2(new_n323), .A3(new_n343), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT10), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n225), .A2(new_n288), .A3(KEYINPUT10), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n341), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G120gat), .B(G148gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(G176gat), .B(G204gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n345), .A2(new_n346), .A3(G230gat), .A4(G233gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n350), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n353), .A2(KEYINPUT101), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n341), .B(KEYINPUT102), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n358), .B1(new_n347), .B2(new_n349), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n357), .B1(new_n359), .B2(new_n355), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n353), .A2(KEYINPUT101), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n360), .A2(KEYINPUT103), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT103), .B1(new_n360), .B2(new_n361), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n356), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n340), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G228gat), .A2(G233gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(G218gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n229), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G211gat), .A2(G218gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT67), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n370), .A2(KEYINPUT67), .A3(new_n371), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OR2_X1    g175(.A1(KEYINPUT66), .A2(KEYINPUT22), .ZN(new_n377));
  NAND2_X1  g176(.A1(KEYINPUT66), .A2(KEYINPUT22), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n371), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G197gat), .B(G204gat), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT68), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n376), .B(new_n381), .Z(new_n382));
  XOR2_X1   g181(.A(G155gat), .B(G162gat), .Z(new_n383));
  INV_X1    g182(.A(KEYINPUT71), .ZN(new_n384));
  INV_X1    g183(.A(G141gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n385), .A2(G148gat), .ZN(new_n386));
  INV_X1    g185(.A(G148gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n387), .A2(G141gat), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n384), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT2), .ZN(new_n390));
  OR2_X1    g189(.A1(new_n390), .A2(KEYINPUT72), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n387), .A2(G141gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n385), .A2(G148gat), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT71), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n390), .A2(KEYINPUT72), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n389), .A2(new_n391), .A3(new_n394), .A4(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n390), .B1(G155gat), .B2(G162gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n397), .A2(KEYINPUT73), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n398), .A2(new_n383), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n397), .A2(KEYINPUT73), .B1(new_n392), .B2(new_n393), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n383), .A2(new_n396), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT29), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT29), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT3), .B1(new_n382), .B2(new_n404), .ZN(new_n405));
  OAI221_X1 g204(.A(new_n368), .B1(new_n382), .B2(new_n403), .C1(new_n405), .C2(new_n401), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT80), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n403), .A2(new_n382), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n379), .A2(new_n380), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n376), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n374), .A2(new_n379), .A3(new_n375), .A4(new_n380), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n404), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n401), .B1(new_n412), .B2(new_n402), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n407), .B(new_n367), .C1(new_n408), .C2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n412), .A2(new_n402), .ZN(new_n416));
  OAI22_X1  g215(.A1(new_n416), .A2(new_n401), .B1(new_n403), .B2(new_n382), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n407), .B1(new_n417), .B2(new_n367), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n406), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G78gat), .B(G106gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT31), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT79), .B(G50gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT81), .B(G22gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n419), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n406), .B(new_n425), .C1(new_n415), .C2(new_n418), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT36), .ZN(new_n431));
  XOR2_X1   g230(.A(KEYINPUT64), .B(KEYINPUT28), .Z(new_n432));
  INV_X1    g231(.A(G190gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT27), .B(G183gat), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  AND2_X1   g234(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n436));
  NOR2_X1   g235(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n433), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(KEYINPUT64), .A3(KEYINPUT28), .ZN(new_n439));
  NAND2_X1  g238(.A1(G183gat), .A2(G190gat), .ZN(new_n440));
  OR3_X1    g239(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(G169gat), .A2(G176gat), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n435), .A2(new_n439), .A3(new_n440), .A4(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT23), .ZN(new_n446));
  INV_X1    g245(.A(G169gat), .ZN(new_n447));
  INV_X1    g246(.A(G176gat), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n244), .A2(new_n433), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(KEYINPUT24), .A3(new_n440), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n440), .A2(KEYINPUT24), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n451), .A2(new_n453), .A3(new_n455), .A4(new_n443), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT25), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n454), .B1(new_n450), .B2(new_n449), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT25), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n458), .A2(new_n459), .A3(new_n443), .A4(new_n453), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  XOR2_X1   g260(.A(G127gat), .B(G134gat), .Z(new_n462));
  NOR2_X1   g261(.A1(new_n462), .A2(KEYINPUT1), .ZN(new_n463));
  AND2_X1   g262(.A1(KEYINPUT65), .A2(G120gat), .ZN(new_n464));
  NOR2_X1   g263(.A1(KEYINPUT65), .A2(G120gat), .ZN(new_n465));
  OAI21_X1  g264(.A(G113gat), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(G120gat), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n466), .B1(G113gat), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT1), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n467), .A2(G113gat), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n467), .A2(G113gat), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n463), .A2(new_n468), .B1(new_n472), .B2(new_n462), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n461), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(G227gat), .A2(G233gat), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n473), .A2(new_n445), .A3(new_n457), .A4(new_n460), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n476), .B1(new_n475), .B2(new_n477), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT32), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT34), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT34), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n479), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G15gat), .B(G43gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(G71gat), .B(G99gat), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n486), .B(new_n487), .Z(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(new_n480), .B2(KEYINPUT33), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  OR3_X1    g289(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT34), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n491), .A2(new_n482), .A3(new_n478), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n485), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n490), .B1(new_n485), .B2(new_n492), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n431), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n485), .A2(new_n492), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n489), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n498), .A2(KEYINPUT36), .A3(new_n493), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n430), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT82), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n396), .A2(new_n383), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n399), .A2(new_n400), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n474), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT76), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n473), .A2(new_n502), .A3(new_n503), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G225gat), .A2(G233gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT74), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n504), .A2(new_n474), .A3(KEYINPUT76), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n508), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT4), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n473), .A2(new_n502), .A3(new_n513), .A4(new_n503), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT75), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT75), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n401), .A2(new_n517), .A3(new_n513), .A4(new_n473), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT3), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n401), .A2(new_n402), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n521), .A3(new_n474), .ZN(new_n522));
  INV_X1    g321(.A(new_n510), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n512), .B(KEYINPUT5), .C1(new_n519), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n516), .A2(new_n514), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(new_n522), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(KEYINPUT78), .B(G1gat), .Z(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G57gat), .B(G85gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(G29gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n532), .B(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n529), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT6), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n525), .A2(new_n535), .A3(new_n528), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n535), .B1(new_n525), .B2(new_n528), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT6), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n501), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n461), .A2(G226gat), .A3(G233gat), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n461), .A2(new_n404), .B1(G226gat), .B2(G233gat), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n382), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n461), .A2(new_n404), .ZN(new_n547));
  NAND2_X1  g346(.A1(G226gat), .A2(G233gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n382), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n461), .A2(G226gat), .A3(G233gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n546), .A2(new_n552), .A3(KEYINPUT69), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT69), .B1(new_n546), .B2(new_n552), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT37), .ZN(new_n555));
  NOR3_X1   g354(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n546), .A2(new_n552), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n555), .ZN(new_n558));
  XNOR2_X1  g357(.A(G8gat), .B(G36gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(G64gat), .B(G92gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT38), .B1(new_n556), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n561), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n557), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT70), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n557), .A2(KEYINPUT70), .A3(new_n564), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n564), .B1(new_n557), .B2(new_n555), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT38), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n546), .A2(new_n552), .A3(KEYINPUT37), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n563), .A2(new_n569), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n542), .A2(new_n501), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NOR3_X1   g375(.A1(new_n543), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT30), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n567), .A2(new_n578), .A3(new_n568), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n553), .A2(new_n554), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n561), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n557), .A2(KEYINPUT30), .A3(new_n564), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n523), .B1(new_n526), .B2(new_n522), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n510), .B1(new_n508), .B2(new_n511), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT39), .ZN(new_n587));
  OR3_X1    g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n536), .B1(new_n585), .B2(new_n587), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT40), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n588), .A2(KEYINPUT40), .A3(new_n589), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(new_n593), .A3(new_n537), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n584), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n500), .B1(new_n577), .B2(new_n595), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n429), .A2(new_n498), .A3(new_n493), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n597), .B(new_n584), .C1(new_n543), .C2(new_n576), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT35), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AND3_X1   g399(.A1(new_n525), .A2(new_n535), .A3(new_n528), .ZN(new_n601));
  NOR3_X1   g400(.A1(new_n601), .A2(new_n541), .A3(KEYINPUT6), .ZN(new_n602));
  INV_X1    g401(.A(new_n542), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n429), .B1(new_n496), .B2(new_n499), .ZN(new_n606));
  AND4_X1   g405(.A1(KEYINPUT35), .A2(new_n429), .A3(new_n498), .A4(new_n493), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n605), .B(new_n584), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n596), .A2(new_n600), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT83), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n584), .A2(new_n594), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT82), .B1(new_n602), .B2(new_n603), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n572), .A2(new_n571), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n567), .B(new_n568), .C1(new_n562), .C2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n580), .A2(KEYINPUT37), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n570), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n615), .B1(new_n617), .B2(KEYINPUT38), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n613), .A2(new_n618), .A3(new_n575), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n612), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n620), .A2(new_n500), .B1(new_n599), .B2(new_n598), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n621), .A2(KEYINPUT83), .A3(new_n608), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n366), .B1(new_n611), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT86), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n624), .B1(new_n322), .B2(new_n239), .ZN(new_n625));
  AOI211_X1 g424(.A(KEYINPUT86), .B(new_n238), .C1(new_n320), .C2(new_n321), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(G229gat), .A2(G233gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n238), .A2(new_n309), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n627), .A2(KEYINPUT18), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  AOI211_X1 g429(.A(new_n316), .B(new_n318), .C1(new_n304), .C2(new_n308), .ZN(new_n631));
  INV_X1    g430(.A(new_n321), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n239), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT86), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n322), .A2(new_n624), .A3(new_n239), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n634), .A2(new_n628), .A3(new_n629), .A4(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT18), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT87), .B1(new_n238), .B2(new_n309), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(new_n629), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n628), .B(KEYINPUT13), .Z(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n630), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G113gat), .B(G141gat), .ZN(new_n644));
  INV_X1    g443(.A(G197gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT11), .B(G169gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n630), .A2(new_n638), .A3(new_n649), .A4(new_n642), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(KEYINPUT88), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT88), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n643), .A2(new_n654), .A3(new_n650), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n623), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n604), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g460(.A1(new_n232), .A2(new_n236), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n623), .A2(new_n657), .A3(new_n583), .A4(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT42), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n232), .A2(new_n236), .ZN(new_n665));
  OR3_X1    g464(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(G8gat), .B1(new_n658), .B2(new_n584), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n664), .B1(new_n663), .B2(new_n665), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n666), .A2(KEYINPUT104), .A3(new_n667), .A4(new_n668), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(G1325gat));
  NOR2_X1   g472(.A1(new_n494), .A2(new_n495), .ZN(new_n674));
  AOI21_X1  g473(.A(G15gat), .B1(new_n659), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  INV_X1    g477(.A(new_n496), .ZN(new_n679));
  INV_X1    g478(.A(new_n499), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(G15gat), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT106), .Z(new_n683));
  AOI22_X1  g482(.A1(new_n677), .A2(new_n678), .B1(new_n659), .B2(new_n683), .ZN(G1326gat));
  NOR2_X1   g483(.A1(new_n658), .A2(new_n429), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT43), .B(G22gat), .Z(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1327gat));
  AOI21_X1  g486(.A(new_n335), .B1(new_n611), .B2(new_n622), .ZN(new_n688));
  INV_X1    g487(.A(new_n268), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n689), .A2(new_n656), .A3(new_n364), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n691), .A2(new_n297), .A3(new_n604), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT107), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT107), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n691), .A2(new_n694), .A3(new_n297), .A4(new_n604), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT45), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT83), .B1(new_n621), .B2(new_n608), .ZN(new_n699));
  AND4_X1   g498(.A1(KEYINPUT83), .A2(new_n596), .A3(new_n600), .A4(new_n608), .ZN(new_n700));
  OAI211_X1 g499(.A(KEYINPUT44), .B(new_n336), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n609), .A2(new_n336), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n690), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT108), .B1(new_n706), .B2(new_n605), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n705), .A2(new_n708), .A3(new_n604), .A4(new_n690), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n707), .A2(new_n709), .A3(G29gat), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n693), .A2(KEYINPUT45), .A3(new_n695), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n698), .A2(new_n710), .A3(new_n711), .ZN(G1328gat));
  NAND3_X1  g511(.A1(new_n691), .A2(new_n298), .A3(new_n583), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n713), .B(KEYINPUT46), .Z(new_n714));
  OAI21_X1  g513(.A(G36gat), .B1(new_n706), .B2(new_n584), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(G1329gat));
  NAND4_X1  g515(.A1(new_n701), .A2(new_n681), .A3(new_n704), .A4(new_n690), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G43gat), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n691), .A2(new_n305), .A3(new_n674), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n720), .A2(KEYINPUT109), .A3(KEYINPUT47), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT47), .B1(new_n720), .B2(KEYINPUT109), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(G1330gat));
  NAND4_X1  g522(.A1(new_n701), .A2(new_n430), .A3(new_n704), .A4(new_n690), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G50gat), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n430), .A2(new_n290), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT110), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n691), .A2(new_n727), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n725), .B(new_n728), .C1(KEYINPUT111), .C2(KEYINPUT48), .ZN(new_n729));
  NAND2_X1  g528(.A1(KEYINPUT111), .A2(KEYINPUT48), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1331gat));
  AOI21_X1  g530(.A(new_n657), .B1(new_n621), .B2(new_n608), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n340), .A2(new_n364), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n605), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(new_n209), .ZN(G1332gat));
  INV_X1    g535(.A(new_n734), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n583), .ZN(new_n738));
  AND2_X1   g537(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n739));
  OR3_X1    g538(.A1(new_n738), .A2(KEYINPUT112), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT112), .B1(new_n738), .B2(new_n739), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n742), .B(new_n744), .ZN(G1333gat));
  INV_X1    g544(.A(new_n681), .ZN(new_n746));
  OAI21_X1  g545(.A(G71gat), .B1(new_n734), .B2(new_n746), .ZN(new_n747));
  OR2_X1    g546(.A1(new_n734), .A2(G71gat), .ZN(new_n748));
  INV_X1    g547(.A(new_n674), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g550(.A1(new_n737), .A2(new_n430), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g552(.A1(new_n689), .A2(new_n657), .A3(new_n365), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n705), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(G85gat), .B1(new_n755), .B2(new_n605), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n689), .A2(new_n657), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n609), .A2(new_n336), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n609), .A2(KEYINPUT51), .A3(new_n336), .A4(new_n757), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n758), .A2(KEYINPUT113), .A3(new_n759), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n763), .A2(KEYINPUT114), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT114), .B1(new_n763), .B2(new_n764), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n364), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n605), .A2(G85gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n756), .B1(new_n767), .B2(new_n768), .ZN(G1336gat));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n705), .A2(new_n583), .A3(new_n754), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n760), .A2(new_n762), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n365), .A2(new_n584), .A3(G92gat), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n771), .A2(G92gat), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n771), .A2(G92gat), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n763), .A2(new_n764), .A3(new_n773), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n770), .ZN(new_n777));
  OAI22_X1  g576(.A1(new_n770), .A2(new_n774), .B1(new_n775), .B2(new_n777), .ZN(G1337gat));
  OAI21_X1  g577(.A(KEYINPUT115), .B1(new_n755), .B2(new_n746), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n705), .A2(new_n780), .A3(new_n681), .A4(new_n754), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(new_n781), .A3(G99gat), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n749), .A2(G99gat), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n767), .B2(new_n783), .ZN(G1338gat));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n701), .A2(new_n430), .A3(new_n704), .A4(new_n754), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G106gat), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n365), .A2(G106gat), .A3(new_n429), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n763), .A2(new_n764), .A3(new_n789), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n772), .A2(new_n789), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n788), .B1(new_n787), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n785), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n786), .A2(G106gat), .B1(new_n772), .B2(new_n789), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n795), .B(KEYINPUT116), .C1(new_n788), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n794), .A2(new_n797), .ZN(G1339gat));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n799), .B(new_n358), .C1(new_n347), .C2(new_n349), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n347), .A2(new_n349), .A3(new_n358), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n350), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT10), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n344), .A2(new_n288), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n323), .B1(new_n225), .B2(new_n343), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n358), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n807), .A2(new_n802), .A3(new_n348), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT54), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n353), .B(new_n800), .C1(new_n803), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT55), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n807), .A2(new_n348), .A3(new_n808), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT117), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n814), .A2(KEYINPUT54), .A3(new_n350), .A4(new_n809), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n815), .A2(new_n816), .A3(new_n353), .A4(new_n800), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n818), .A2(new_n653), .A3(new_n655), .A4(new_n356), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n628), .B1(new_n627), .B2(new_n629), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n640), .A2(new_n641), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n648), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n652), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n364), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n336), .B1(new_n819), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n356), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n826), .B1(new_n812), .B2(new_n817), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n336), .A2(new_n827), .A3(new_n823), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n268), .B1(new_n825), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n337), .A2(new_n656), .A3(new_n339), .A4(new_n365), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n832), .A2(new_n597), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n605), .A2(new_n583), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(new_n656), .ZN(new_n836));
  XOR2_X1   g635(.A(KEYINPUT118), .B(G113gat), .Z(new_n837));
  XNOR2_X1  g636(.A(new_n836), .B(new_n837), .ZN(G1340gat));
  INV_X1    g637(.A(new_n835), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n364), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(G120gat), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n464), .A2(new_n465), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n841), .B1(new_n842), .B2(new_n840), .ZN(G1341gat));
  NOR2_X1   g642(.A1(new_n835), .A2(new_n268), .ZN(new_n844));
  NOR2_X1   g643(.A1(KEYINPUT119), .A2(G127gat), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n844), .B(new_n845), .ZN(G1342gat));
  NAND2_X1  g645(.A1(new_n839), .A2(new_n336), .ZN(new_n847));
  OR3_X1    g646(.A1(new_n847), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(G134gat), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT56), .B1(new_n847), .B2(G134gat), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(G1343gat));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n852), .B1(new_n832), .B2(new_n430), .ZN(new_n853));
  AOI211_X1 g652(.A(KEYINPUT57), .B(new_n429), .C1(new_n830), .C2(new_n831), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n746), .A2(new_n834), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n385), .B1(new_n856), .B2(new_n657), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n819), .A2(new_n824), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n335), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n689), .B1(new_n859), .B2(new_n828), .ZN(new_n860));
  INV_X1    g659(.A(new_n831), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n604), .B(new_n606), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT121), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n656), .A2(G141gat), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n832), .A2(KEYINPUT121), .A3(new_n604), .A4(new_n606), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n864), .A2(new_n584), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT122), .B1(new_n857), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n832), .A2(new_n430), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT57), .ZN(new_n872));
  INV_X1    g671(.A(new_n855), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n832), .A2(new_n852), .A3(new_n430), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(G141gat), .B1(new_n875), .B2(new_n656), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n876), .A2(new_n877), .A3(new_n868), .A4(new_n867), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n870), .A2(new_n878), .ZN(new_n879));
  NOR4_X1   g678(.A1(new_n862), .A2(G141gat), .A3(new_n656), .A4(new_n583), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n853), .A2(new_n854), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT120), .B1(new_n881), .B2(new_n873), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n883));
  NOR4_X1   g682(.A1(new_n853), .A2(new_n854), .A3(new_n883), .A4(new_n855), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n657), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n880), .B1(new_n885), .B2(G141gat), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n879), .B1(new_n886), .B2(new_n868), .ZN(G1344gat));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n864), .A2(new_n584), .A3(new_n866), .ZN(new_n889));
  AOI211_X1 g688(.A(new_n888), .B(G148gat), .C1(new_n889), .C2(new_n364), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n831), .A2(KEYINPUT123), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n831), .A2(KEYINPUT123), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n830), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n852), .A3(new_n430), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n894), .A2(new_n364), .A3(new_n872), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(KEYINPUT59), .A3(new_n873), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n875), .A2(new_n883), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n881), .A2(KEYINPUT120), .A3(new_n873), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n365), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n896), .B1(new_n899), .B2(KEYINPUT59), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n890), .B1(new_n900), .B2(G148gat), .ZN(G1345gat));
  AOI21_X1  g700(.A(G155gat), .B1(new_n889), .B2(new_n689), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n882), .A2(new_n884), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n903), .A2(new_n268), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n902), .B1(new_n904), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g704(.A(G162gat), .B1(new_n889), .B2(new_n336), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n903), .A2(new_n335), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g707(.A1(new_n604), .A2(new_n584), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n833), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n447), .A3(new_n657), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n909), .B(KEYINPUT124), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n833), .A2(new_n913), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n914), .A2(new_n657), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n912), .B1(new_n915), .B2(new_n447), .ZN(G1348gat));
  AOI21_X1  g715(.A(G176gat), .B1(new_n911), .B2(new_n364), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n365), .A2(new_n448), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n914), .B2(new_n918), .ZN(G1349gat));
  NAND2_X1  g718(.A1(new_n914), .A2(new_n689), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n689), .A2(new_n434), .ZN(new_n921));
  AOI22_X1  g720(.A1(new_n920), .A2(G183gat), .B1(new_n911), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT60), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n922), .B(new_n923), .ZN(G1350gat));
  NAND3_X1  g723(.A1(new_n911), .A2(new_n433), .A3(new_n336), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n832), .A2(new_n597), .A3(new_n336), .A4(new_n913), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(G190gat), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT125), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n926), .A2(new_n930), .A3(G190gat), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n929), .B1(new_n928), .B2(new_n931), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n925), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI211_X1 g735(.A(KEYINPUT126), .B(new_n925), .C1(new_n932), .C2(new_n933), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1351gat));
  AND2_X1   g737(.A1(new_n913), .A2(new_n746), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n894), .A2(new_n872), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n657), .A2(G197gat), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n832), .A2(new_n606), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n909), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n645), .B1(new_n944), .B2(new_n656), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n942), .A2(KEYINPUT127), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT127), .B1(new_n942), .B2(new_n945), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n946), .A2(new_n947), .ZN(G1352gat));
  NOR3_X1   g747(.A1(new_n944), .A2(G204gat), .A3(new_n365), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT62), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n895), .A2(new_n939), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(G204gat), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1353gat));
  INV_X1    g752(.A(new_n944), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n954), .A2(new_n229), .A3(new_n689), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n894), .A2(new_n689), .A3(new_n872), .A4(new_n939), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  OAI21_X1  g758(.A(G218gat), .B1(new_n940), .B2(new_n335), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n954), .A2(new_n369), .A3(new_n336), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1355gat));
endmodule


