//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT78), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT78), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G104), .ZN(new_n193));
  AOI21_X1  g007(.A(G107), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G107), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G104), .ZN(new_n196));
  OAI211_X1 g010(.A(KEYINPUT81), .B(G101), .C1(new_n194), .C2(new_n196), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n191), .B(new_n193), .C1(KEYINPUT3), .C2(G107), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT3), .A2(G107), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT3), .A2(G107), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n199), .B1(G104), .B2(new_n200), .ZN(new_n201));
  XOR2_X1   g015(.A(KEYINPUT80), .B(G101), .Z(new_n202));
  NAND3_X1  g016(.A1(new_n198), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n197), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n196), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT78), .B(G104), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(G107), .ZN(new_n207));
  AOI21_X1  g021(.A(KEYINPUT81), .B1(new_n207), .B2(G101), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n215), .B1(G143), .B2(new_n210), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n214), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G143), .B(G146), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT67), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AND4_X1   g035(.A1(KEYINPUT67), .A2(new_n220), .A3(new_n211), .A4(new_n213), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n218), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT82), .B1(new_n209), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT81), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n191), .A2(new_n193), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n196), .B1(new_n226), .B2(new_n195), .ZN(new_n227));
  INV_X1    g041(.A(G101), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n225), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n223), .A2(new_n229), .A3(new_n203), .A4(new_n197), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT82), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT68), .B(G128), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n214), .B1(new_n233), .B2(new_n216), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n234), .B1(new_n221), .B2(new_n222), .ZN(new_n235));
  OAI22_X1  g049(.A1(new_n224), .A2(new_n232), .B1(new_n235), .B2(new_n209), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT11), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(KEYINPUT65), .ZN(new_n238));
  INV_X1    g052(.A(G134), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(G137), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(KEYINPUT65), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n238), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(G137), .ZN(new_n243));
  INV_X1    g057(.A(G137), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G134), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT11), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n243), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(G131), .B1(new_n242), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n246), .A2(KEYINPUT11), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n247), .B1(new_n250), .B2(new_n245), .ZN(new_n251));
  INV_X1    g065(.A(G131), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n240), .A2(new_n238), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n251), .A2(new_n252), .A3(new_n243), .A4(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n236), .A2(KEYINPUT12), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT12), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n230), .A2(new_n231), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n197), .A2(new_n203), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n259), .A2(KEYINPUT82), .A3(new_n223), .A4(new_n229), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n220), .A2(new_n211), .A3(new_n213), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n219), .A2(KEYINPUT67), .A3(new_n220), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n217), .A2(KEYINPUT68), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G128), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n263), .A2(new_n264), .B1(new_n270), .B2(new_n214), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n259), .A2(new_n229), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n258), .A2(new_n260), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n255), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n257), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n256), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(G110), .B(G140), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n277), .B(KEYINPUT77), .ZN(new_n278));
  INV_X1    g092(.A(G953), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n279), .A2(G227), .ZN(new_n280));
  XOR2_X1   g094(.A(new_n278), .B(new_n280), .Z(new_n281));
  AOI21_X1  g095(.A(KEYINPUT10), .B1(new_n258), .B2(new_n260), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT83), .B1(new_n204), .B2(new_n208), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT83), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n229), .A2(new_n284), .A3(new_n203), .A4(new_n197), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT10), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n271), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n283), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT0), .A4(G128), .ZN(new_n289));
  OR2_X1    g103(.A1(KEYINPUT0), .A2(G128), .ZN(new_n290));
  NAND2_X1  g104(.A1(KEYINPUT0), .A2(G128), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n289), .B1(new_n219), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n228), .B1(new_n198), .B2(new_n201), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT4), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g111(.A(KEYINPUT4), .B(new_n203), .C1(new_n295), .C2(KEYINPUT79), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n295), .A2(KEYINPUT79), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n294), .B(new_n297), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n288), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n282), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT84), .B1(new_n302), .B2(new_n274), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT84), .ZN(new_n304));
  NOR4_X1   g118(.A1(new_n282), .A2(new_n301), .A3(new_n304), .A4(new_n255), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n276), .B(new_n281), .C1(new_n303), .C2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n255), .B1(new_n282), .B2(new_n301), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n286), .B1(new_n224), .B2(new_n232), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n288), .A2(new_n300), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(new_n274), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n304), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n302), .A2(KEYINPUT84), .A3(new_n274), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n308), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n306), .B1(new_n314), .B2(new_n281), .ZN(new_n315));
  INV_X1    g129(.A(G469), .ZN(new_n316));
  INV_X1    g130(.A(G902), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT85), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n307), .B1(new_n303), .B2(new_n305), .ZN(new_n321));
  INV_X1    g135(.A(new_n281), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(G902), .B1(new_n323), .B2(new_n306), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(KEYINPUT85), .A3(new_n316), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n276), .B1(new_n303), .B2(new_n305), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n322), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n307), .B(new_n281), .C1(new_n303), .C2(new_n305), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(G469), .B1(new_n331), .B2(G902), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n189), .B1(new_n326), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT2), .B(G113), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(G116), .B(G119), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n336), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n244), .A2(G134), .ZN(new_n340));
  OAI21_X1  g154(.A(G131), .B1(new_n340), .B2(new_n240), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n235), .A2(new_n341), .A3(new_n254), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n242), .A2(new_n248), .A3(G131), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n340), .B1(new_n240), .B2(new_n238), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n252), .B1(new_n344), .B2(new_n251), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n294), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(new_n346), .A3(KEYINPUT30), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n293), .B1(new_n249), .B2(new_n254), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n254), .A2(new_n341), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n263), .A2(new_n264), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n349), .A2(KEYINPUT66), .B1(new_n350), .B2(new_n234), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT66), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n254), .A2(new_n352), .A3(new_n341), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n348), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n339), .B(new_n347), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT31), .ZN(new_n357));
  INV_X1    g171(.A(new_n339), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n342), .A2(new_n358), .A3(new_n346), .ZN(new_n359));
  NOR2_X1   g173(.A1(G237), .A2(G953), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G210), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(KEYINPUT27), .ZN(new_n362));
  XNOR2_X1  g176(.A(KEYINPUT26), .B(G101), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n362), .B(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n356), .A2(new_n357), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT69), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT69), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n356), .A2(new_n368), .A3(new_n357), .A4(new_n365), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n254), .A2(new_n341), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n371), .A2(new_n235), .B1(new_n255), .B2(new_n294), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT28), .B1(new_n372), .B2(new_n358), .ZN(new_n373));
  AND4_X1   g187(.A1(KEYINPUT28), .A2(new_n342), .A3(new_n358), .A4(new_n346), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n349), .A2(KEYINPUT66), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n235), .A3(new_n353), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n346), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n339), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n364), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n357), .B1(new_n356), .B2(new_n365), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n370), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(G472), .A2(G902), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT32), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G472), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n356), .A2(new_n359), .ZN(new_n387));
  INV_X1    g201(.A(new_n364), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT70), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(KEYINPUT70), .A3(new_n388), .ZN(new_n392));
  INV_X1    g206(.A(new_n374), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT28), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n359), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n379), .A2(new_n393), .A3(new_n364), .A4(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT29), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n391), .A2(new_n392), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT71), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n372), .A2(new_n401), .A3(new_n358), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n359), .A2(KEYINPUT71), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n402), .B(new_n403), .C1(new_n358), .C2(new_n372), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n373), .B1(new_n404), .B2(KEYINPUT28), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n388), .A2(new_n397), .ZN(new_n406));
  AOI21_X1  g220(.A(G902), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n386), .B1(new_n400), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT32), .ZN(new_n409));
  INV_X1    g223(.A(new_n384), .ZN(new_n410));
  AOI211_X1 g224(.A(new_n409), .B(new_n410), .C1(new_n370), .C2(new_n382), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n385), .A2(new_n408), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT76), .ZN(new_n413));
  INV_X1    g227(.A(G217), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n414), .B1(G234), .B2(new_n317), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT74), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n265), .A2(new_n267), .A3(G119), .ZN(new_n418));
  INV_X1    g232(.A(G119), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G128), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT72), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT72), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n418), .A2(new_n423), .A3(new_n420), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT24), .B(G110), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n422), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT16), .ZN(new_n428));
  INV_X1    g242(.A(G140), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n429), .A3(G125), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(G125), .ZN(new_n431));
  INV_X1    g245(.A(G125), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G140), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n430), .B1(new_n434), .B2(new_n428), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n210), .ZN(new_n436));
  OAI211_X1 g250(.A(G146), .B(new_n430), .C1(new_n434), .C2(new_n428), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT23), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n439), .B1(new_n419), .B2(G128), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n420), .B(new_n440), .C1(new_n418), .C2(new_n439), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G110), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n427), .A2(new_n438), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT73), .B1(new_n434), .B2(G146), .ZN(new_n445));
  XNOR2_X1  g259(.A(G125), .B(G140), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT73), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(new_n210), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n437), .ZN(new_n450));
  OR2_X1    g264(.A1(new_n441), .A2(G110), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n418), .A2(new_n423), .A3(new_n420), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n423), .B1(new_n418), .B2(new_n420), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n425), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n450), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n417), .B1(new_n444), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n426), .B1(new_n422), .B2(new_n424), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n441), .A2(G110), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n443), .B(KEYINPUT74), .C1(new_n459), .C2(new_n450), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT22), .B(G137), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n279), .A2(G221), .A3(G234), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n461), .B(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(KEYINPUT75), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n456), .A2(new_n460), .A3(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n443), .B(new_n463), .C1(new_n459), .C2(new_n450), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n317), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT25), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT25), .A4(new_n317), .ZN(new_n470));
  AOI211_X1 g284(.A(new_n413), .B(new_n416), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n469), .A2(new_n470), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n415), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n413), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n465), .A2(new_n466), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n415), .A2(G902), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n472), .B(new_n475), .C1(new_n476), .C2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n412), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n212), .A2(KEYINPUT13), .A3(G128), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT96), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n233), .A2(G143), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n217), .A2(G143), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n482), .B(new_n483), .C1(KEYINPUT13), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G134), .ZN(new_n486));
  INV_X1    g300(.A(G122), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n487), .A2(KEYINPUT95), .A3(G116), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT95), .B1(new_n487), .B2(G116), .ZN(new_n489));
  OAI22_X1  g303(.A1(new_n488), .A2(new_n489), .B1(G116), .B2(new_n487), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(G107), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n212), .A2(G128), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n483), .A2(new_n239), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n486), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT97), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT97), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n486), .A2(new_n491), .A3(new_n496), .A4(new_n493), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n483), .A2(new_n492), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G134), .ZN(new_n499));
  INV_X1    g313(.A(new_n490), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n195), .A2(KEYINPUT14), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n499), .A2(new_n493), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT14), .B1(new_n488), .B2(new_n489), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n490), .A2(new_n503), .A3(G107), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n495), .A2(new_n497), .A3(new_n505), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n187), .A2(new_n414), .A3(G953), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n494), .A2(KEYINPUT97), .B1(new_n502), .B2(new_n504), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n497), .A3(new_n507), .ZN(new_n511));
  AOI21_X1  g325(.A(G902), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G478), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(KEYINPUT15), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n512), .B(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n360), .A2(G214), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT91), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n517), .A3(new_n212), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n360), .B(G214), .C1(KEYINPUT91), .C2(G143), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G131), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT17), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n518), .A2(new_n252), .A3(new_n519), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n252), .B1(new_n518), .B2(new_n519), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT17), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n524), .A2(new_n436), .A3(new_n437), .A4(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n434), .A2(G146), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n518), .A2(new_n519), .ZN(new_n529));
  NAND2_X1  g343(.A1(KEYINPUT92), .A2(KEYINPUT18), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n449), .A2(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n518), .A2(new_n252), .A3(new_n519), .ZN(new_n532));
  OAI211_X1 g346(.A(KEYINPUT92), .B(KEYINPUT18), .C1(new_n532), .C2(new_n525), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(G113), .B(G122), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(new_n190), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n527), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n536), .B1(new_n527), .B2(new_n534), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n317), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT94), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(KEYINPUT94), .B(new_n317), .C1(new_n537), .C2(new_n538), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(G475), .A3(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(G475), .A2(G902), .ZN(new_n544));
  AND2_X1   g358(.A1(KEYINPUT93), .A2(KEYINPUT19), .ZN(new_n545));
  NOR2_X1   g359(.A1(KEYINPUT93), .A2(KEYINPUT19), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n446), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n547), .B1(new_n446), .B2(new_n546), .ZN(new_n548));
  OAI221_X1 g362(.A(new_n437), .B1(new_n548), .B2(G146), .C1(new_n525), .C2(new_n532), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n536), .B1(new_n534), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n544), .B1(new_n537), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT20), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT20), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n553), .B(new_n544), .C1(new_n537), .C2(new_n550), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n543), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n279), .A2(G952), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(G234), .B2(G237), .ZN(new_n558));
  AOI211_X1 g372(.A(new_n317), .B(new_n279), .C1(G234), .C2(G237), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT21), .B(G898), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n515), .A2(new_n556), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(G210), .B1(G237), .B2(G902), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n419), .A2(G116), .ZN(new_n566));
  INV_X1    g380(.A(G116), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G119), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n568), .A3(KEYINPUT5), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT87), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n336), .A2(KEYINPUT87), .A3(KEYINPUT5), .ZN(new_n572));
  INV_X1    g386(.A(G113), .ZN(new_n573));
  INV_X1    g387(.A(new_n566), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT5), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n571), .A2(new_n572), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n338), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n259), .A2(new_n229), .A3(new_n578), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n576), .A2(new_n569), .B1(new_n335), .B2(new_n336), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n580), .B1(new_n204), .B2(new_n208), .ZN(new_n581));
  XNOR2_X1  g395(.A(G110), .B(G122), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(KEYINPUT8), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n579), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n350), .A2(new_n432), .A3(new_n234), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n293), .A2(G125), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(G224), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(G953), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT88), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n589), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n587), .A2(new_n592), .B1(KEYINPUT7), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(KEYINPUT7), .ZN(new_n595));
  AOI211_X1 g409(.A(new_n591), .B(new_n595), .C1(new_n585), .C2(new_n586), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n584), .B(KEYINPUT89), .C1(new_n594), .C2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n283), .A2(new_n285), .A3(new_n580), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n339), .B(new_n297), .C1(new_n298), .C2(new_n299), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n582), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n587), .A2(new_n590), .A3(KEYINPUT7), .A4(new_n593), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n214), .A2(new_n291), .A3(new_n290), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n432), .B1(new_n603), .B2(new_n289), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n271), .B2(new_n432), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n595), .B1(new_n605), .B2(new_n591), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(KEYINPUT89), .B1(new_n607), .B2(new_n584), .ZN(new_n608));
  OAI211_X1 g422(.A(KEYINPUT90), .B(new_n317), .C1(new_n601), .C2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n598), .A2(new_n599), .ZN(new_n610));
  INV_X1    g424(.A(new_n582), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(KEYINPUT6), .A3(new_n600), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n605), .B(KEYINPUT86), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n589), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT86), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n605), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n593), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT6), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n610), .A2(new_n620), .A3(new_n611), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n613), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n609), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n584), .B1(new_n594), .B2(new_n596), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT89), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n626), .A2(new_n600), .A3(new_n597), .ZN(new_n627));
  AOI21_X1  g441(.A(KEYINPUT90), .B1(new_n627), .B2(new_n317), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n565), .B1(new_n623), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n317), .B1(new_n601), .B2(new_n608), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT90), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n632), .A2(new_n564), .A3(new_n622), .A4(new_n609), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(G214), .B1(G237), .B2(G902), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n563), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n333), .A2(new_n480), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT98), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(new_n202), .ZN(G3));
  NAND2_X1  g453(.A1(new_n383), .A2(new_n317), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(G472), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n640), .B(new_n642), .Z(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n479), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n333), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n645), .B(KEYINPUT100), .Z(new_n646));
  NOR2_X1   g460(.A1(new_n513), .A2(new_n317), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n512), .B2(new_n513), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n510), .A2(new_n497), .A3(new_n507), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n507), .B1(new_n510), .B2(new_n497), .ZN(new_n650));
  OAI21_X1  g464(.A(KEYINPUT33), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT33), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n509), .A2(new_n652), .A3(new_n511), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n651), .A2(G478), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n655), .A2(new_n556), .A3(new_n561), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n629), .A2(KEYINPUT101), .A3(new_n633), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT101), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n658), .B(new_n565), .C1(new_n623), .C2(new_n628), .ZN(new_n659));
  AND4_X1   g473(.A1(new_n635), .A2(new_n656), .A3(new_n657), .A4(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n646), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT34), .B(G104), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G6));
  NAND2_X1  g478(.A1(new_n543), .A2(new_n555), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n561), .B(KEYINPUT102), .Z(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n515), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  AND4_X1   g482(.A1(new_n635), .A2(new_n668), .A3(new_n657), .A4(new_n659), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n646), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT35), .B(G107), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  AOI21_X1  g487(.A(KEYINPUT76), .B1(new_n473), .B2(new_n415), .ZN(new_n674));
  OR2_X1    g488(.A1(new_n464), .A2(KEYINPUT36), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n456), .A2(new_n460), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n675), .B1(new_n456), .B2(new_n460), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n477), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n674), .A2(new_n471), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n643), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n333), .A2(new_n682), .A3(new_n636), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT103), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT37), .B(G110), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G12));
  XOR2_X1   g500(.A(new_n558), .B(KEYINPUT104), .Z(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(G900), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n688), .B1(new_n689), .B2(new_n559), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n515), .A2(new_n665), .A3(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n691), .A2(new_n657), .A3(new_n635), .A4(new_n659), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n692), .A2(new_n412), .A3(new_n681), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n333), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G128), .ZN(G30));
  NOR2_X1   g509(.A1(new_n385), .A2(new_n411), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n317), .B1(new_n404), .B2(new_n364), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n388), .B1(new_n356), .B2(new_n359), .ZN(new_n698));
  OAI21_X1  g512(.A(G472), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n634), .B(KEYINPUT38), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n515), .A2(new_n556), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n681), .A2(new_n635), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n701), .B1(new_n703), .B2(KEYINPUT105), .ZN(new_n704));
  AOI211_X1 g518(.A(new_n700), .B(new_n704), .C1(KEYINPUT105), .C2(new_n703), .ZN(new_n705));
  XOR2_X1   g519(.A(new_n690), .B(KEYINPUT39), .Z(new_n706));
  NAND2_X1  g520(.A1(new_n333), .A2(new_n706), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n707), .A2(KEYINPUT40), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(KEYINPUT40), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n705), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G143), .ZN(G45));
  NOR2_X1   g525(.A1(new_n655), .A2(new_n556), .ZN(new_n712));
  INV_X1    g526(.A(new_n690), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n412), .A2(new_n681), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(KEYINPUT85), .B1(new_n324), .B2(new_n316), .ZN(new_n716));
  AND4_X1   g530(.A1(KEYINPUT85), .A2(new_n315), .A3(new_n316), .A4(new_n317), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n332), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n657), .A2(new_n635), .A3(new_n659), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n715), .A2(new_n718), .A3(new_n188), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G146), .ZN(G48));
  OAI21_X1  g535(.A(new_n188), .B1(new_n324), .B2(new_n316), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n320), .B2(new_n325), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n480), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n661), .ZN(new_n725));
  XOR2_X1   g539(.A(KEYINPUT41), .B(G113), .Z(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G15));
  NOR2_X1   g541(.A1(new_n724), .A2(new_n670), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(new_n567), .ZN(G18));
  INV_X1    g543(.A(new_n722), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n719), .A2(new_n326), .A3(new_n730), .ZN(new_n731));
  AOI211_X1 g545(.A(new_n381), .B(new_n380), .C1(new_n367), .C2(new_n369), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n409), .B1(new_n732), .B2(new_n410), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n383), .A2(KEYINPUT32), .A3(new_n384), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT70), .B1(new_n387), .B2(new_n388), .ZN(new_n735));
  AOI211_X1 g549(.A(new_n390), .B(new_n364), .C1(new_n356), .C2(new_n359), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n735), .A2(new_n736), .A3(new_n398), .ZN(new_n737));
  INV_X1    g551(.A(new_n407), .ZN(new_n738));
  OAI21_X1  g552(.A(G472), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n733), .A2(new_n734), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n472), .A2(new_n475), .A3(new_n679), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n740), .A2(new_n563), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n731), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G119), .ZN(G21));
  NAND2_X1  g558(.A1(new_n640), .A2(G472), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n381), .B1(new_n367), .B2(new_n369), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n405), .A2(KEYINPUT106), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n388), .B1(new_n405), .B2(KEYINPUT106), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n384), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n702), .A2(new_n666), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n479), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n731), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G122), .ZN(G24));
  NOR3_X1   g569(.A1(new_n751), .A2(new_n714), .A3(new_n681), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n723), .A3(new_n719), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G125), .ZN(G27));
  NAND2_X1  g572(.A1(G469), .A2(G902), .ZN(new_n759));
  XOR2_X1   g573(.A(new_n759), .B(KEYINPUT107), .Z(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n761), .B1(new_n330), .B2(new_n316), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n326), .A2(new_n763), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n655), .A2(new_n556), .A3(new_n690), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n629), .A2(new_n635), .A3(new_n633), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n189), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n764), .A2(new_n480), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT42), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n765), .A2(KEYINPUT42), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n764), .A2(new_n767), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT108), .B1(new_n412), .B2(new_n479), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT108), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n476), .A2(new_n478), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n674), .A2(new_n471), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n740), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT109), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n773), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n762), .B1(new_n320), .B2(new_n325), .ZN(new_n782));
  INV_X1    g596(.A(new_n766), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n188), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n782), .A2(new_n784), .A3(new_n771), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n740), .A2(new_n775), .A3(new_n777), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n775), .B1(new_n740), .B2(new_n777), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT109), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n770), .B1(new_n781), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G131), .ZN(G33));
  NAND4_X1  g605(.A1(new_n764), .A2(new_n480), .A3(new_n691), .A4(new_n767), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G134), .ZN(G36));
  NAND2_X1  g607(.A1(new_n331), .A2(KEYINPUT45), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n316), .B1(new_n330), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n761), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT46), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n797), .A2(KEYINPUT46), .A3(new_n761), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(new_n326), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n188), .A3(new_n706), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT110), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n802), .A2(KEYINPUT110), .A3(new_n188), .A4(new_n706), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n556), .A2(new_n654), .A3(new_n648), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT43), .ZN(new_n808));
  OR3_X1    g622(.A1(new_n655), .A2(KEYINPUT43), .A3(new_n665), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n643), .A2(new_n741), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT44), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n812), .A2(new_n813), .A3(new_n766), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n805), .A2(new_n806), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G137), .ZN(G39));
  NOR4_X1   g630(.A1(new_n740), .A2(new_n714), .A3(new_n777), .A4(new_n766), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n802), .A2(KEYINPUT47), .A3(new_n188), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT47), .B1(new_n802), .B2(new_n188), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n817), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G140), .ZN(G42));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n668), .A2(new_n634), .A3(new_n635), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT111), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT111), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n668), .A2(new_n634), .A3(new_n826), .A4(new_n635), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n634), .A2(new_n712), .A3(new_n635), .A4(new_n666), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n825), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n333), .A3(new_n644), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n830), .A2(new_n637), .A3(new_n683), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n719), .B(new_n723), .C1(new_n753), .C2(new_n742), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n723), .B(new_n480), .C1(new_n660), .C2(new_n669), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n764), .A2(new_n756), .A3(new_n767), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n681), .B1(new_n696), .B2(new_n739), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n515), .A2(new_n556), .A3(new_n713), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n766), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n718), .A2(new_n836), .A3(new_n188), .A4(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n792), .A2(new_n835), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n834), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n790), .A2(new_n831), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n690), .A2(new_n189), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n472), .A2(new_n475), .A3(new_n679), .A4(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n696), .B2(new_n699), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n764), .A2(new_n845), .A3(new_n719), .A4(new_n702), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n694), .A2(new_n720), .A3(new_n846), .A4(new_n757), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT52), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n731), .A2(new_n756), .B1(new_n693), .B2(new_n333), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n849), .A2(new_n850), .A3(new_n720), .A4(new_n846), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n823), .B1(new_n842), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT112), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n850), .B1(new_n694), .B2(new_n757), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n792), .A2(new_n835), .A3(new_n839), .A4(KEYINPUT53), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n790), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n834), .A2(KEYINPUT113), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT113), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n832), .A2(new_n833), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n831), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n852), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n853), .A2(new_n854), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n830), .A2(new_n637), .A3(new_n683), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n867), .A2(new_n834), .A3(new_n840), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n868), .A2(new_n790), .A3(new_n848), .A4(new_n851), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(KEYINPUT112), .A3(new_n823), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n865), .A2(new_n866), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n855), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n869), .B1(new_n823), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n853), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT54), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n809), .A2(new_n808), .A3(new_n688), .ZN(new_n877));
  AND4_X1   g691(.A1(new_n777), .A2(new_n877), .A3(new_n745), .A4(new_n750), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n819), .A2(new_n820), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n326), .B1(new_n316), .B2(new_n324), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n880), .A2(new_n188), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n783), .B(new_n878), .C1(new_n879), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n723), .A2(new_n783), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n700), .A2(new_n777), .A3(new_n558), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n665), .B1(new_n654), .B2(new_n648), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT117), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n886), .A2(new_n890), .A3(new_n887), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n884), .A2(new_n877), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT116), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n741), .A2(new_n745), .A3(new_n750), .ZN(new_n894));
  OR3_X1    g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n893), .B1(new_n892), .B2(new_n894), .ZN(new_n896));
  AOI22_X1  g710(.A1(new_n889), .A2(new_n891), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n882), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n701), .A2(new_n635), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n878), .A2(new_n723), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT50), .B1(new_n900), .B2(KEYINPUT114), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n900), .A2(KEYINPUT114), .A3(KEYINPUT50), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT115), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n904), .B(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT51), .B1(new_n898), .B2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n904), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n882), .A2(new_n897), .A3(KEYINPUT51), .A4(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n892), .A2(new_n779), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT48), .Z(new_n911));
  NAND2_X1  g725(.A1(new_n878), .A2(new_n731), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT118), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n557), .B1(new_n886), .B2(new_n712), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n909), .A2(new_n911), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n876), .A2(new_n907), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(G952), .A2(G953), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n880), .A2(KEYINPUT49), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n880), .A2(KEYINPUT49), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n188), .A2(new_n635), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n701), .A2(new_n807), .A3(new_n920), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n919), .A2(new_n921), .A3(new_n777), .A4(new_n700), .ZN(new_n922));
  OAI22_X1  g736(.A1(new_n916), .A2(new_n917), .B1(new_n918), .B2(new_n922), .ZN(G75));
  NAND2_X1  g737(.A1(new_n853), .A2(new_n854), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n863), .A2(new_n864), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(new_n925), .A3(new_n870), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n926), .A2(G210), .A3(G902), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT56), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n613), .A2(new_n621), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(new_n619), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT55), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n927), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n931), .B1(new_n927), .B2(new_n928), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n279), .A2(G952), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(G51));
  XNOR2_X1  g749(.A(new_n760), .B(KEYINPUT57), .ZN(new_n936));
  AND4_X1   g750(.A1(new_n866), .A2(new_n924), .A3(new_n925), .A4(new_n870), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n866), .B1(new_n865), .B2(new_n870), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n315), .B(KEYINPUT119), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n926), .A2(G902), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n942), .A2(new_n797), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n934), .B1(new_n941), .B2(new_n943), .ZN(G54));
  NOR2_X1   g758(.A1(new_n537), .A2(new_n550), .ZN(new_n945));
  NAND2_X1  g759(.A1(KEYINPUT58), .A2(G475), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n945), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n934), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n942), .A2(new_n945), .A3(new_n946), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(G60));
  NAND2_X1  g765(.A1(new_n651), .A2(new_n653), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n647), .B(KEYINPUT59), .Z(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n876), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n952), .A2(new_n953), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n926), .A2(KEYINPUT54), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n955), .B1(new_n956), .B2(new_n871), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n954), .A2(new_n934), .A3(new_n957), .ZN(G63));
  NAND2_X1  g772(.A1(G217), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT120), .Z(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT60), .Z(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(new_n865), .B2(new_n870), .ZN(new_n963));
  INV_X1    g777(.A(new_n476), .ZN(new_n964));
  OAI21_X1  g778(.A(KEYINPUT121), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n934), .B1(new_n963), .B2(new_n678), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n926), .A2(new_n961), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT121), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n967), .A2(new_n968), .A3(new_n476), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n965), .A2(new_n966), .A3(new_n969), .A4(KEYINPUT61), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n926), .A2(new_n678), .A3(new_n961), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n948), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n963), .A2(new_n964), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n970), .A2(new_n975), .ZN(G66));
  OAI21_X1  g790(.A(G953), .B1(new_n560), .B2(new_n588), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n867), .A2(new_n834), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n977), .B1(new_n978), .B2(G953), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n929), .B1(G898), .B2(new_n279), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(G69));
  OAI21_X1  g795(.A(new_n347), .B1(new_n354), .B2(new_n355), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(new_n548), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n515), .A2(new_n665), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n480), .B(new_n783), .C1(new_n712), .C2(new_n984), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n707), .A2(new_n985), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n815), .A2(new_n821), .A3(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n694), .A2(new_n720), .A3(new_n757), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT122), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n710), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(KEYINPUT62), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT62), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n989), .A2(new_n992), .A3(new_n710), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n987), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n983), .B1(new_n994), .B2(new_n279), .ZN(new_n995));
  INV_X1    g809(.A(new_n983), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n788), .A2(new_n719), .A3(new_n702), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n805), .B(new_n806), .C1(new_n814), .C2(new_n997), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n790), .A2(new_n792), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n998), .A2(new_n999), .A3(new_n821), .A4(new_n989), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n279), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n279), .A2(G900), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT123), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n996), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n995), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n279), .B1(G227), .B2(G900), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT124), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1006), .B1(new_n996), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1005), .B(new_n1008), .ZN(G72));
  NOR2_X1   g823(.A1(new_n387), .A2(new_n364), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n821), .A2(new_n989), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1012), .A2(new_n978), .A3(new_n999), .A4(new_n998), .ZN(new_n1013));
  NAND2_X1  g827(.A1(G472), .A2(G902), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT63), .Z(new_n1015));
  AOI21_X1  g829(.A(new_n1011), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(KEYINPUT126), .B1(new_n1016), .B2(new_n934), .ZN(new_n1017));
  INV_X1    g831(.A(new_n978), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1015), .B1(new_n1000), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n1010), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT126), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1020), .A2(new_n1021), .A3(new_n948), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1017), .A2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n987), .A2(new_n991), .A3(new_n978), .A4(new_n993), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1024), .A2(new_n1015), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT125), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1024), .A2(KEYINPUT125), .A3(new_n1015), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1027), .A2(new_n698), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n356), .A2(new_n365), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n391), .A2(new_n1030), .A3(new_n392), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1031), .A2(new_n1015), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1032), .B(KEYINPUT127), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1033), .B1(new_n873), .B2(new_n874), .ZN(new_n1034));
  AND3_X1   g848(.A1(new_n1023), .A2(new_n1029), .A3(new_n1034), .ZN(G57));
endmodule


