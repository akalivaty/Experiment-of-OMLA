//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966;
  XNOR2_X1  g000(.A(G71gat), .B(G78gat), .ZN(new_n202));
  XOR2_X1   g001(.A(G57gat), .B(G64gat), .Z(new_n203));
  AOI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(KEYINPUT9), .ZN(new_n204));
  AOI21_X1  g003(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT95), .ZN(new_n206));
  AND3_X1   g005(.A1(new_n203), .A2(new_n202), .A3(new_n206), .ZN(new_n207));
  OR2_X1    g006(.A1(new_n205), .A2(KEYINPUT95), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n204), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n209), .A2(KEYINPUT21), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n211));
  XOR2_X1   g010(.A(new_n210), .B(new_n211), .Z(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G15gat), .B(G22gat), .ZN(new_n214));
  INV_X1    g013(.A(G1gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT16), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G1gat), .B2(new_n214), .ZN(new_n218));
  INV_X1    g017(.A(G8gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n209), .A2(KEYINPUT21), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G183gat), .ZN(new_n223));
  INV_X1    g022(.A(G183gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n220), .A2(new_n221), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT96), .ZN(new_n227));
  INV_X1    g026(.A(G231gat), .ZN(new_n228));
  INV_X1    g027(.A(G233gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT96), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n223), .A2(new_n231), .A3(new_n225), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n227), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n230), .B1(new_n227), .B2(new_n232), .ZN(new_n235));
  XNOR2_X1  g034(.A(G127gat), .B(G155gat), .ZN(new_n236));
  INV_X1    g035(.A(G211gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  NOR3_X1   g037(.A1(new_n234), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n238), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n227), .A2(new_n232), .ZN(new_n241));
  INV_X1    g040(.A(new_n230), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n240), .B1(new_n243), .B2(new_n233), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n213), .B1(new_n239), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n238), .B1(new_n234), .B2(new_n235), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n243), .A2(new_n233), .A3(new_n240), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n247), .A3(new_n212), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G134gat), .B(G162gat), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT14), .ZN(new_n252));
  NOR2_X1   g051(.A1(G29gat), .A2(G36gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT89), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT89), .B1(G29gat), .B2(G36gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n255), .B(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT15), .ZN(new_n259));
  XOR2_X1   g058(.A(G43gat), .B(G50gat), .Z(new_n260));
  XOR2_X1   g059(.A(KEYINPUT90), .B(G36gat), .Z(new_n261));
  AOI22_X1  g060(.A1(new_n259), .A2(new_n260), .B1(new_n261), .B2(G29gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n260), .A2(new_n259), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n258), .B(new_n262), .C1(new_n259), .C2(new_n260), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(KEYINPUT91), .A2(KEYINPUT17), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  OR2_X1    g069(.A1(KEYINPUT91), .A2(KEYINPUT17), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n265), .A2(new_n266), .A3(new_n271), .A4(new_n268), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G85gat), .A2(G92gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT98), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT97), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n276), .A2(KEYINPUT7), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n276), .B(KEYINPUT7), .C1(KEYINPUT97), .C2(new_n274), .ZN(new_n278));
  INV_X1    g077(.A(G85gat), .ZN(new_n279));
  INV_X1    g078(.A(G92gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G99gat), .A2(G106gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT8), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n277), .A2(new_n278), .A3(new_n281), .A4(new_n283), .ZN(new_n284));
  XOR2_X1   g083(.A(G99gat), .B(G106gat), .Z(new_n285));
  OR2_X1    g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n285), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AND2_X1   g087(.A1(G232gat), .A2(G233gat), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n273), .A2(new_n288), .B1(KEYINPUT41), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n288), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n267), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n251), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n289), .A2(KEYINPUT41), .ZN(new_n295));
  XNOR2_X1  g094(.A(G190gat), .B(G218gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n290), .A2(new_n251), .A3(new_n292), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n294), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n297), .B1(new_n294), .B2(new_n298), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n249), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT99), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n284), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(new_n209), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT10), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n286), .A2(new_n209), .A3(new_n287), .A4(new_n304), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n291), .A2(KEYINPUT10), .A3(new_n209), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n309), .A2(new_n310), .B1(G230gat), .B2(G233gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G230gat), .A2(G233gat), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n313), .B1(new_n306), .B2(new_n308), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n312), .A2(KEYINPUT100), .A3(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G176gat), .B(G204gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT101), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(G120gat), .ZN(new_n319));
  INV_X1    g118(.A(G148gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n316), .B(new_n321), .C1(KEYINPUT100), .C2(new_n315), .ZN(new_n322));
  INV_X1    g121(.A(new_n321), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT100), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n311), .A2(new_n324), .A3(new_n314), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n315), .A2(KEYINPUT100), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n323), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n302), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(KEYINPUT102), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n331));
  INV_X1    g130(.A(G141gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G148gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n320), .A2(G141gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT2), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G155gat), .B(G162gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n335), .A2(new_n339), .A3(new_n337), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n331), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G211gat), .A2(G218gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT22), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g146(.A1(G197gat), .A2(G204gat), .ZN(new_n348));
  AND2_X1   g147(.A1(G197gat), .A2(G204gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n345), .ZN(new_n351));
  NOR2_X1   g150(.A1(G211gat), .A2(G218gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT78), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  OR2_X1    g153(.A1(G197gat), .A2(G204gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(G197gat), .A2(G204gat), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n355), .A2(new_n356), .B1(new_n346), .B2(new_n345), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT78), .ZN(new_n358));
  XNOR2_X1  g157(.A(G211gat), .B(G218gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n354), .A2(new_n360), .A3(KEYINPUT80), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT80), .B1(new_n354), .B2(new_n360), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n357), .A2(new_n359), .ZN(new_n363));
  NOR3_X1   g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT29), .B1(new_n341), .B2(new_n342), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n344), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT81), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n354), .A2(new_n360), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n350), .A2(KEYINPUT77), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT77), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n347), .B(new_n371), .C1(new_n348), .C2(new_n349), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n353), .A3(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n341), .A2(new_n342), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(KEYINPUT3), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT80), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n369), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n363), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n354), .A2(new_n360), .A3(KEYINPUT80), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n365), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(new_n344), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n378), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G228gat), .A2(G233gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(G22gat), .ZN(new_n390));
  OAI211_X1 g189(.A(KEYINPUT82), .B(new_n344), .C1(new_n374), .C2(new_n366), .ZN(new_n391));
  INV_X1    g190(.A(new_n388), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n369), .A2(new_n373), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n343), .B1(new_n394), .B2(new_n365), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n378), .B1(new_n395), .B2(KEYINPUT82), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT83), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n395), .A2(KEYINPUT82), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n388), .B1(new_n395), .B2(KEYINPUT82), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT83), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n398), .A2(new_n399), .A3(new_n400), .A4(new_n378), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n389), .A2(new_n390), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n390), .B1(new_n389), .B2(new_n402), .ZN(new_n404));
  XNOR2_X1  g203(.A(G78gat), .B(G106gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(KEYINPUT31), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(G50gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(KEYINPUT84), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n403), .A2(new_n404), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n385), .B1(new_n384), .B2(new_n344), .ZN(new_n411));
  AOI211_X1 g210(.A(KEYINPUT81), .B(new_n343), .C1(new_n383), .C2(new_n365), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n392), .B1(new_n413), .B2(new_n378), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n397), .A2(new_n401), .ZN(new_n415));
  OAI211_X1 g214(.A(G22gat), .B(new_n409), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n389), .A2(new_n390), .A3(new_n402), .A4(new_n407), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n410), .A2(new_n418), .ZN(new_n419));
  XOR2_X1   g218(.A(G8gat), .B(G36gat), .Z(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(G64gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(new_n280), .ZN(new_n422));
  INV_X1    g221(.A(G190gat), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT27), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT68), .B1(new_n424), .B2(G183gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT27), .B(G183gat), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n423), .B(new_n425), .C1(new_n426), .C2(KEYINPUT68), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT69), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT28), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT68), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n424), .A2(G183gat), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n224), .A2(KEYINPUT27), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n434), .A2(KEYINPUT69), .A3(new_n423), .A4(new_n425), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n429), .A2(new_n430), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n426), .A2(KEYINPUT28), .A3(new_n423), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT26), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NOR3_X1   g240(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(G169gat), .A2(G176gat), .ZN(new_n444));
  NOR2_X1   g243(.A1(G169gat), .A2(G176gat), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT70), .B1(new_n445), .B2(new_n439), .ZN(new_n446));
  OR3_X1    g245(.A1(new_n445), .A2(KEYINPUT70), .A3(new_n439), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n443), .A2(new_n444), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(G183gat), .A2(G190gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n438), .A2(new_n451), .ZN(new_n452));
  OR3_X1    g251(.A1(KEYINPUT67), .A2(G183gat), .A3(G190gat), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT24), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n453), .A2(new_n455), .A3(new_n456), .A4(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT23), .B1(new_n441), .B2(new_n442), .ZN(new_n459));
  AND4_X1   g258(.A1(KEYINPUT25), .A2(new_n458), .A3(new_n444), .A4(new_n459), .ZN(new_n460));
  OR2_X1    g259(.A1(new_n445), .A2(KEYINPUT23), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OR3_X1    g261(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n463), .A2(new_n455), .A3(new_n456), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n445), .A2(KEYINPUT23), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n465), .A2(new_n444), .A3(new_n466), .A4(new_n461), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT25), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n462), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(G226gat), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(new_n229), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n452), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n450), .B1(new_n436), .B2(new_n437), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n460), .A2(new_n461), .B1(new_n468), .B2(new_n467), .ZN(new_n476));
  OAI22_X1  g275(.A1(new_n475), .A2(new_n476), .B1(KEYINPUT29), .B2(new_n472), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n474), .A2(new_n477), .A3(new_n394), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n394), .B1(new_n474), .B2(new_n477), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n422), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n474), .A2(new_n477), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n374), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n474), .A2(new_n477), .A3(new_n394), .ZN(new_n483));
  INV_X1    g282(.A(new_n422), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n480), .A2(new_n485), .A3(KEYINPUT30), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT30), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n482), .A2(new_n483), .A3(new_n487), .A4(new_n484), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT40), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT39), .ZN(new_n491));
  INV_X1    g290(.A(new_n376), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT72), .ZN(new_n493));
  INV_X1    g292(.A(G113gat), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT71), .ZN(new_n495));
  INV_X1    g294(.A(G120gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n496), .A2(G113gat), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n493), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT1), .ZN(new_n502));
  XOR2_X1   g301(.A(G127gat), .B(G134gat), .Z(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  AND2_X1   g303(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n506));
  OAI21_X1  g305(.A(G113gat), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n500), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(KEYINPUT72), .A3(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n501), .A2(new_n502), .A3(new_n504), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT73), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n507), .A2(new_n508), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n503), .B1(new_n512), .B2(new_n493), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT73), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n513), .A2(new_n514), .A3(new_n502), .A4(new_n509), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  XOR2_X1   g315(.A(G113gat), .B(G120gat), .Z(new_n517));
  AOI21_X1  g316(.A(new_n504), .B1(new_n517), .B2(new_n502), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n492), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  AOI211_X1 g319(.A(new_n518), .B(new_n376), .C1(new_n511), .C2(new_n515), .ZN(new_n521));
  NAND2_X1  g320(.A1(G225gat), .A2(G233gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT4), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n516), .A2(new_n519), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n525), .B1(new_n526), .B2(new_n376), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n518), .B1(new_n511), .B2(new_n515), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n528), .A2(KEYINPUT4), .A3(new_n492), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n492), .A2(new_n331), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n526), .A2(new_n530), .A3(new_n344), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n527), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  AOI211_X1 g331(.A(new_n491), .B(new_n524), .C1(new_n523), .C2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(new_n491), .A3(new_n523), .ZN(new_n534));
  XOR2_X1   g333(.A(G1gat), .B(G29gat), .Z(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G57gat), .B(G85gat), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n537), .B(new_n538), .Z(new_n539));
  NAND2_X1  g338(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n490), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n523), .A2(KEYINPUT5), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n527), .A2(new_n531), .A3(new_n529), .A4(new_n542), .ZN(new_n543));
  OAI22_X1  g342(.A1(new_n526), .A2(new_n376), .B1(new_n525), .B2(new_n523), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n544), .A2(new_n529), .A3(new_n531), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n523), .B1(new_n520), .B2(new_n521), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT5), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n543), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n539), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n523), .ZN(new_n551));
  INV_X1    g350(.A(new_n524), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(new_n552), .A3(KEYINPUT39), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n553), .A2(KEYINPUT40), .A3(new_n539), .A4(new_n534), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n489), .A2(new_n541), .A3(new_n550), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n482), .A2(new_n483), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n484), .B1(new_n556), .B2(KEYINPUT37), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT37), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n482), .A2(new_n558), .A3(new_n483), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT85), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT85), .A4(new_n558), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n557), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT38), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT86), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n563), .A2(KEYINPUT86), .A3(KEYINPUT38), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT6), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n543), .B(new_n539), .C1(new_n545), .C2(new_n547), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n550), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n548), .A2(KEYINPUT6), .A3(new_n549), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT38), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n557), .A2(new_n561), .A3(new_n573), .A4(new_n562), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n571), .A2(new_n572), .A3(new_n485), .A4(new_n574), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n419), .B(new_n555), .C1(new_n568), .C2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n489), .B1(new_n571), .B2(new_n572), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(G22gat), .B1(new_n414), .B2(new_n415), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n389), .A2(new_n390), .A3(new_n402), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n580), .A3(new_n408), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n581), .A2(new_n417), .A3(new_n416), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT76), .ZN(new_n584));
  XNOR2_X1  g383(.A(KEYINPUT75), .B(G15gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G43gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(G71gat), .B(G99gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G227gat), .A2(G233gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT64), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n528), .A2(new_n452), .A3(new_n470), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n528), .B1(new_n452), .B2(new_n470), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n588), .B1(new_n593), .B2(KEYINPUT32), .ZN(new_n594));
  INV_X1    g393(.A(new_n590), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n511), .A2(new_n515), .ZN(new_n596));
  OAI22_X1  g395(.A1(new_n596), .A2(new_n518), .B1(new_n475), .B2(new_n476), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n528), .A2(new_n452), .A3(new_n470), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT74), .B1(new_n599), .B2(KEYINPUT33), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT74), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT33), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n593), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n594), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n593), .B(KEYINPUT32), .C1(new_n602), .C2(new_n588), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n597), .A2(new_n595), .A3(new_n598), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT34), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n604), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n608), .B1(new_n604), .B2(new_n605), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n584), .B(KEYINPUT36), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n584), .B1(new_n609), .B2(new_n610), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT36), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n576), .A2(new_n583), .A3(new_n611), .A4(new_n614), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n582), .A2(new_n609), .A3(new_n610), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT35), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT87), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n617), .A2(KEYINPUT87), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n616), .A2(new_n577), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n621));
  INV_X1    g420(.A(new_n608), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n416), .A2(new_n417), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n604), .A2(new_n605), .A3(new_n608), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n581), .A4(new_n625), .ZN(new_n626));
  OAI211_X1 g425(.A(KEYINPUT87), .B(new_n617), .C1(new_n578), .C2(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n620), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n330), .B1(new_n615), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n273), .A2(new_n220), .ZN(new_n630));
  NAND2_X1  g429(.A1(G229gat), .A2(G233gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n220), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n267), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n630), .A2(KEYINPUT18), .A3(new_n631), .A4(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n220), .A2(new_n265), .A3(new_n266), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n633), .A2(KEYINPUT93), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n631), .B(KEYINPUT13), .Z(new_n637));
  INV_X1    g436(.A(KEYINPUT93), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n267), .A2(new_n632), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n634), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT11), .B(G169gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G197gat), .ZN(new_n643));
  XOR2_X1   g442(.A(G113gat), .B(G141gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT12), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT18), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n641), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT92), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n647), .A2(KEYINPUT92), .A3(new_n648), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n652), .A2(new_n641), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n646), .B(KEYINPUT88), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n654), .A2(KEYINPUT94), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT94), .B1(new_n654), .B2(new_n656), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n650), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n629), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n571), .A2(new_n572), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(new_n215), .ZN(G1324gat));
  INV_X1    g462(.A(new_n660), .ZN(new_n664));
  NAND2_X1  g463(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n665));
  OR2_X1    g464(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n664), .A2(new_n489), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT42), .ZN(new_n668));
  OR3_X1    g467(.A1(new_n667), .A2(KEYINPUT103), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n219), .B1(new_n664), .B2(new_n489), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n670), .B1(new_n668), .B2(new_n667), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT103), .B1(new_n667), .B2(new_n668), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(G1325gat));
  NAND2_X1  g472(.A1(new_n623), .A2(new_n625), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(G15gat), .B1(new_n664), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n614), .A2(new_n611), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n660), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n676), .B1(G15gat), .B2(new_n679), .ZN(G1326gat));
  NOR2_X1   g479(.A1(new_n660), .A2(new_n419), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT43), .B(G22gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT104), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n681), .B(new_n683), .ZN(G1327gat));
  AOI21_X1  g483(.A(new_n301), .B1(new_n628), .B2(new_n615), .ZN(new_n685));
  INV_X1    g484(.A(new_n650), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT94), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n647), .A2(KEYINPUT92), .A3(new_n648), .ZN(new_n688));
  AOI21_X1  g487(.A(KEYINPUT92), .B1(new_n647), .B2(new_n648), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n634), .A2(new_n640), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n687), .B1(new_n691), .B2(new_n655), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n654), .A2(KEYINPUT94), .A3(new_n656), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n686), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n694), .A2(new_n249), .A3(new_n328), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n685), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(G29gat), .ZN(new_n697));
  INV_X1    g496(.A(new_n661), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT45), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT105), .B1(new_n685), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n301), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n419), .A2(new_n555), .ZN(new_n704));
  INV_X1    g503(.A(new_n575), .ZN(new_n705));
  INV_X1    g504(.A(new_n567), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT86), .B1(new_n563), .B2(KEYINPUT38), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n704), .B1(new_n705), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n577), .A2(new_n419), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n709), .A2(new_n677), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n620), .A2(new_n627), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n703), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(new_n714), .A3(KEYINPUT44), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n678), .A2(new_n576), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n710), .B(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n628), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n719), .A2(new_n701), .A3(new_n703), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n702), .A2(new_n715), .A3(new_n720), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n721), .A2(new_n698), .A3(new_n695), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n700), .B1(new_n697), .B2(new_n722), .ZN(G1328gat));
  INV_X1    g522(.A(new_n261), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n696), .A2(new_n724), .A3(new_n489), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT107), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT46), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n721), .A2(new_n489), .A3(new_n695), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n261), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(G1329gat));
  INV_X1    g529(.A(new_n696), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n731), .A2(G43gat), .A3(new_n674), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n721), .A2(new_n677), .A3(new_n695), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n732), .B1(new_n733), .B2(G43gat), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g534(.A1(new_n731), .A2(G50gat), .A3(new_n419), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n582), .A3(new_n695), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(G50gat), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n739), .B1(new_n737), .B2(G50gat), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT48), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n738), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  AOI221_X4 g541(.A(new_n736), .B1(new_n739), .B2(KEYINPUT48), .C1(new_n737), .C2(G50gat), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(G1331gat));
  NOR2_X1   g543(.A1(new_n659), .A2(new_n302), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n719), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n328), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(new_n661), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT109), .B(G57gat), .Z(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1332gat));
  INV_X1    g549(.A(new_n489), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n751), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT110), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n746), .A2(new_n328), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n754), .B(new_n755), .Z(G1333gat));
  OAI21_X1  g555(.A(G71gat), .B1(new_n747), .B2(new_n678), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n747), .A2(G71gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n758), .B2(new_n674), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n759), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g559(.A1(new_n747), .A2(new_n419), .ZN(new_n761));
  XNOR2_X1  g560(.A(KEYINPUT111), .B(G78gat), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1335gat));
  AND2_X1   g562(.A1(new_n245), .A2(new_n248), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n694), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n328), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT112), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n721), .A2(new_n698), .A3(new_n768), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n769), .A2(KEYINPUT113), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(KEYINPUT113), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n770), .A2(G85gat), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n719), .A2(new_n703), .A3(new_n766), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT114), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n773), .A2(new_n774), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n698), .A2(new_n279), .A3(new_n328), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT115), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n777), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n772), .A2(new_n782), .ZN(G1336gat));
  AND2_X1   g582(.A1(new_n322), .A2(new_n327), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n784), .A2(G92gat), .A3(new_n751), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n777), .A2(new_n779), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n721), .A2(new_n489), .A3(new_n768), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G92gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n788), .A2(new_n791), .A3(G92gat), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n791), .B1(new_n788), .B2(G92gat), .ZN(new_n793));
  INV_X1    g592(.A(new_n785), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n775), .B2(new_n778), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n792), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n790), .B1(new_n796), .B2(new_n787), .ZN(G1337gat));
  NOR2_X1   g596(.A1(new_n674), .A2(G99gat), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n777), .A2(new_n328), .A3(new_n779), .A4(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n721), .A2(new_n677), .A3(new_n768), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G99gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(G1338gat));
  NOR3_X1   g601(.A1(new_n419), .A2(new_n784), .A3(G106gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n777), .A2(new_n779), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n721), .A2(new_n582), .A3(new_n768), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(G106gat), .ZN(new_n806));
  XNOR2_X1  g605(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n804), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n803), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(KEYINPUT117), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n775), .B2(new_n778), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(KEYINPUT117), .ZN(new_n812));
  AOI22_X1  g611(.A1(new_n811), .A2(new_n812), .B1(new_n805), .B2(G106gat), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n808), .B1(new_n813), .B2(new_n814), .ZN(G1339gat));
  AOI21_X1  g614(.A(new_n631), .B1(new_n630), .B2(new_n633), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n637), .B1(new_n636), .B2(new_n639), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n645), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n650), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n328), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n323), .B1(new_n311), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n309), .A2(new_n310), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT54), .B1(new_n824), .B2(new_n313), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n823), .B1(new_n311), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n823), .B(KEYINPUT55), .C1(new_n311), .C2(new_n825), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(new_n327), .A3(new_n829), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n301), .B(new_n821), .C1(new_n694), .C2(new_n830), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n828), .A2(new_n327), .A3(new_n829), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n820), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n249), .B1(new_n833), .B2(new_n703), .ZN(new_n834));
  AOI22_X1  g633(.A1(new_n831), .A2(new_n834), .B1(new_n745), .B2(new_n784), .ZN(new_n835));
  NOR4_X1   g634(.A1(new_n835), .A2(new_n661), .A3(new_n489), .A4(new_n626), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n659), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n328), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(G120gat), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n505), .A2(new_n506), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(new_n839), .ZN(G1341gat));
  NAND2_X1  g641(.A1(new_n836), .A2(new_n249), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g643(.A1(new_n836), .A2(new_n703), .ZN(new_n845));
  OR3_X1    g644(.A1(new_n845), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(G134gat), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT56), .B1(new_n845), .B2(G134gat), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(G1343gat));
  OAI21_X1  g648(.A(KEYINPUT57), .B1(new_n835), .B2(new_n419), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n419), .A2(KEYINPUT57), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n830), .A2(new_n819), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n764), .B1(new_n852), .B2(new_n301), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n784), .A2(new_n819), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n854), .B1(new_n659), .B2(new_n832), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n853), .B1(new_n855), .B2(new_n301), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n694), .A2(new_n249), .A3(new_n301), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(new_n328), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n851), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n677), .A2(new_n661), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n489), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n850), .A2(new_n659), .A3(new_n859), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(G141gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n582), .B1(new_n856), .B2(new_n858), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n694), .A2(G141gat), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n862), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT119), .B1(new_n869), .B2(KEYINPUT58), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  AOI211_X1 g671(.A(new_n871), .B(new_n872), .C1(new_n864), .C2(new_n868), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT58), .B1(new_n863), .B2(G141gat), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT120), .B1(new_n865), .B2(new_n861), .ZN(new_n875));
  INV_X1    g674(.A(new_n835), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n876), .A2(new_n877), .A3(new_n582), .A4(new_n860), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n875), .A2(new_n751), .A3(new_n867), .A4(new_n878), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n874), .A2(KEYINPUT121), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT121), .B1(new_n874), .B2(new_n879), .ZN(new_n881));
  OAI22_X1  g680(.A1(new_n870), .A2(new_n873), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n879), .A2(new_n864), .A3(new_n872), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT121), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n874), .A2(KEYINPUT121), .A3(new_n879), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n889), .B(KEYINPUT122), .C1(new_n870), .C2(new_n873), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n884), .A2(new_n890), .ZN(G1344gat));
  AND2_X1   g690(.A1(new_n875), .A2(new_n751), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n878), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n320), .A3(new_n328), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n330), .A2(new_n659), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n851), .B1(new_n897), .B2(new_n856), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n850), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n328), .A3(new_n862), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n896), .B1(new_n901), .B2(G148gat), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n850), .A2(new_n862), .A3(new_n859), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n896), .B1(new_n903), .B2(new_n784), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n904), .A2(new_n320), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n895), .B1(new_n902), .B2(new_n905), .ZN(G1345gat));
  AOI21_X1  g705(.A(G155gat), .B1(new_n894), .B2(new_n249), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n903), .A2(new_n764), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(G155gat), .B2(new_n908), .ZN(G1346gat));
  OAI21_X1  g708(.A(G162gat), .B1(new_n903), .B2(new_n301), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n301), .A2(G162gat), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n910), .B1(new_n893), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT123), .ZN(G1347gat));
  NOR2_X1   g713(.A1(new_n835), .A2(new_n626), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n698), .A2(new_n751), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(G169gat), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n917), .A2(new_n918), .A3(new_n659), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(KEYINPUT124), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n915), .A2(new_n916), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n924), .A2(new_n659), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n919), .B1(new_n925), .B2(new_n918), .ZN(G1348gat));
  AOI21_X1  g725(.A(G176gat), .B1(new_n917), .B2(new_n328), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n924), .A2(new_n328), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(G176gat), .ZN(G1349gat));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n930), .A2(KEYINPUT60), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n920), .A2(new_n249), .A3(new_n923), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(G183gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n917), .A2(new_n249), .A3(new_n426), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n930), .A2(KEYINPUT60), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n935), .B(new_n936), .ZN(G1350gat));
  NAND3_X1  g736(.A1(new_n917), .A2(new_n423), .A3(new_n703), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n703), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(G190gat), .ZN(new_n941));
  AOI211_X1 g740(.A(KEYINPUT61), .B(new_n423), .C1(new_n924), .C2(new_n703), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(G1351gat));
  NOR3_X1   g742(.A1(new_n677), .A2(new_n698), .A3(new_n751), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n866), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(G197gat), .B1(new_n945), .B2(new_n659), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n944), .B(KEYINPUT126), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n899), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n659), .A2(G197gat), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(G1352gat));
  INV_X1    g749(.A(G204gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n945), .A2(new_n951), .A3(new_n328), .ZN(new_n952));
  XOR2_X1   g751(.A(new_n952), .B(KEYINPUT62), .Z(new_n953));
  NAND2_X1  g752(.A1(new_n900), .A2(new_n328), .ZN(new_n954));
  OAI21_X1  g753(.A(G204gat), .B1(new_n954), .B2(new_n947), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n955), .ZN(G1353gat));
  NAND3_X1  g755(.A1(new_n945), .A2(new_n237), .A3(new_n249), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n900), .A2(new_n249), .A3(new_n944), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT63), .B1(new_n958), .B2(G211gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(G1354gat));
  NAND3_X1  g760(.A1(new_n948), .A2(G218gat), .A3(new_n703), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n703), .ZN(new_n963));
  INV_X1    g762(.A(G218gat), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


