//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G104), .ZN(new_n193));
  INV_X1    g007(.A(G101), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n189), .A2(G107), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n190), .A2(new_n193), .A3(new_n194), .A4(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n189), .A2(G107), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n192), .A2(G104), .ZN(new_n198));
  OAI21_X1  g012(.A(G101), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT76), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n196), .A2(new_n199), .A3(KEYINPUT76), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT10), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n205), .B1(G143), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n206), .A2(G143), .ZN(new_n211));
  OAI22_X1  g025(.A1(new_n207), .A2(new_n208), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n213), .B1(new_n209), .B2(G146), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n206), .A2(KEYINPUT64), .A3(G143), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n209), .A2(G146), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n204), .B1(new_n212), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n202), .A2(new_n203), .A3(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n190), .A2(new_n193), .A3(new_n195), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G101), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(KEYINPUT4), .A3(new_n196), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  OR2_X1    g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n224), .B(new_n225), .C1(new_n210), .C2(new_n211), .ZN(new_n226));
  INV_X1    g040(.A(new_n224), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n214), .A2(new_n215), .A3(new_n217), .A4(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n221), .A2(new_n230), .A3(G101), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n223), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n214), .A2(new_n215), .A3(new_n217), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT1), .B1(new_n209), .B2(G146), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT75), .ZN(new_n235));
  OAI21_X1  g049(.A(G128), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n206), .A2(G143), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT75), .B1(new_n237), .B2(KEYINPUT1), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n233), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n200), .B1(new_n239), .B2(new_n218), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n220), .B(new_n232), .C1(KEYINPUT10), .C2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G137), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT65), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G137), .ZN(new_n245));
  AND2_X1   g059(.A1(KEYINPUT11), .A2(G134), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(KEYINPUT11), .A2(G134), .ZN(new_n248));
  NOR2_X1   g062(.A1(KEYINPUT11), .A2(G134), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(G137), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G131), .ZN(new_n252));
  INV_X1    g066(.A(G131), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n247), .A2(new_n253), .A3(new_n250), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n255), .B(KEYINPUT77), .ZN(new_n256));
  OR2_X1    g070(.A1(new_n241), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(G110), .B(G140), .ZN(new_n258));
  INV_X1    g072(.A(G953), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n259), .A2(G227), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n258), .B(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT79), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n241), .A2(new_n263), .A3(new_n255), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n263), .B1(new_n241), .B2(new_n255), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n257), .B(new_n262), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  AND2_X1   g080(.A1(KEYINPUT78), .A2(KEYINPUT12), .ZN(new_n267));
  OR2_X1    g081(.A1(new_n267), .A2(KEYINPUT12), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT78), .B1(new_n252), .B2(new_n254), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n200), .A2(new_n218), .A3(new_n212), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n268), .B(new_n269), .C1(new_n240), .C2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n200), .A2(new_n218), .A3(new_n212), .ZN(new_n273));
  AND4_X1   g087(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n234), .A2(new_n235), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n237), .A2(KEYINPUT75), .A3(KEYINPUT1), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(G128), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n274), .B1(new_n277), .B2(new_n233), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n273), .B1(new_n278), .B2(new_n200), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n268), .B1(new_n279), .B2(new_n269), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n272), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n241), .A2(new_n256), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n261), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n266), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT80), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT80), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n266), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n285), .A2(G469), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G469), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT70), .B(G902), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n241), .A2(new_n255), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT79), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n241), .A2(new_n263), .A3(new_n255), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n262), .B1(new_n294), .B2(new_n257), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n262), .B1(new_n241), .B2(new_n256), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n281), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n289), .B(new_n290), .C1(new_n295), .C2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n289), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n188), .B1(new_n288), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT81), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n290), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n257), .B1(new_n264), .B2(new_n265), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n261), .ZN(new_n308));
  INV_X1    g122(.A(new_n297), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n306), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n300), .B1(new_n310), .B2(new_n289), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n285), .A2(G469), .A3(new_n287), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(KEYINPUT81), .A3(new_n188), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n305), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G140), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G125), .ZN(new_n317));
  INV_X1    g131(.A(G125), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G140), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT16), .ZN(new_n320));
  OR3_X1    g134(.A1(new_n318), .A2(KEYINPUT16), .A3(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n206), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT72), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n320), .A2(new_n321), .A3(G146), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G119), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G128), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n208), .A2(G119), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XOR2_X1   g144(.A(KEYINPUT24), .B(G110), .Z(new_n331));
  INV_X1    g145(.A(KEYINPUT71), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n328), .A2(new_n329), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT24), .B(G110), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT71), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT23), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n337), .B1(new_n327), .B2(G128), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n208), .A2(KEYINPUT23), .A3(G119), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n339), .A3(new_n328), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n333), .A2(new_n336), .B1(G110), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n322), .A2(KEYINPUT72), .A3(new_n206), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n326), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(G125), .B(G140), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n206), .ZN(new_n345));
  INV_X1    g159(.A(G110), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n338), .A2(new_n339), .A3(new_n346), .A4(new_n328), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT73), .ZN(new_n348));
  OAI22_X1  g162(.A1(new_n347), .A2(new_n348), .B1(new_n330), .B2(new_n331), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n347), .A2(new_n348), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n325), .B(new_n345), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n343), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT22), .B(G137), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n259), .A2(G221), .A3(G234), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n353), .B(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n343), .A2(new_n351), .A3(new_n355), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT25), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(KEYINPUT74), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n306), .B1(KEYINPUT74), .B2(new_n360), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n359), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G217), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(new_n290), .B2(G234), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n357), .A2(new_n358), .A3(new_n363), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n367), .B1(new_n368), .B2(new_n361), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n364), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n366), .A2(G902), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n359), .A2(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT69), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n327), .A2(G116), .ZN(new_n376));
  INV_X1    g190(.A(G116), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G119), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G113), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT2), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT2), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G113), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n379), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n383), .ZN(new_n385));
  XNOR2_X1  g199(.A(G116), .B(G119), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n387), .A3(KEYINPUT66), .ZN(new_n388));
  OR3_X1    g202(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT66), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G134), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n243), .A2(new_n245), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n253), .B1(G134), .B2(G137), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n234), .A2(G128), .B1(new_n237), .B2(new_n217), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n254), .B(new_n394), .C1(new_n274), .C2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n226), .A2(new_n228), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n398), .B1(new_n252), .B2(new_n254), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT30), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n247), .A2(new_n253), .A3(new_n250), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n253), .B1(new_n247), .B2(new_n250), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n228), .B(new_n226), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT30), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(new_n404), .A3(new_n396), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n390), .B1(new_n400), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n403), .A2(new_n396), .A3(new_n390), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT26), .B(G101), .ZN(new_n410));
  INV_X1    g224(.A(G237), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n411), .A2(new_n259), .A3(G210), .ZN(new_n412));
  OR2_X1    g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n410), .A2(new_n412), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n414), .B1(new_n413), .B2(new_n415), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n375), .B1(new_n409), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT28), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n388), .A2(new_n389), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n397), .B2(new_n399), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n420), .B1(new_n422), .B2(new_n407), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n407), .A2(new_n420), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT29), .B1(new_n425), .B2(new_n418), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n403), .A2(new_n404), .A3(new_n396), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n404), .B1(new_n403), .B2(new_n396), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n421), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n407), .ZN(new_n430));
  INV_X1    g244(.A(new_n418), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(KEYINPUT69), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n419), .A2(new_n426), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n425), .A2(KEYINPUT29), .A3(new_n418), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n434), .A2(new_n290), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT32), .ZN(new_n437));
  NOR2_X1   g251(.A1(G472), .A2(G902), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT31), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT68), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n407), .A2(new_n418), .A3(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n406), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n407), .A2(new_n418), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT68), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n439), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n407), .A2(new_n418), .A3(new_n440), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n429), .A2(new_n444), .A3(new_n439), .A4(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n431), .B1(new_n423), .B2(new_n424), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n438), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n436), .A2(G472), .B1(new_n437), .B2(new_n450), .ZN(new_n451));
  OAI211_X1 g265(.A(KEYINPUT32), .B(new_n438), .C1(new_n445), .C2(new_n449), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n374), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT89), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n209), .B2(G128), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n208), .A2(KEYINPUT89), .A3(G143), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n209), .A2(G128), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT91), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n455), .A2(new_n456), .B1(G128), .B2(new_n209), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT91), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n391), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n460), .A2(G134), .A3(new_n463), .ZN(new_n466));
  OAI21_X1  g280(.A(KEYINPUT87), .B1(new_n377), .B2(G122), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT87), .ZN(new_n468));
  INV_X1    g282(.A(G122), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n469), .A3(G116), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n377), .A2(G122), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(KEYINPUT14), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n474), .A3(G107), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n471), .B(new_n472), .C1(KEYINPUT14), .C2(new_n192), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n465), .A2(new_n466), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  XOR2_X1   g291(.A(KEYINPUT88), .B(KEYINPUT13), .Z(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n457), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n461), .B1(new_n479), .B2(G134), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT88), .B(KEYINPUT13), .ZN(new_n481));
  AND4_X1   g295(.A1(G134), .A2(new_n457), .A3(new_n458), .A4(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n473), .A2(new_n192), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n471), .A2(G107), .A3(new_n472), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n483), .A2(new_n486), .A3(KEYINPUT90), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT90), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n481), .B1(new_n455), .B2(new_n456), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n459), .B1(new_n489), .B2(new_n391), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n479), .A2(G134), .A3(new_n461), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n484), .A2(new_n485), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n488), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n477), .B1(new_n487), .B2(new_n494), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n187), .A2(new_n365), .A3(G953), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT92), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT90), .B1(new_n483), .B2(new_n486), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n492), .A2(new_n493), .A3(new_n488), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(new_n497), .A3(new_n477), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n499), .A2(new_n290), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT93), .ZN(new_n505));
  INV_X1    g319(.A(G478), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n506), .A2(KEYINPUT15), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT93), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n499), .A2(new_n508), .A3(new_n290), .A4(new_n503), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n505), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n504), .A2(new_n507), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n259), .A2(G952), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(G234), .B2(G237), .ZN(new_n513));
  AOI211_X1 g327(.A(new_n259), .B(new_n290), .C1(G234), .C2(G237), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT21), .B(G898), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n510), .A2(new_n511), .A3(new_n517), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n223), .A2(new_n389), .A3(new_n388), .A4(new_n231), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n386), .A2(KEYINPUT5), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n377), .A2(G119), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT5), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n380), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n520), .A2(new_n523), .B1(new_n386), .B2(new_n385), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n202), .A2(new_n203), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(G110), .B(G122), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n519), .A2(new_n525), .A3(new_n527), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(KEYINPUT6), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT6), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n526), .A2(new_n532), .A3(new_n528), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n212), .A2(new_n218), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(G125), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n318), .B1(new_n226), .B2(new_n228), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n259), .A2(G224), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n531), .A2(new_n533), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n536), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n541), .B(new_n543), .C1(G125), .C2(new_n534), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n542), .B1(new_n535), .B2(new_n536), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n527), .B(KEYINPUT8), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n196), .A2(new_n199), .A3(KEYINPUT83), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n547), .B1(new_n524), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n379), .A2(new_n522), .ZN(new_n550));
  OAI21_X1  g364(.A(G113), .B1(new_n376), .B2(KEYINPUT5), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n387), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT83), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n552), .B1(new_n553), .B2(new_n200), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n549), .B1(new_n554), .B2(new_n548), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n546), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(G902), .B1(new_n556), .B2(new_n530), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n540), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(G210), .B1(G237), .B2(G902), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n540), .A2(new_n557), .A3(new_n559), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(G214), .B1(G237), .B2(G902), .ZN(new_n564));
  XOR2_X1   g378(.A(new_n564), .B(KEYINPUT82), .Z(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(G237), .A2(G953), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n568), .A2(G143), .A3(G214), .ZN(new_n569));
  AOI21_X1  g383(.A(G143), .B1(new_n568), .B2(G214), .ZN(new_n570));
  OAI21_X1  g384(.A(G131), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT17), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n411), .A2(new_n259), .A3(G214), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n209), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n568), .A2(G143), .A3(G214), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n253), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n571), .A2(new_n572), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n575), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(KEYINPUT17), .A3(G131), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n326), .A2(new_n342), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n578), .A2(KEYINPUT18), .A3(G131), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n344), .B(new_n206), .ZN(new_n584));
  NAND2_X1  g398(.A1(KEYINPUT18), .A2(G131), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n574), .A2(new_n575), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(G113), .B(G122), .Z(new_n588));
  XOR2_X1   g402(.A(KEYINPUT84), .B(G104), .Z(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n582), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n592), .B1(new_n580), .B2(new_n581), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(new_n590), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n299), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(KEYINPUT86), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT86), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n597), .B(new_n299), .C1(new_n591), .C2(new_n594), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(G475), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT20), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n571), .A2(new_n576), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT19), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT19), .B1(new_n317), .B2(new_n319), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n206), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n601), .A2(new_n325), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n590), .B1(new_n605), .B2(new_n587), .ZN(new_n606));
  AOI211_X1 g420(.A(KEYINPUT85), .B(new_n606), .C1(new_n593), .C2(new_n590), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT85), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n582), .A2(new_n587), .A3(new_n590), .ZN(new_n609));
  INV_X1    g423(.A(new_n606), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(G475), .A2(G902), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n600), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n609), .A2(new_n610), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(new_n600), .A3(new_n613), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n599), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n518), .A2(new_n567), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n315), .A2(new_n453), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT94), .B(G101), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G3));
  INV_X1    g436(.A(new_n562), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n559), .B1(new_n540), .B2(new_n557), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n564), .B(new_n517), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT95), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n306), .A2(new_n506), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n495), .A2(new_n498), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n497), .B1(new_n502), .B2(new_n477), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT33), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(KEYINPUT33), .B1(new_n499), .B2(new_n503), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n627), .B(new_n628), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n505), .A2(new_n506), .A3(new_n509), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n631), .B1(new_n629), .B2(new_n630), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n499), .A2(KEYINPUT33), .A3(new_n503), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n627), .B1(new_n639), .B2(new_n628), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n626), .B(new_n618), .C1(new_n636), .C2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n290), .B1(new_n445), .B2(new_n449), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(G472), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n450), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n374), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n315), .A2(new_n642), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT34), .B(G104), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  NAND2_X1  g463(.A1(new_n510), .A2(new_n511), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n615), .A2(KEYINPUT85), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n609), .A2(new_n608), .A3(new_n610), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n651), .A2(new_n613), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(KEYINPUT20), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n612), .A2(new_n600), .A3(new_n613), .ZN(new_n655));
  INV_X1    g469(.A(G475), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n656), .B1(new_n595), .B2(KEYINPUT86), .ZN(new_n657));
  AOI22_X1  g471(.A1(new_n654), .A2(new_n655), .B1(new_n598), .B2(new_n657), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n626), .A2(new_n650), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n315), .A2(new_n646), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT35), .B(G107), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  NOR2_X1   g476(.A1(new_n356), .A2(KEYINPUT36), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n352), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n371), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n370), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT96), .ZN(new_n667));
  AOI22_X1  g481(.A1(new_n364), .A2(new_n369), .B1(new_n371), .B2(new_n664), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT96), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n671), .A2(new_n645), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n315), .A2(new_n619), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT97), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT37), .B(G110), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  NAND2_X1  g490(.A1(new_n450), .A2(new_n437), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n434), .A2(new_n290), .ZN(new_n678));
  AOI21_X1  g492(.A(KEYINPUT69), .B1(new_n430), .B2(new_n431), .ZN(new_n679));
  AOI211_X1 g493(.A(new_n375), .B(new_n418), .C1(new_n429), .C2(new_n407), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n678), .B1(new_n681), .B2(new_n426), .ZN(new_n682));
  INV_X1    g496(.A(G472), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n677), .B(new_n452), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n668), .B(KEYINPUT96), .ZN(new_n685));
  INV_X1    g499(.A(new_n564), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n686), .B1(new_n561), .B2(new_n562), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n684), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n513), .ZN(new_n689));
  INV_X1    g503(.A(new_n514), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n689), .B1(new_n690), .B2(G900), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n658), .A2(new_n650), .A3(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n315), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G128), .ZN(G30));
  XNOR2_X1  g509(.A(new_n691), .B(KEYINPUT39), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n315), .A2(new_n696), .ZN(new_n697));
  OR2_X1    g511(.A1(new_n697), .A2(KEYINPUT40), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(KEYINPUT40), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n650), .A2(new_n618), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n700), .A2(new_n686), .A3(new_n666), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n442), .A2(new_n444), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n418), .B1(new_n422), .B2(new_n407), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n299), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G472), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n677), .A3(new_n452), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n563), .B(KEYINPUT38), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n701), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n698), .A2(new_n699), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G143), .ZN(G45));
  AND3_X1   g525(.A1(new_n684), .A2(new_n687), .A3(new_n685), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n618), .B(new_n691), .C1(new_n636), .C2(new_n640), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT81), .B1(new_n313), .B2(new_n188), .ZN(new_n715));
  INV_X1    g529(.A(new_n188), .ZN(new_n716));
  AOI211_X1 g530(.A(new_n304), .B(new_n716), .C1(new_n311), .C2(new_n312), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n712), .B(new_n714), .C1(new_n715), .C2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G146), .ZN(G48));
  AOI21_X1  g533(.A(new_n297), .B1(new_n307), .B2(new_n261), .ZN(new_n720));
  OAI21_X1  g534(.A(G469), .B1(new_n720), .B2(new_n306), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n721), .A2(new_n298), .A3(new_n188), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n684), .A2(new_n722), .A3(new_n373), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n642), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NAND2_X1  g540(.A1(new_n723), .A2(new_n659), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G116), .ZN(G18));
  NAND3_X1  g542(.A1(new_n721), .A2(new_n298), .A3(new_n188), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n729), .A2(new_n518), .A3(new_n618), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n712), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G119), .ZN(G21));
  NAND3_X1  g546(.A1(new_n650), .A2(new_n618), .A3(new_n687), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n721), .A2(new_n298), .A3(new_n188), .A4(new_n517), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n438), .B(KEYINPUT98), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n735), .B1(new_n445), .B2(new_n449), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n644), .A2(new_n373), .A3(new_n736), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n733), .A2(new_n734), .A3(new_n737), .ZN(new_n738));
  XOR2_X1   g552(.A(KEYINPUT99), .B(G122), .Z(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G24));
  NAND3_X1  g554(.A1(new_n644), .A2(new_n666), .A3(new_n736), .ZN(new_n741));
  INV_X1    g555(.A(new_n687), .ZN(new_n742));
  NOR4_X1   g556(.A1(new_n713), .A2(new_n741), .A3(new_n742), .A4(new_n729), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(new_n318), .ZN(G27));
  AOI22_X1  g558(.A1(new_n654), .A2(new_n616), .B1(new_n657), .B2(new_n598), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n634), .A2(new_n635), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n639), .A2(new_n628), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT95), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n745), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n436), .A2(G472), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n445), .A2(new_n449), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT103), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n751), .A2(new_n752), .A3(KEYINPUT32), .A4(new_n438), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n452), .A2(KEYINPUT103), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n750), .A2(new_n753), .A3(new_n677), .A4(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n749), .A2(new_n755), .A3(new_n373), .A4(new_n691), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT100), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n283), .A2(new_n757), .ZN(new_n758));
  OAI211_X1 g572(.A(KEYINPUT100), .B(new_n261), .C1(new_n281), .C2(new_n282), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n758), .A2(G469), .A3(new_n266), .A4(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n298), .A2(new_n301), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT101), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n298), .A2(KEYINPUT101), .A3(new_n301), .A4(new_n760), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT102), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT102), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n561), .A2(new_n768), .A3(new_n562), .A4(new_n564), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n767), .A2(new_n188), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n765), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT42), .B1(new_n756), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n770), .B1(new_n763), .B2(new_n764), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n713), .A2(KEYINPUT42), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n453), .A3(new_n775), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G131), .ZN(G33));
  INV_X1    g592(.A(new_n692), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n774), .A2(new_n453), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G134), .ZN(G36));
  NAND3_X1  g595(.A1(new_n748), .A2(new_n635), .A3(new_n634), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n745), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n783), .A2(KEYINPUT43), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(KEYINPUT43), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n668), .B1(new_n644), .B2(new_n450), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT105), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n767), .A2(new_n769), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n784), .A2(KEYINPUT44), .A3(new_n785), .A4(new_n786), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n789), .A2(new_n790), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT45), .B1(new_n285), .B2(new_n287), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n758), .A2(KEYINPUT45), .A3(new_n266), .A4(new_n759), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(G469), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(new_n300), .ZN(new_n799));
  OAI21_X1  g613(.A(KEYINPUT104), .B1(new_n799), .B2(KEYINPUT46), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT104), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT46), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n801), .B(new_n802), .C1(new_n798), .C2(new_n300), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n799), .A2(KEYINPUT46), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n800), .A2(new_n298), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n805), .A2(new_n188), .A3(new_n696), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n794), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n791), .B1(new_n787), .B2(new_n788), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n790), .B1(new_n809), .B2(new_n793), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G137), .ZN(G39));
  NOR4_X1   g627(.A1(new_n713), .A2(new_n791), .A3(new_n684), .A4(new_n373), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n805), .A2(KEYINPUT47), .A3(new_n188), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT47), .B1(new_n805), .B2(new_n188), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G140), .ZN(G42));
  NAND3_X1  g632(.A1(new_n373), .A2(new_n188), .A3(new_n566), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n819), .B(KEYINPUT106), .Z(new_n820));
  INV_X1    g634(.A(new_n783), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT49), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n721), .A2(new_n298), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n820), .B(new_n821), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT107), .ZN(new_n825));
  AOI211_X1 g639(.A(new_n707), .B(new_n708), .C1(new_n823), .C2(new_n822), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n737), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n784), .A2(new_n513), .A3(new_n828), .A4(new_n785), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT50), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n722), .A2(new_n686), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT110), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n708), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n833), .B1(new_n832), .B2(new_n831), .ZN(new_n834));
  OR3_X1    g648(.A1(new_n829), .A2(new_n830), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n830), .B1(new_n829), .B2(new_n834), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n791), .A2(new_n729), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n784), .A2(new_n513), .A3(new_n785), .A4(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n741), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n707), .A2(new_n374), .A3(new_n689), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n838), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n842), .A2(new_n618), .A3(new_n782), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n837), .A2(KEYINPUT51), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n815), .A2(new_n816), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n823), .A2(new_n716), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n829), .A2(new_n791), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n847), .B1(new_n846), .B2(new_n848), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n845), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n512), .B(KEYINPUT113), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n782), .A2(new_n618), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n854), .B1(new_n842), .B2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n829), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n729), .A2(new_n742), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT48), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n860), .A2(KEYINPUT114), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n755), .A2(new_n373), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n862), .B1(KEYINPUT114), .B2(new_n860), .ZN(new_n863));
  OR3_X1    g677(.A1(new_n839), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n861), .B1(new_n839), .B2(new_n863), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n859), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT115), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT111), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n837), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n835), .A2(KEYINPUT111), .A3(new_n836), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(new_n844), .A3(new_n870), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n791), .B(new_n829), .C1(new_n846), .C2(new_n848), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n853), .B(new_n867), .C1(new_n873), .C2(KEYINPUT51), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT109), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n713), .A2(new_n741), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n774), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n876), .B1(new_n774), .B2(new_n877), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n773), .B(new_n776), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n659), .A2(new_n723), .B1(new_n712), .B2(new_n730), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n738), .B1(new_n642), .B2(new_n723), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n658), .A2(new_n691), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n791), .A2(new_n883), .A3(new_n650), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n671), .B1(new_n451), .B2(new_n452), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n884), .B(new_n885), .C1(new_n715), .C2(new_n717), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n881), .A2(new_n780), .A3(new_n882), .A4(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n563), .A2(new_n566), .A3(new_n517), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n782), .A2(new_n618), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT108), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n889), .A2(new_n891), .A3(new_n745), .A4(new_n650), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n650), .A2(new_n745), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT108), .B1(new_n893), .B2(new_n888), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n890), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(new_n315), .A3(new_n646), .ZN(new_n896));
  OAI221_X1 g710(.A(new_n619), .B1(new_n453), .B2(new_n672), .C1(new_n715), .C2(new_n717), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n880), .A2(new_n887), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n877), .A2(new_n858), .ZN(new_n900));
  INV_X1    g714(.A(new_n733), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n668), .A2(new_n188), .A3(new_n691), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n765), .A2(new_n901), .A3(new_n707), .A4(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n694), .A2(new_n718), .A3(new_n900), .A4(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT52), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n743), .B1(new_n693), .B2(new_n315), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n907), .A2(KEYINPUT52), .A3(new_n718), .A4(new_n903), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n899), .A2(KEYINPUT53), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT53), .B1(new_n899), .B2(new_n909), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n875), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT53), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n906), .A2(new_n908), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n882), .A2(new_n727), .A3(new_n731), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n886), .A2(new_n780), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n896), .A2(new_n897), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n878), .A2(new_n879), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n917), .A2(new_n918), .A3(new_n919), .A4(new_n777), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n913), .B1(new_n914), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n899), .A2(new_n909), .A3(KEYINPUT53), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n921), .A2(KEYINPUT54), .A3(new_n922), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n912), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n874), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(G952), .A2(G953), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n827), .B1(new_n925), .B2(new_n926), .ZN(G75));
  OR2_X1    g741(.A1(new_n259), .A2(G952), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT118), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n290), .B1(new_n921), .B2(new_n922), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n560), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT56), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n531), .A2(new_n533), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n539), .ZN(new_n936));
  XNOR2_X1  g750(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n930), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n932), .A2(KEYINPUT117), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT117), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n931), .A2(new_n941), .A3(new_n560), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n938), .A2(KEYINPUT56), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n939), .A2(new_n944), .ZN(G51));
  XNOR2_X1  g759(.A(new_n300), .B(KEYINPUT57), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n912), .A2(new_n923), .A3(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n720), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(KEYINPUT119), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n931), .A2(new_n798), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n947), .A2(new_n948), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT119), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n930), .B1(new_n951), .B2(new_n954), .ZN(G54));
  NAND2_X1  g769(.A1(KEYINPUT58), .A2(G475), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT120), .Z(new_n957));
  NAND2_X1  g771(.A1(new_n931), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n958), .A2(new_n612), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n612), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n930), .B1(new_n959), .B2(new_n960), .ZN(G60));
  NAND2_X1  g775(.A1(G478), .A2(G902), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT59), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n912), .A2(new_n923), .A3(new_n639), .A4(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT121), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n964), .A2(new_n965), .A3(new_n929), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n639), .B1(new_n924), .B2(new_n963), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n965), .B1(new_n964), .B2(new_n929), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(G63));
  NAND2_X1  g783(.A1(G217), .A2(G902), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT60), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n921), .B2(new_n922), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n664), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n973), .B(new_n929), .C1(new_n359), .C2(new_n972), .ZN(new_n974));
  AOI21_X1  g788(.A(KEYINPUT61), .B1(new_n973), .B2(KEYINPUT122), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(G66));
  INV_X1    g790(.A(G224), .ZN(new_n977));
  OAI21_X1  g791(.A(G953), .B1(new_n515), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n898), .A2(new_n915), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n978), .B1(new_n979), .B2(G953), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n935), .B1(G898), .B2(new_n259), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(G69));
  AND2_X1   g796(.A1(new_n907), .A2(new_n718), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n710), .A2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT62), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n984), .B(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n453), .A2(new_n792), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n855), .A2(new_n893), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n987), .B1(KEYINPUT124), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n989), .B1(KEYINPUT124), .B2(new_n988), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n990), .A2(new_n697), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n991), .B1(new_n808), .B2(new_n811), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n986), .A2(new_n817), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n259), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n400), .A2(new_n405), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n602), .A2(new_n603), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n995), .B(new_n996), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT123), .Z(new_n998));
  NAND2_X1  g812(.A1(new_n994), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n259), .B1(G227), .B2(G900), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n806), .A2(new_n901), .A3(new_n862), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n817), .A2(new_n1002), .A3(new_n777), .A4(new_n780), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n983), .B1(new_n807), .B2(new_n810), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT125), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g820(.A(KEYINPUT125), .B(new_n983), .C1(new_n807), .C2(new_n810), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1003), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n1008), .A2(new_n259), .ZN(new_n1009));
  INV_X1    g823(.A(new_n997), .ZN(new_n1010));
  INV_X1    g824(.A(G900), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1010), .B1(new_n1011), .B2(new_n259), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n999), .B(new_n1001), .C1(new_n1009), .C2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1012), .B1(new_n1008), .B2(new_n259), .ZN(new_n1014));
  INV_X1    g828(.A(new_n998), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(new_n993), .B2(new_n259), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1000), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1013), .A2(new_n1017), .ZN(G72));
  NAND2_X1  g832(.A1(new_n430), .A2(new_n418), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT126), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n984), .B(KEYINPUT62), .ZN(new_n1021));
  INV_X1    g835(.A(new_n979), .ZN(new_n1022));
  INV_X1    g836(.A(new_n991), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n817), .B(new_n1023), .C1(new_n807), .C2(new_n810), .ZN(new_n1024));
  NOR3_X1   g838(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT63), .Z(new_n1027));
  INV_X1    g841(.A(new_n1027), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1020), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  OAI211_X1 g843(.A(KEYINPUT126), .B(new_n1027), .C1(new_n993), .C2(new_n1022), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1019), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n921), .A2(new_n922), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1028), .B1(new_n681), .B2(new_n702), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n930), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1028), .B1(new_n1008), .B2(new_n979), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n430), .A2(new_n418), .ZN(new_n1036));
  XNOR2_X1  g850(.A(new_n1036), .B(KEYINPUT127), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1034), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g852(.A1(new_n1031), .A2(new_n1038), .ZN(G57));
endmodule


