//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n187));
  INV_X1    g001(.A(G137), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(KEYINPUT11), .A3(G134), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G137), .ZN(new_n191));
  AND2_X1   g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G131), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n194), .B1(new_n190), .B2(G137), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT67), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT67), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n197), .B(new_n194), .C1(new_n190), .C2(G137), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n192), .A2(new_n193), .A3(new_n196), .A4(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n189), .A3(new_n191), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n188), .A2(G134), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n197), .B1(new_n201), .B2(new_n194), .ZN(new_n202));
  OAI21_X1  g016(.A(G131), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT65), .B1(new_n204), .B2(G146), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n204), .A2(G146), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT1), .B1(new_n204), .B2(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G128), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(KEYINPUT1), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n205), .A2(new_n208), .A3(new_n209), .A4(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G101), .ZN(new_n218));
  INV_X1    g032(.A(G104), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G107), .ZN(new_n220));
  INV_X1    g034(.A(G107), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n221), .A2(KEYINPUT3), .A3(G104), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT3), .B1(new_n221), .B2(G104), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n218), .B(new_n220), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT80), .B1(new_n221), .B2(G104), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT80), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n219), .A3(G107), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n221), .A2(G104), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G101), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n217), .A2(new_n224), .A3(new_n230), .ZN(new_n231));
  AND4_X1   g045(.A1(new_n205), .A2(new_n208), .A3(new_n209), .A4(new_n215), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n207), .A2(G143), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n211), .A2(G128), .B1(new_n233), .B2(new_n209), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n230), .A2(new_n224), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI221_X4 g051(.A(KEYINPUT12), .B1(new_n199), .B2(new_n203), .C1(new_n231), .C2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT12), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n231), .A2(new_n237), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n203), .A2(new_n199), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n220), .B1(new_n222), .B2(new_n223), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n218), .A2(KEYINPUT4), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(KEYINPUT79), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT79), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n221), .A2(G104), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT3), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n249), .B1(new_n219), .B2(G107), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n221), .A2(KEYINPUT3), .A3(G104), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n245), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n247), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(new_n252), .B2(new_n218), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n244), .A2(G101), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n246), .A2(new_n254), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  OR2_X1    g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n204), .A2(G146), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n207), .A2(G143), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n259), .B(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n259), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n205), .A2(new_n208), .A3(new_n264), .A4(new_n209), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n263), .A2(new_n265), .A3(KEYINPUT70), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT70), .B1(new_n263), .B2(new_n265), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n261), .A2(new_n262), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n214), .B1(new_n233), .B2(KEYINPUT1), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n216), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n271), .A2(KEYINPUT10), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n230), .A2(new_n224), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n258), .A2(new_n268), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n241), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT82), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n276), .B1(new_n231), .B2(new_n278), .ZN(new_n279));
  AOI211_X1 g093(.A(KEYINPUT82), .B(new_n277), .C1(new_n273), .C2(new_n217), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n274), .B(new_n275), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n243), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(G110), .B(G140), .ZN(new_n283));
  INV_X1    g097(.A(G953), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n284), .A2(G227), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n283), .B(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n286), .B(KEYINPUT78), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n282), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT83), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n274), .B1(new_n280), .B2(new_n279), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n241), .ZN(new_n292));
  INV_X1    g106(.A(new_n286), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n281), .A3(new_n293), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n289), .A2(new_n290), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n290), .B1(new_n289), .B2(new_n294), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n295), .A2(new_n296), .A3(G902), .ZN(new_n297));
  INV_X1    g111(.A(G469), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n187), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n281), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n232), .B1(new_n210), .B2(new_n212), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n278), .B1(new_n301), .B2(new_n236), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT82), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n231), .A2(new_n276), .A3(new_n278), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n275), .B1(new_n305), .B2(new_n274), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n300), .A2(new_n306), .A3(new_n286), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n287), .B1(new_n243), .B2(new_n281), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT83), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G902), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n289), .A2(new_n290), .A3(new_n294), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(KEYINPUT84), .A3(G469), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n243), .A2(new_n281), .A3(new_n293), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n286), .B1(new_n300), .B2(new_n306), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT85), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n282), .A2(KEYINPUT85), .A3(new_n286), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n298), .B(new_n310), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n299), .A2(new_n313), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G221), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT9), .B(G234), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n321), .B1(new_n323), .B2(new_n310), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(G214), .B1(G237), .B2(G902), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(KEYINPUT86), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n263), .A2(new_n265), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G125), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n330), .B1(G125), .B2(new_n271), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n284), .A2(G224), .ZN(new_n332));
  XOR2_X1   g146(.A(new_n332), .B(KEYINPUT90), .Z(new_n333));
  XNOR2_X1  g147(.A(new_n331), .B(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT2), .B(G113), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G116), .B(G119), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G119), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G116), .ZN(new_n340));
  INV_X1    g154(.A(G116), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G119), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n342), .A3(KEYINPUT5), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT5), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n339), .A3(G116), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT87), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT87), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n347), .A2(new_n344), .A3(new_n339), .A4(G116), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n343), .A2(new_n346), .A3(G113), .A4(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n273), .A2(new_n338), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT68), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT69), .B1(new_n337), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n340), .A2(new_n342), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT69), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(KEYINPUT68), .A3(new_n354), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n352), .A2(new_n355), .A3(new_n335), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n335), .B1(new_n352), .B2(new_n355), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT79), .B1(new_n244), .B2(new_n245), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n252), .A2(new_n247), .A3(new_n253), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n224), .A2(KEYINPUT4), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n252), .A2(new_n218), .ZN(new_n362));
  OAI22_X1  g176(.A1(new_n359), .A2(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n350), .B1(new_n358), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(G110), .B(G122), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n349), .A2(new_n338), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(new_n236), .ZN(new_n369));
  NOR3_X1   g183(.A1(new_n337), .A2(new_n351), .A3(KEYINPUT69), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n354), .B1(new_n353), .B2(KEYINPUT68), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n336), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n352), .A2(new_n355), .A3(new_n335), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n369), .B1(new_n258), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n365), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n367), .A2(new_n376), .A3(KEYINPUT6), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n258), .A2(new_n374), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n365), .B1(new_n378), .B2(new_n350), .ZN(new_n379));
  XOR2_X1   g193(.A(KEYINPUT88), .B(KEYINPUT6), .Z(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT89), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT89), .ZN(new_n383));
  NOR4_X1   g197(.A1(new_n375), .A2(new_n383), .A3(new_n365), .A4(new_n380), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n334), .B(new_n377), .C1(new_n382), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n332), .A2(KEYINPUT7), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n331), .A2(new_n386), .ZN(new_n387));
  XOR2_X1   g201(.A(new_n365), .B(KEYINPUT8), .Z(new_n388));
  NAND2_X1  g202(.A1(new_n368), .A2(new_n236), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n388), .B1(new_n350), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n331), .A2(new_n386), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n387), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(G902), .B1(new_n392), .B2(new_n376), .ZN(new_n393));
  OAI21_X1  g207(.A(G210), .B1(G237), .B2(G902), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n385), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n394), .B1(new_n385), .B2(new_n393), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n328), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT94), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT91), .ZN(new_n399));
  INV_X1    g213(.A(G125), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(G140), .ZN(new_n401));
  INV_X1    g215(.A(G140), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(G125), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n399), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(G125), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n400), .A2(G140), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT91), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(KEYINPUT19), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(G125), .B(G140), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT19), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT92), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n410), .A2(KEYINPUT92), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n409), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n408), .A2(new_n207), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G237), .ZN(new_n415));
  AND4_X1   g229(.A1(G143), .A2(new_n415), .A3(new_n284), .A4(G214), .ZN(new_n416));
  NOR2_X1   g230(.A1(G237), .A2(G953), .ZN(new_n417));
  AOI21_X1  g231(.A(G143), .B1(new_n417), .B2(G214), .ZN(new_n418));
  OAI21_X1  g232(.A(G131), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n415), .A2(new_n284), .A3(G214), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n204), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n417), .A2(G143), .A3(G214), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n193), .A3(new_n422), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n400), .A2(KEYINPUT16), .A3(G140), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n424), .B1(new_n409), .B2(KEYINPUT16), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n419), .A2(new_n423), .B1(new_n425), .B2(G146), .ZN(new_n426));
  NAND2_X1  g240(.A1(KEYINPUT18), .A2(G131), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n421), .A2(new_n422), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n427), .B1(new_n421), .B2(new_n422), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n404), .A2(G146), .A3(new_n407), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n409), .A2(new_n207), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n414), .A2(new_n426), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  XOR2_X1   g248(.A(G113), .B(G122), .Z(new_n435));
  XOR2_X1   g249(.A(KEYINPUT93), .B(G104), .Z(new_n436));
  XOR2_X1   g250(.A(new_n435), .B(new_n436), .Z(new_n437));
  OAI21_X1  g251(.A(new_n398), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n426), .A2(new_n414), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n430), .A2(new_n433), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n437), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n441), .A2(KEYINPUT94), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n425), .A2(G146), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT16), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT16), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n401), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n207), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT95), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n444), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n445), .A2(G146), .A3(new_n447), .ZN(new_n452));
  AOI21_X1  g266(.A(G146), .B1(new_n445), .B2(new_n447), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT95), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT17), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n419), .A2(new_n456), .A3(new_n423), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n456), .B2(new_n419), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n437), .B(new_n440), .C1(new_n455), .C2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n438), .A2(new_n443), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT96), .ZN(new_n461));
  NOR2_X1   g275(.A1(G475), .A2(G902), .ZN(new_n462));
  XOR2_X1   g276(.A(new_n462), .B(KEYINPUT97), .Z(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT96), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n438), .A2(new_n443), .A3(new_n465), .A4(new_n459), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n461), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT20), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n463), .A2(KEYINPUT20), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n460), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n455), .A2(new_n458), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n437), .B1(new_n472), .B2(new_n440), .ZN(new_n473));
  INV_X1    g287(.A(new_n459), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n310), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n341), .A2(G122), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n341), .A2(G122), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n478), .B1(new_n479), .B2(KEYINPUT14), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT14), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n341), .A3(G122), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(KEYINPUT101), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT101), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n484), .B(new_n478), .C1(new_n479), .C2(KEYINPUT14), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(G107), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT102), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT102), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n483), .A2(new_n488), .A3(G107), .A4(new_n485), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n204), .A2(G128), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n214), .A2(G143), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n190), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT100), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n491), .A2(new_n492), .A3(new_n190), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n496), .ZN(new_n498));
  OAI21_X1  g312(.A(KEYINPUT100), .B1(new_n498), .B2(new_n493), .ZN(new_n499));
  INV_X1    g313(.A(new_n479), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(new_n478), .A3(new_n221), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n490), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n204), .A2(KEYINPUT13), .A3(G128), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n204), .A2(G128), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n505), .B1(new_n506), .B2(KEYINPUT99), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(KEYINPUT99), .B2(new_n505), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT13), .B1(new_n204), .B2(G128), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT98), .ZN(new_n510));
  OAI21_X1  g324(.A(G134), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n500), .A2(new_n478), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G107), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n498), .B1(new_n513), .B2(new_n501), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G217), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n322), .A2(new_n516), .A3(G953), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n504), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n517), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n502), .B1(new_n487), .B2(new_n489), .ZN(new_n520));
  INV_X1    g334(.A(new_n515), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(G902), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(G478), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n523), .B1(KEYINPUT15), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n517), .B1(new_n504), .B2(new_n515), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n520), .A2(new_n521), .A3(new_n519), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n310), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n524), .A2(KEYINPUT15), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI211_X1 g344(.A(new_n310), .B(new_n284), .C1(G234), .C2(G237), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT21), .B(G898), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n284), .A2(G952), .ZN(new_n534));
  INV_X1    g348(.A(G234), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n534), .B1(new_n535), .B2(new_n415), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n525), .A2(new_n530), .A3(new_n537), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n397), .A2(new_n477), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n320), .A2(new_n325), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT74), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT66), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n203), .A2(new_n199), .B1(new_n329), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n263), .A2(new_n265), .A3(KEYINPUT66), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n201), .A2(new_n191), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G131), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n271), .A2(new_n199), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n358), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT28), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n199), .A2(new_n547), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n268), .A2(new_n241), .B1(new_n552), .B2(new_n271), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n551), .B1(new_n553), .B2(new_n358), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT70), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n329), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n263), .A2(new_n265), .A3(KEYINPUT70), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n241), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n558), .A2(new_n358), .A3(new_n551), .A4(new_n548), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n550), .B1(new_n554), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT73), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n417), .A2(G210), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT27), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT26), .B(G101), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n561), .A2(new_n562), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n558), .A2(new_n358), .A3(new_n548), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT28), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n549), .B1(new_n570), .B2(new_n559), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT73), .B1(new_n571), .B2(new_n566), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n558), .A2(KEYINPUT30), .A3(new_n548), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n543), .A2(new_n544), .B1(new_n552), .B2(new_n271), .ZN(new_n575));
  XOR2_X1   g389(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n576));
  OAI211_X1 g390(.A(new_n574), .B(new_n374), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(new_n569), .A3(new_n566), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT31), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT71), .ZN(new_n580));
  XOR2_X1   g394(.A(KEYINPUT72), .B(KEYINPUT31), .Z(new_n581));
  OR2_X1    g395(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT71), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n578), .A2(new_n583), .A3(KEYINPUT31), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n573), .A2(new_n580), .A3(new_n582), .A4(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(G472), .A2(G902), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT32), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT29), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n571), .A2(new_n567), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n566), .B1(new_n553), .B2(new_n358), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n577), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n591), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n553), .A2(new_n358), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n570), .B2(new_n559), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n567), .A2(new_n591), .ZN(new_n598));
  AOI21_X1  g412(.A(G902), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G472), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n590), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT32), .B1(new_n585), .B2(new_n586), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n541), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n585), .A2(new_n586), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n588), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n585), .A2(new_n589), .B1(new_n600), .B2(G472), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n607), .A3(KEYINPUT74), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n516), .B1(G234), .B2(new_n310), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT22), .B(G137), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n321), .A2(new_n535), .A3(G953), .ZN(new_n611));
  XOR2_X1   g425(.A(new_n610), .B(new_n611), .Z(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(G119), .B(G128), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT24), .B(G110), .Z(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(KEYINPUT75), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT24), .B(G110), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT75), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n614), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n339), .A2(G128), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT76), .B1(new_n214), .B2(G119), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT23), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI211_X1 g438(.A(KEYINPUT76), .B(KEYINPUT23), .C1(new_n214), .C2(G119), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n624), .A2(G110), .A3(new_n625), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n444), .B(new_n432), .C1(new_n620), .C2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n616), .A2(new_n614), .A3(new_n619), .ZN(new_n628));
  OAI21_X1  g442(.A(G110), .B1(new_n624), .B2(new_n625), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n628), .B(new_n629), .C1(new_n453), .C2(new_n452), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(KEYINPUT77), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT77), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n627), .B2(new_n630), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n613), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n631), .A2(new_n612), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(KEYINPUT25), .B1(new_n637), .B2(new_n310), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT25), .ZN(new_n639));
  AOI211_X1 g453(.A(new_n639), .B(G902), .C1(new_n635), .C2(new_n636), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n609), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n609), .A2(G902), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n604), .A2(new_n608), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n540), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT103), .B(G101), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G3));
  AND2_X1   g462(.A1(new_n313), .A2(new_n319), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n324), .B1(new_n649), .B2(new_n299), .ZN(new_n650));
  INV_X1    g464(.A(G472), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n585), .B2(new_n310), .ZN(new_n652));
  INV_X1    g466(.A(new_n579), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n653), .A2(new_n583), .B1(new_n568), .B2(new_n572), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n578), .A2(new_n581), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(KEYINPUT71), .B2(new_n579), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n587), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n641), .A2(new_n643), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n652), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(KEYINPUT33), .B1(new_n526), .B2(new_n527), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT33), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n518), .A2(new_n522), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n660), .A2(G478), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n524), .A2(new_n310), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n664), .B1(new_n523), .B2(new_n524), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  AOI22_X1  g481(.A1(new_n467), .A2(KEYINPUT20), .B1(new_n460), .B2(new_n469), .ZN(new_n668));
  INV_X1    g482(.A(new_n476), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n667), .B(new_n537), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n397), .A2(KEYINPUT104), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n672), .B(new_n328), .C1(new_n395), .C2(new_n396), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n670), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n650), .A2(new_n659), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(KEYINPUT105), .Z(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT34), .B(G104), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G6));
  NAND2_X1  g492(.A1(new_n468), .A2(KEYINPUT106), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n467), .A2(new_n680), .A3(KEYINPUT20), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n461), .A2(new_n466), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n469), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n679), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n525), .A2(new_n530), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n476), .A3(new_n537), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n671), .B2(new_n673), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n650), .A2(new_n659), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT35), .B(G107), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G9));
  XNOR2_X1  g506(.A(new_n631), .B(KEYINPUT77), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n693), .B1(KEYINPUT36), .B2(new_n613), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n632), .A2(new_n634), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n613), .A2(KEYINPUT36), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI211_X1 g511(.A(G902), .B(new_n609), .C1(new_n694), .C2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n636), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n693), .B2(new_n613), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n639), .B1(new_n700), .B2(G902), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n637), .A2(KEYINPUT25), .A3(new_n310), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n698), .B1(new_n703), .B2(new_n609), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n652), .A2(new_n704), .A3(new_n657), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n320), .A2(new_n705), .A3(new_n325), .A4(new_n539), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT37), .B(G110), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G12));
  NOR3_X1   g522(.A1(new_n602), .A2(new_n541), .A3(new_n603), .ZN(new_n709));
  AOI21_X1  g523(.A(KEYINPUT74), .B1(new_n606), .B2(new_n607), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n694), .A2(new_n697), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n642), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n641), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n385), .A2(new_n393), .ZN(new_n715));
  INV_X1    g529(.A(new_n394), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n385), .A2(new_n393), .A3(new_n394), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n672), .B1(new_n719), .B2(new_n328), .ZN(new_n720));
  INV_X1    g534(.A(new_n673), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n714), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n685), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n669), .ZN(new_n724));
  INV_X1    g538(.A(new_n536), .ZN(new_n725));
  INV_X1    g539(.A(G900), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n725), .B1(new_n531), .B2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n684), .A2(new_n724), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n722), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n711), .A2(new_n730), .A3(new_n650), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G128), .ZN(G30));
  XOR2_X1   g546(.A(new_n727), .B(KEYINPUT39), .Z(new_n733));
  NAND2_X1  g547(.A1(new_n650), .A2(new_n733), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n734), .A2(KEYINPUT40), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(KEYINPUT40), .ZN(new_n736));
  INV_X1    g550(.A(new_n593), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n310), .B1(new_n737), .B2(new_n596), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n567), .B1(new_n577), .B2(new_n569), .ZN(new_n739));
  OAI21_X1  g553(.A(G472), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n606), .A2(new_n590), .A3(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n719), .B(KEYINPUT38), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n477), .A2(new_n685), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n704), .A2(new_n328), .ZN(new_n746));
  NOR4_X1   g560(.A1(new_n742), .A2(new_n744), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n735), .A2(new_n736), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G143), .ZN(G45));
  OAI211_X1 g563(.A(new_n667), .B(new_n728), .C1(new_n668), .C2(new_n669), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n722), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n711), .A2(new_n751), .A3(new_n650), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G146), .ZN(G48));
  OAI21_X1  g567(.A(new_n310), .B1(new_n317), .B2(new_n318), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(G469), .ZN(new_n755));
  AND4_X1   g569(.A1(new_n644), .A2(new_n755), .A3(new_n325), .A4(new_n319), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(new_n604), .A3(new_n674), .A4(new_n608), .ZN(new_n757));
  XNOR2_X1  g571(.A(KEYINPUT41), .B(G113), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G15));
  NAND4_X1  g573(.A1(new_n689), .A2(new_n756), .A3(new_n604), .A4(new_n608), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G116), .ZN(G18));
  NOR3_X1   g575(.A1(new_n668), .A2(new_n538), .A3(new_n669), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n755), .A2(new_n762), .A3(new_n325), .A4(new_n319), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n722), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n711), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n763), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n704), .B1(new_n671), .B2(new_n673), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n767), .A2(new_n604), .A3(new_n768), .A4(new_n608), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT107), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G119), .ZN(G21));
  AOI21_X1  g586(.A(new_n745), .B1(new_n671), .B2(new_n673), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n755), .A2(new_n325), .A3(new_n319), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n597), .A2(new_n566), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n653), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n587), .B1(new_n776), .B2(new_n582), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n652), .A2(new_n777), .A3(new_n658), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n773), .A2(new_n537), .A3(new_n774), .A4(new_n778), .ZN(new_n779));
  XOR2_X1   g593(.A(KEYINPUT108), .B(G122), .Z(new_n780));
  XNOR2_X1  g594(.A(new_n779), .B(new_n780), .ZN(G24));
  NAND2_X1  g595(.A1(new_n671), .A2(new_n673), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n652), .A2(new_n704), .A3(new_n777), .ZN(new_n783));
  INV_X1    g597(.A(new_n750), .ZN(new_n784));
  AND4_X1   g598(.A1(new_n782), .A2(new_n774), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(new_n400), .ZN(G27));
  INV_X1    g600(.A(new_n645), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n298), .A2(new_n310), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n294), .A2(KEYINPUT109), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT109), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n292), .A2(new_n790), .A3(new_n281), .A4(new_n293), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n308), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n788), .B1(new_n792), .B2(G469), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n324), .B1(new_n793), .B2(new_n319), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n717), .A2(new_n328), .A3(new_n718), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n794), .A2(new_n784), .A3(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(KEYINPUT42), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n658), .B1(new_n606), .B2(new_n607), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n799), .A2(new_n784), .A3(new_n796), .A4(new_n794), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n787), .A2(new_n798), .B1(new_n800), .B2(KEYINPUT42), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G131), .ZN(G33));
  INV_X1    g616(.A(new_n729), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(new_n796), .A3(new_n794), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n645), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(new_n190), .ZN(G36));
  NOR2_X1   g620(.A1(new_n477), .A2(new_n666), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT110), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n807), .B1(new_n808), .B2(KEYINPUT43), .ZN(new_n809));
  XOR2_X1   g623(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n810));
  OAI21_X1  g624(.A(new_n810), .B1(new_n477), .B2(new_n666), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n812), .B(new_n714), .C1(new_n657), .C2(new_n652), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT44), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT111), .ZN(new_n816));
  OR3_X1    g630(.A1(new_n295), .A2(new_n296), .A3(KEYINPUT45), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n298), .B1(new_n792), .B2(KEYINPUT45), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n788), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n819), .A2(KEYINPUT46), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n319), .B1(new_n819), .B2(KEYINPUT46), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n325), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n733), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n796), .B1(new_n813), .B2(new_n814), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n816), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G137), .ZN(G39));
  INV_X1    g642(.A(KEYINPUT47), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n822), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n822), .A2(new_n829), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n711), .A2(new_n644), .A3(new_n750), .A4(new_n795), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(G140), .ZN(G42));
  NAND2_X1  g649(.A1(new_n755), .A2(new_n319), .ZN(new_n836));
  XOR2_X1   g650(.A(new_n836), .B(KEYINPUT49), .Z(new_n837));
  AND4_X1   g651(.A1(new_n644), .A2(new_n807), .A3(new_n325), .A4(new_n328), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n742), .A3(new_n744), .A4(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n760), .A2(new_n757), .A3(new_n779), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n771), .A2(new_n840), .A3(KEYINPUT112), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT112), .B1(new_n771), .B2(new_n840), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n719), .A2(new_n328), .A3(new_n537), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n845), .B1(new_n477), .B2(new_n723), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n668), .A2(new_n669), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(KEYINPUT113), .A3(new_n685), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n844), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n320), .A3(new_n325), .A4(new_n659), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n706), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT114), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n670), .A2(new_n397), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n320), .A2(new_n325), .A3(new_n659), .A4(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n854), .B1(new_n540), .B2(new_n645), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n850), .A2(new_n857), .A3(new_n706), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n852), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n783), .ZN(new_n860));
  OAI22_X1  g674(.A1(new_n645), .A2(new_n804), .B1(new_n860), .B2(new_n797), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n604), .A2(new_n608), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n313), .A2(new_n319), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT84), .B1(new_n312), .B2(G469), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n325), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n723), .A2(new_n476), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n704), .A2(new_n795), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(new_n684), .A3(new_n728), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n863), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n801), .A2(new_n862), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n859), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT116), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n714), .A2(new_n727), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n794), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n874), .B1(new_n794), .B2(new_n875), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n741), .B(new_n773), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n755), .A2(new_n325), .A3(new_n319), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n879), .B1(new_n671), .B2(new_n673), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n784), .A3(new_n783), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n731), .A2(new_n752), .A3(new_n878), .A4(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT52), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n863), .A2(new_n866), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n785), .B1(new_n885), .B2(new_n730), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n886), .A2(KEYINPUT52), .A3(new_n752), .A4(new_n878), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n843), .A2(KEYINPUT53), .A3(new_n873), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT117), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n857), .B1(new_n850), .B2(new_n706), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n855), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n861), .A2(new_n870), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n892), .A2(new_n801), .A3(new_n893), .A4(new_n858), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n894), .A2(new_n841), .A3(new_n842), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT53), .A4(new_n888), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n890), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n884), .A2(new_n887), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n771), .A2(new_n840), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT112), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n858), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n903), .A2(new_n891), .A3(new_n855), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n800), .A2(KEYINPUT42), .ZN(new_n905));
  INV_X1    g719(.A(new_n798), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n905), .B1(new_n906), .B2(new_n645), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n907), .A2(new_n870), .A3(new_n861), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n771), .A2(new_n840), .A3(KEYINPUT112), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n902), .A2(new_n904), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n899), .B1(new_n910), .B2(KEYINPUT115), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT115), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n843), .A2(new_n912), .A3(new_n873), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT53), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT54), .B1(new_n898), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT53), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(new_n910), .B2(new_n899), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT118), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n916), .B1(new_n900), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n771), .A2(new_n840), .A3(KEYINPUT118), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n873), .A2(new_n888), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(KEYINPUT54), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n536), .B1(new_n809), .B2(new_n811), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n879), .A2(new_n795), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n927), .A2(new_n799), .ZN(new_n928));
  OR2_X1    g742(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n929));
  NAND2_X1  g743(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n928), .B2(new_n929), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n926), .A2(new_n742), .A3(new_n644), .A4(new_n725), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n847), .A2(new_n666), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n925), .A2(new_n778), .ZN(new_n936));
  INV_X1    g750(.A(new_n880), .ZN(new_n937));
  OAI221_X1 g751(.A(new_n534), .B1(new_n933), .B2(new_n935), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n932), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n936), .A2(new_n795), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n836), .A2(new_n325), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n940), .B1(new_n832), .B2(new_n941), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n743), .A2(new_n879), .A3(new_n328), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n925), .A2(new_n943), .A3(new_n778), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT50), .Z(new_n945));
  NOR3_X1   g759(.A1(new_n933), .A2(new_n477), .A3(new_n667), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n783), .B2(new_n927), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n942), .A2(KEYINPUT51), .A3(new_n945), .A4(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n939), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT119), .ZN(new_n950));
  OAI22_X1  g764(.A1(new_n832), .A2(new_n950), .B1(new_n325), .B2(new_n836), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT119), .B1(new_n830), .B2(new_n831), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n940), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n953), .A2(new_n945), .A3(new_n947), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT51), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n949), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n915), .A2(new_n924), .A3(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(G952), .A2(G953), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n839), .B1(new_n957), .B2(new_n958), .ZN(G75));
  NOR2_X1   g773(.A1(new_n284), .A2(G952), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n310), .B1(new_n917), .B2(new_n921), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT56), .B1(new_n962), .B2(G210), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n377), .B1(new_n382), .B2(new_n384), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(new_n334), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT55), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n961), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g781(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n962), .A2(G210), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n969), .B1(new_n970), .B2(KEYINPUT121), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n922), .A2(G902), .ZN(new_n972));
  INV_X1    g786(.A(G210), .ZN(new_n973));
  OR3_X1    g787(.A1(new_n972), .A2(KEYINPUT121), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n967), .B1(new_n971), .B2(new_n974), .ZN(G51));
  INV_X1    g789(.A(KEYINPUT54), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n917), .B2(new_n921), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n923), .A2(new_n977), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n788), .B(KEYINPUT57), .Z(new_n979));
  OAI22_X1  g793(.A1(new_n978), .A2(new_n979), .B1(new_n317), .B2(new_n318), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n962), .A2(new_n817), .A3(new_n818), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n960), .B1(new_n980), .B2(new_n981), .ZN(G54));
  NAND2_X1  g796(.A1(KEYINPUT58), .A2(G475), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT123), .Z(new_n984));
  NAND3_X1  g798(.A1(new_n922), .A2(G902), .A3(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n682), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n962), .A2(new_n682), .A3(new_n984), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n987), .A2(new_n961), .A3(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT124), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n987), .A2(KEYINPUT124), .A3(new_n961), .A4(new_n988), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(G60));
  NAND2_X1  g807(.A1(new_n660), .A2(new_n662), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n664), .B(KEYINPUT59), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n997), .B1(new_n923), .B2(new_n977), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n961), .ZN(new_n999));
  INV_X1    g813(.A(new_n996), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n890), .A2(new_n897), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n910), .A2(KEYINPUT115), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n1002), .A2(new_n913), .A3(new_n888), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n916), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n976), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1000), .B1(new_n1005), .B2(new_n923), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n999), .B1(new_n1006), .B2(new_n995), .ZN(G63));
  XNOR2_X1  g821(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n516), .A2(new_n310), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n922), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n700), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n922), .A2(new_n712), .A3(new_n1010), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1012), .A2(new_n961), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT61), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1012), .A2(KEYINPUT61), .A3(new_n961), .A4(new_n1013), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(G66));
  NAND2_X1  g832(.A1(new_n843), .A2(new_n904), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n284), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT126), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(G224), .ZN(new_n1023));
  OAI21_X1  g837(.A(G953), .B1(new_n532), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  OR2_X1    g839(.A1(new_n284), .A2(G898), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n964), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1025), .B(new_n1027), .ZN(G69));
  INV_X1    g842(.A(KEYINPUT127), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n408), .A2(new_n413), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1030), .B(new_n1031), .Z(new_n1032));
  AOI21_X1  g846(.A(new_n1032), .B1(G900), .B2(G953), .ZN(new_n1033));
  AOI22_X1  g847(.A1(new_n816), .A2(new_n826), .B1(new_n832), .B2(new_n833), .ZN(new_n1034));
  INV_X1    g848(.A(new_n824), .ZN(new_n1035));
  AND2_X1   g849(.A1(new_n773), .A2(new_n799), .ZN(new_n1036));
  AOI211_X1 g850(.A(new_n907), .B(new_n805), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g851(.A1(new_n1034), .A2(new_n752), .A3(new_n886), .A4(new_n1037), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1033), .B1(new_n1038), .B2(G953), .ZN(new_n1039));
  INV_X1    g853(.A(new_n748), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n886), .A2(new_n752), .ZN(new_n1041));
  OR3_X1    g855(.A1(new_n1040), .A2(KEYINPUT62), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g856(.A(KEYINPUT62), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1043));
  AND2_X1   g857(.A1(new_n846), .A2(new_n848), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n795), .B1(new_n1044), .B2(new_n935), .ZN(new_n1045));
  NAND4_X1  g859(.A1(new_n787), .A2(new_n1045), .A3(new_n650), .A4(new_n733), .ZN(new_n1046));
  NAND4_X1  g860(.A1(new_n1042), .A2(new_n1034), .A3(new_n1043), .A4(new_n1046), .ZN(new_n1047));
  AND2_X1   g861(.A1(new_n1047), .A2(new_n284), .ZN(new_n1048));
  INV_X1    g862(.A(new_n1032), .ZN(new_n1049));
  OAI211_X1 g863(.A(new_n1029), .B(new_n1039), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n284), .B1(G227), .B2(G900), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AND2_X1   g866(.A1(new_n1039), .A2(new_n1029), .ZN(new_n1053));
  INV_X1    g867(.A(new_n1051), .ZN(new_n1054));
  OAI211_X1 g868(.A(new_n1053), .B(new_n1054), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1052), .A2(new_n1055), .ZN(G72));
  NAND2_X1  g870(.A1(G472), .A2(G902), .ZN(new_n1057));
  XOR2_X1   g871(.A(new_n1057), .B(KEYINPUT63), .Z(new_n1058));
  OAI21_X1  g872(.A(new_n1058), .B1(new_n1038), .B2(new_n1019), .ZN(new_n1059));
  AOI21_X1  g873(.A(new_n960), .B1(new_n1059), .B2(new_n594), .ZN(new_n1060));
  OAI21_X1  g874(.A(new_n1058), .B1(new_n1047), .B2(new_n1019), .ZN(new_n1061));
  NAND2_X1  g875(.A1(new_n1061), .A2(new_n739), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g877(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1064));
  INV_X1    g878(.A(new_n1058), .ZN(new_n1065));
  NOR3_X1   g879(.A1(new_n594), .A2(new_n739), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g880(.A(new_n1063), .B1(new_n1064), .B2(new_n1066), .ZN(G57));
endmodule


