//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 0 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1264, new_n1265, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  OAI21_X1  g0007(.A(G50), .B1(G58), .B2(G68), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT64), .Z(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G107), .A2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(G87), .B2(G250), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT66), .B(G244), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n222), .B(new_n223), .C1(new_n202), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT65), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n214), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n213), .B(new_n217), .C1(new_n228), .C2(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT67), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G68), .Z(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  XNOR2_X1  g0046(.A(KEYINPUT69), .B(G1), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(G13), .A3(G20), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT25), .ZN(new_n249));
  NOR3_X1   g0049(.A1(new_n248), .A2(new_n249), .A3(G107), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n249), .B1(new_n248), .B2(G107), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n210), .B1(new_n214), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n247), .A2(G33), .ZN(new_n256));
  AND3_X1   g0056(.A1(new_n248), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n251), .A2(new_n252), .B1(G107), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT70), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n261), .A2(G33), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(new_n266), .A3(KEYINPUT70), .ZN(new_n267));
  INV_X1    g0067(.A(G87), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n268), .A2(KEYINPUT22), .A3(G20), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n264), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n265), .A2(new_n266), .A3(new_n211), .A4(G87), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT22), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT86), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n270), .A2(KEYINPUT86), .A3(new_n272), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n211), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT23), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n280), .B1(new_n211), .B2(G107), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n205), .A2(KEYINPUT23), .A3(G20), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n279), .A2(G116), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(KEYINPUT87), .B1(new_n277), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT24), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n255), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AND3_X1   g0086(.A1(new_n270), .A2(KEYINPUT86), .A3(new_n272), .ZN(new_n287));
  AOI21_X1  g0087(.A(KEYINPUT86), .B1(new_n270), .B2(new_n272), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n283), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT87), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(KEYINPUT87), .B(new_n283), .C1(new_n287), .C2(new_n288), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(KEYINPUT24), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n259), .B1(new_n286), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G41), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(G1), .A3(G13), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n265), .A2(new_n266), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT71), .B(G1698), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G250), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G257), .A2(G1698), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G294), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n253), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n297), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT5), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G41), .ZN(new_n307));
  INV_X1    g0107(.A(G41), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT5), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n247), .A2(G45), .A3(new_n307), .A4(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G274), .ZN(new_n311));
  AND2_X1   g0111(.A1(G1), .A2(G13), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n311), .B1(new_n312), .B2(new_n295), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n310), .A2(G264), .A3(new_n296), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n305), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(G179), .B2(new_n318), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT88), .B1(new_n294), .B2(new_n321), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n291), .A2(KEYINPUT24), .A3(new_n292), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n254), .B1(new_n291), .B2(KEYINPUT24), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n258), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT88), .ZN(new_n326));
  INV_X1    g0126(.A(new_n321), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G190), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n318), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(G200), .B2(new_n318), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n258), .B(new_n331), .C1(new_n323), .C2(new_n324), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n322), .A2(new_n328), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G45), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n308), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n247), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(G238), .A3(new_n296), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT68), .ZN(new_n338));
  AOI21_X1  g0138(.A(G1), .B1(new_n308), .B2(new_n334), .ZN(new_n339));
  AND4_X1   g0139(.A1(new_n338), .A2(new_n339), .A3(new_n296), .A4(G274), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n338), .B1(new_n313), .B2(new_n339), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n337), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n264), .A2(G232), .A3(G1698), .A4(new_n267), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n264), .A2(G226), .A3(new_n267), .A4(new_n299), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G33), .A2(G97), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI211_X1 g0146(.A(KEYINPUT13), .B(new_n342), .C1(new_n297), .C2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT13), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n297), .ZN(new_n349));
  INV_X1    g0149(.A(new_n342), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(G169), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT14), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n349), .A2(new_n350), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT13), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n349), .A2(new_n348), .A3(new_n350), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(G179), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT14), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(G169), .C1(new_n347), .C2(new_n351), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n353), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n278), .A2(new_n202), .B1(new_n211), .B2(G68), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n211), .A2(new_n253), .ZN(new_n362));
  INV_X1    g0162(.A(G50), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n254), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT11), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n247), .A2(G13), .A3(G20), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n367), .A2(new_n254), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n247), .A2(G20), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(G68), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n248), .A2(G68), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n372), .B(KEYINPUT12), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n360), .A2(new_n375), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n265), .A2(new_n266), .A3(KEYINPUT70), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT70), .B1(new_n265), .B2(new_n266), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n379), .A2(G222), .A3(new_n299), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(G1698), .ZN(new_n381));
  INV_X1    g0181(.A(G223), .ZN(new_n382));
  OAI221_X1 g0182(.A(new_n380), .B1(new_n202), .B2(new_n379), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n297), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n313), .A2(new_n339), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT68), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n313), .A2(new_n338), .A3(new_n339), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n297), .B1(new_n247), .B2(new_n335), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G226), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n384), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n393), .A2(KEYINPUT74), .A3(G200), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT74), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n391), .B1(new_n383), .B2(new_n297), .ZN(new_n396));
  INV_X1    g0196(.A(G200), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n396), .A2(G190), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT10), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n368), .A2(G50), .A3(new_n369), .ZN(new_n402));
  NOR2_X1   g0202(.A1(G20), .A2(G33), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G150), .ZN(new_n404));
  XNOR2_X1  g0204(.A(KEYINPUT8), .B(G58), .ZN(new_n405));
  OAI221_X1 g0205(.A(new_n404), .B1(new_n201), .B2(new_n211), .C1(new_n405), .C2(new_n278), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n406), .A2(new_n254), .B1(new_n367), .B2(new_n363), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT9), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n402), .A2(KEYINPUT9), .A3(new_n407), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n400), .A2(new_n401), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT75), .B1(new_n399), .B2(new_n412), .ZN(new_n413));
  AOI211_X1 g0213(.A(new_n329), .B(new_n391), .C1(new_n383), .C2(new_n297), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n410), .A2(new_n411), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n414), .A2(KEYINPUT10), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT75), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n416), .A2(new_n417), .A3(new_n394), .A4(new_n398), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n414), .A2(new_n415), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n397), .B2(new_n396), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT10), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G58), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(new_n219), .ZN(new_n425));
  NOR2_X1   g0225(.A1(G58), .A2(G68), .ZN(new_n426));
  OAI21_X1  g0226(.A(G20), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(G159), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n362), .A2(KEYINPUT76), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT76), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n430), .B1(new_n403), .B2(G159), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n427), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT7), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT3), .B(G33), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n433), .B1(new_n434), .B2(G20), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n298), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n432), .B1(new_n437), .B2(G68), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n255), .B1(new_n438), .B2(KEYINPUT16), .ZN(new_n439));
  AOI21_X1  g0239(.A(G20), .B1(new_n264), .B2(new_n267), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n436), .B1(new_n440), .B2(KEYINPUT7), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n432), .B1(new_n441), .B2(G68), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n439), .B1(new_n442), .B2(KEYINPUT16), .ZN(new_n443));
  INV_X1    g0243(.A(new_n405), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n369), .A2(new_n444), .ZN(new_n445));
  AOI211_X1 g0245(.A(new_n254), .B(new_n367), .C1(KEYINPUT77), .C2(new_n445), .ZN(new_n446));
  OR2_X1    g0246(.A1(new_n445), .A2(KEYINPUT77), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n446), .A2(new_n447), .B1(new_n367), .B2(new_n405), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n443), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(G1698), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT71), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT71), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G1698), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(new_n453), .A3(G223), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G226), .A2(G1698), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n298), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n253), .A2(new_n268), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n297), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n389), .A2(G232), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n388), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G169), .ZN(new_n461));
  INV_X1    g0261(.A(G179), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n461), .B1(new_n462), .B2(new_n460), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n449), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT18), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT18), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n449), .A2(new_n466), .A3(new_n463), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT78), .B1(new_n460), .B2(G190), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n460), .A2(new_n397), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n386), .A2(new_n387), .B1(new_n389), .B2(G232), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT78), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n471), .A2(new_n472), .A3(new_n329), .A4(new_n458), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n469), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(new_n443), .A3(new_n448), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT17), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n474), .A2(KEYINPUT17), .A3(new_n443), .A4(new_n448), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n468), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n355), .A2(G190), .A3(new_n356), .ZN(new_n481));
  OAI21_X1  g0281(.A(G200), .B1(new_n347), .B2(new_n351), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(new_n482), .A3(new_n374), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n393), .A2(G179), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n408), .B1(new_n396), .B2(G169), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT15), .B(G87), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n488), .A2(KEYINPUT72), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(KEYINPUT72), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n279), .ZN(new_n492));
  OAI22_X1  g0292(.A1(new_n405), .A2(new_n362), .B1(new_n211), .B2(new_n202), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n255), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n248), .A2(new_n369), .A3(G77), .A4(new_n255), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n248), .A2(KEYINPUT73), .A3(G77), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT73), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n367), .B2(new_n202), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n496), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OR2_X1    g0300(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n224), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n389), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n388), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n379), .A2(G232), .A3(new_n299), .ZN(new_n505));
  OAI221_X1 g0305(.A(new_n505), .B1(new_n205), .B2(new_n379), .C1(new_n381), .C2(new_n220), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n504), .B1(new_n506), .B2(new_n297), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n501), .B1(new_n507), .B2(G169), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n462), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OR2_X1    g0311(.A1(new_n507), .A2(new_n397), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n501), .B1(new_n507), .B2(G190), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AND4_X1   g0314(.A1(new_n483), .A2(new_n487), .A3(new_n511), .A4(new_n514), .ZN(new_n515));
  AND4_X1   g0315(.A1(new_n376), .A2(new_n423), .A3(new_n480), .A4(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(G257), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n310), .A2(new_n296), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n316), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n379), .A2(KEYINPUT79), .A3(G250), .A4(G1698), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n264), .A2(G250), .A3(G1698), .A4(new_n267), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT79), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g0323(.A1(KEYINPUT4), .A2(G244), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n264), .A2(new_n267), .A3(new_n299), .A4(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n434), .A2(new_n299), .A3(G244), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT4), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n526), .A2(new_n527), .B1(G33), .B2(G283), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n520), .A2(new_n523), .A3(new_n525), .A4(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n519), .B1(new_n529), .B2(new_n297), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G190), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n257), .A2(G97), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n367), .A2(new_n204), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT6), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n535), .A2(new_n204), .A3(G107), .ZN(new_n536));
  XNOR2_X1  g0336(.A(G97), .B(G107), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n536), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  OAI22_X1  g0338(.A1(new_n538), .A2(new_n211), .B1(new_n202), .B2(new_n362), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n436), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n211), .B1(new_n377), .B2(new_n378), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n541), .B1(new_n542), .B2(new_n433), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n540), .B1(new_n543), .B2(new_n205), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n534), .B1(new_n544), .B2(new_n254), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT80), .ZN(new_n546));
  OAI21_X1  g0346(.A(G200), .B1(new_n530), .B2(new_n546), .ZN(new_n547));
  AOI211_X1 g0347(.A(KEYINPUT80), .B(new_n519), .C1(new_n529), .C2(new_n297), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n531), .B(new_n545), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n529), .A2(new_n297), .ZN(new_n550));
  INV_X1    g0350(.A(new_n519), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n550), .A2(new_n462), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n539), .B1(new_n441), .B2(G107), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n533), .B(new_n532), .C1(new_n553), .C2(new_n255), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n552), .B(new_n554), .C1(G169), .C2(new_n530), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n451), .A2(new_n453), .A3(G238), .ZN(new_n556));
  NAND2_X1  g0356(.A1(G244), .A2(G1698), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n298), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(G116), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n253), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n297), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n313), .A2(G45), .A3(new_n247), .ZN(new_n562));
  INV_X1    g0362(.A(G1), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT69), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT69), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G1), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n566), .A3(G45), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT81), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n247), .A2(KEYINPUT81), .A3(G45), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(G250), .A4(new_n296), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n561), .A2(new_n562), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n462), .ZN(new_n574));
  XNOR2_X1  g0374(.A(new_n488), .B(KEYINPUT72), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT19), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n211), .B1(new_n345), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(G87), .B2(new_n206), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n265), .A2(new_n266), .A3(new_n211), .A4(G68), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n576), .B1(new_n278), .B2(new_n204), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n367), .A2(new_n575), .B1(new_n581), .B2(new_n254), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n257), .A2(new_n491), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n319), .A2(new_n572), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n581), .A2(new_n254), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n367), .B1(new_n489), .B2(new_n490), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n248), .A2(new_n256), .A3(G87), .A4(new_n255), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(G200), .B2(new_n572), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n573), .A2(G190), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n574), .A2(new_n584), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n549), .A2(new_n555), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT82), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n549), .A2(KEYINPUT82), .A3(new_n555), .A4(new_n591), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n307), .A2(new_n309), .ZN(new_n597));
  OAI211_X1 g0397(.A(G270), .B(new_n296), .C1(new_n567), .C2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT83), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT83), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n310), .A2(new_n600), .A3(G270), .A4(new_n296), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(G303), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n603), .B1(new_n264), .B2(new_n267), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n451), .A2(new_n453), .A3(G257), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G264), .A2(G1698), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n298), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n297), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n602), .A2(new_n608), .A3(new_n316), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(G200), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n248), .A2(new_n256), .A3(G116), .A4(new_n255), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n367), .A2(new_n559), .ZN(new_n612));
  NAND2_X1  g0412(.A1(G33), .A2(G283), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n613), .B(new_n211), .C1(G33), .C2(new_n204), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n559), .A2(G20), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(new_n254), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT20), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n611), .B(new_n612), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n610), .B(new_n621), .C1(new_n329), .C2(new_n609), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n622), .B(KEYINPUT85), .ZN(new_n623));
  OAI21_X1  g0423(.A(G303), .B1(new_n377), .B2(new_n378), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n605), .A2(new_n606), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n434), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n315), .B1(new_n627), .B2(new_n297), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n319), .B1(new_n628), .B2(new_n602), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n629), .A2(KEYINPUT84), .A3(KEYINPUT21), .A4(new_n620), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n609), .A2(KEYINPUT21), .A3(G169), .A4(new_n620), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT84), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n609), .A2(G169), .A3(new_n620), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT21), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n602), .A2(new_n608), .A3(G179), .A4(new_n316), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n635), .A2(new_n636), .B1(new_n638), .B2(new_n620), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n623), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n333), .A2(new_n516), .A3(new_n596), .A4(new_n642), .ZN(G372));
  INV_X1    g0443(.A(KEYINPUT90), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n286), .A2(new_n293), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n321), .B1(new_n645), .B2(new_n258), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n631), .A2(new_n632), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n631), .A2(new_n632), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n639), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT89), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT89), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n634), .A2(new_n651), .A3(new_n639), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n646), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n332), .A2(new_n549), .A3(new_n555), .A4(new_n591), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n644), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n325), .A2(new_n327), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n634), .A2(new_n651), .A3(new_n639), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n651), .B1(new_n634), .B2(new_n639), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AND4_X1   g0459(.A1(new_n332), .A2(new_n549), .A3(new_n555), .A4(new_n591), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(new_n660), .A3(KEYINPUT90), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n584), .A2(new_n574), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n589), .A2(new_n590), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n662), .B1(new_n555), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT91), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n550), .A2(new_n551), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n545), .B1(new_n668), .B2(new_n319), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n669), .A2(new_n591), .A3(KEYINPUT26), .A4(new_n552), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n666), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  OAI211_X1 g0471(.A(KEYINPUT91), .B(new_n662), .C1(new_n555), .C2(new_n665), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n671), .A2(new_n663), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n655), .A2(new_n661), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n516), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n508), .B1(new_n462), .B2(new_n507), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n483), .A2(new_n676), .B1(new_n360), .B2(new_n375), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n465), .B(new_n467), .C1(new_n677), .C2(new_n479), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n486), .B1(new_n678), .B2(new_n423), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n675), .A2(new_n679), .ZN(G369));
  INV_X1    g0480(.A(new_n333), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n211), .A2(G13), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n247), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n683), .A2(KEYINPUT27), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(KEYINPUT27), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(G213), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(G343), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n325), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT92), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n681), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n688), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n656), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n692), .A2(new_n621), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n650), .A2(new_n652), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n641), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n649), .A2(new_n692), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AOI22_X1  g0502(.A1(new_n691), .A2(new_n702), .B1(new_n646), .B2(new_n692), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n700), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n215), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(G1), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n208), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n674), .A2(new_n692), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n322), .A2(new_n328), .A3(new_n640), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT93), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(new_n716), .A3(new_n660), .ZN(new_n717));
  AOI22_X1  g0517(.A1(new_n666), .A2(new_n670), .B1(new_n574), .B2(new_n584), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n716), .B1(new_n715), .B2(new_n660), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT29), .B(new_n692), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n714), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n641), .A2(new_n688), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n596), .A2(new_n333), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n305), .A2(new_n317), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n572), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n530), .A2(new_n638), .A3(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n530), .A2(new_n638), .A3(KEYINPUT30), .A4(new_n726), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n573), .A2(G179), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n668), .A2(new_n318), .A3(new_n609), .A4(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n688), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT31), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n733), .A2(KEYINPUT31), .A3(new_n688), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n724), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G330), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n722), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT94), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n740), .A2(new_n741), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n711), .B1(new_n746), .B2(G1), .ZN(G364));
  AOI21_X1  g0547(.A(new_n563), .B1(new_n682), .B2(G45), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n706), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n705), .A2(new_n434), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n245), .A2(new_n334), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n753), .B(new_n754), .C1(new_n334), .C2(new_n209), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n379), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n705), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n758), .A2(G355), .B1(new_n559), .B2(new_n705), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n210), .B1(G20), .B2(new_n319), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n751), .B1(new_n760), .B2(new_n765), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n766), .A2(KEYINPUT95), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(KEYINPUT95), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n211), .A2(new_n329), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(G179), .A3(new_n397), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n397), .A2(G179), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n770), .A2(new_n424), .B1(new_n772), .B2(new_n268), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n211), .A2(G190), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n771), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n773), .B1(G107), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G179), .A2(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n428), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT32), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n774), .A2(G179), .A3(new_n397), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n782), .A2(KEYINPUT96), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(KEYINPUT96), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n777), .B(new_n781), .C1(new_n202), .C2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n329), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(G190), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G50), .A2(new_n788), .B1(new_n789), .B2(G68), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n211), .B1(new_n778), .B2(G190), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G97), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n379), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n786), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n770), .ZN(new_n796));
  INV_X1    g0596(.A(new_n779), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n796), .A2(G322), .B1(new_n797), .B2(G329), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n799), .B2(new_n775), .ZN(new_n800));
  INV_X1    g0600(.A(G317), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n801), .A2(KEYINPUT33), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(KEYINPUT33), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n789), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n788), .A2(G326), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n804), .B(new_n805), .C1(new_n303), .C2(new_n791), .ZN(new_n806));
  INV_X1    g0606(.A(G311), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n807), .A2(new_n782), .B1(new_n772), .B2(new_n603), .ZN(new_n808));
  NOR4_X1   g0608(.A1(new_n800), .A2(new_n379), .A3(new_n806), .A4(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n764), .B1(new_n795), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n767), .A2(new_n768), .A3(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT97), .ZN(new_n812));
  INV_X1    g0612(.A(new_n763), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n812), .B1(new_n697), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n750), .B1(new_n697), .B2(G330), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(G330), .B2(new_n697), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G396));
  INV_X1    g0618(.A(KEYINPUT101), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n501), .A2(new_n688), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n514), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n511), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n509), .A2(new_n510), .A3(new_n692), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n819), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n512), .A2(new_n513), .B1(new_n501), .B2(new_n688), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n819), .B(new_n823), .C1(new_n825), .C2(new_n676), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n712), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n674), .A2(new_n692), .A3(new_n828), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n750), .B1(new_n832), .B2(new_n739), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n739), .B2(new_n832), .ZN(new_n834));
  INV_X1    g0634(.A(new_n764), .ZN(new_n835));
  INV_X1    g0635(.A(new_n789), .ZN(new_n836));
  INV_X1    g0636(.A(G150), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(G137), .ZN(new_n839));
  INV_X1    g0639(.A(new_n788), .ZN(new_n840));
  INV_X1    g0640(.A(G143), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n839), .A2(new_n840), .B1(new_n770), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n785), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n838), .B(new_n842), .C1(new_n843), .C2(G159), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT34), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n434), .B1(new_n772), .B2(new_n363), .ZN(new_n846));
  INV_X1    g0646(.A(G132), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n775), .A2(new_n219), .B1(new_n779), .B2(new_n847), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n846), .B(new_n848), .C1(G58), .C2(new_n792), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n844), .A2(KEYINPUT34), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n757), .B1(new_n205), .B2(new_n772), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT99), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n776), .A2(G87), .B1(new_n797), .B2(G311), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n854), .B1(new_n303), .B2(new_n770), .C1(new_n785), .C2(new_n559), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n793), .B1(new_n840), .B2(new_n603), .C1(new_n799), .C2(new_n836), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n850), .A2(new_n851), .B1(new_n853), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n835), .B1(new_n858), .B2(KEYINPUT100), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(KEYINPUT100), .B2(new_n858), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n764), .A2(new_n761), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n750), .B1(G77), .B2(new_n862), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT98), .Z(new_n864));
  OAI211_X1 g0664(.A(new_n860), .B(new_n864), .C1(new_n828), .C2(new_n762), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n834), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(G384));
  INV_X1    g0667(.A(new_n538), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n868), .A2(KEYINPUT35), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(KEYINPUT35), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n869), .A2(G116), .A3(new_n212), .A4(new_n870), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n871), .B(KEYINPUT36), .Z(new_n872));
  OAI21_X1  g0672(.A(G77), .B1(new_n424), .B2(new_n219), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n873), .A2(new_n208), .B1(G50), .B2(new_n219), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n247), .A2(G13), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n872), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(G330), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n596), .A2(new_n333), .A3(new_n723), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n737), .A2(KEYINPUT108), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n736), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n734), .A2(KEYINPUT108), .A3(new_n735), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT109), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT109), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n724), .A2(new_n884), .A3(new_n880), .A4(new_n881), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n516), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT110), .Z(new_n888));
  XNOR2_X1  g0688(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n464), .A2(new_n475), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT37), .ZN(new_n892));
  INV_X1    g0692(.A(new_n686), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n449), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n891), .A2(KEYINPUT107), .A3(new_n892), .A4(new_n894), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n464), .A2(new_n894), .A3(new_n475), .A4(new_n892), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT107), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n464), .A2(new_n894), .A3(new_n475), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT37), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n895), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n449), .B(new_n893), .C1(new_n468), .C2(new_n479), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n890), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n439), .B1(KEYINPUT16), .B2(new_n438), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n686), .B1(new_n904), .B2(new_n448), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n468), .B2(new_n479), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n448), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n463), .B2(new_n893), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n908), .A2(new_n475), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n896), .B1(new_n909), .B2(new_n892), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n906), .A2(KEYINPUT38), .A3(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n903), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT105), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n483), .A2(new_n353), .A3(new_n357), .A4(new_n359), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT104), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n374), .A2(new_n692), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n916), .B1(new_n915), .B2(new_n917), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n359), .A2(new_n357), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n355), .A2(new_n356), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n358), .B1(new_n922), .B2(G169), .ZN(new_n923));
  OAI211_X1 g0723(.A(KEYINPUT103), .B(new_n375), .C1(new_n921), .C2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT103), .B1(new_n360), .B2(new_n375), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n483), .B1(new_n374), .B2(new_n692), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n914), .B1(new_n920), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n915), .A2(new_n917), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT104), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n926), .ZN(new_n934));
  INV_X1    g0734(.A(new_n927), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(new_n924), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n933), .A2(new_n936), .A3(KEYINPUT105), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n829), .B1(new_n929), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n886), .A2(new_n913), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT40), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT38), .B1(new_n906), .B2(new_n910), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n912), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n942), .A2(KEYINPUT40), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n886), .A2(new_n938), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n877), .B1(new_n888), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n888), .B2(new_n945), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n823), .B(KEYINPUT102), .Z(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  AOI221_X4 g0749(.A(new_n942), .B1(new_n929), .B2(new_n937), .C1(new_n831), .C2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT39), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n903), .B2(new_n912), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n688), .B1(new_n934), .B2(new_n924), .ZN(new_n953));
  INV_X1    g0753(.A(new_n941), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(KEYINPUT39), .A3(new_n911), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n468), .A2(new_n686), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n950), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n714), .A2(new_n516), .A3(new_n721), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n960), .A2(new_n679), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n959), .B(new_n961), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n947), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT111), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n964), .B1(new_n247), .B2(new_n682), .C1(new_n962), .C2(new_n947), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n963), .A2(KEYINPUT111), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n876), .B1(new_n965), .B2(new_n966), .ZN(G367));
  OR2_X1    g0767(.A1(new_n234), .A2(new_n753), .ZN(new_n968));
  INV_X1    g0768(.A(new_n765), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n491), .B2(new_n705), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n751), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n688), .A2(new_n588), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n591), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n663), .B2(new_n972), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n775), .A2(new_n202), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n770), .A2(new_n837), .B1(new_n779), .B2(new_n839), .ZN(new_n976));
  INV_X1    g0776(.A(new_n772), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n975), .B(new_n976), .C1(G58), .C2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n843), .A2(G50), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n757), .B1(G143), .B2(new_n788), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n791), .A2(new_n219), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n789), .B2(G159), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n978), .A2(new_n979), .A3(new_n980), .A4(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n772), .A2(new_n559), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n984), .A2(KEYINPUT46), .B1(G294), .B2(new_n789), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(KEYINPUT46), .B2(new_n984), .C1(new_n807), .C2(new_n840), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n775), .A2(new_n204), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G303), .B2(new_n796), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n988), .B(new_n298), .C1(new_n801), .C2(new_n779), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n843), .A2(G283), .B1(G107), .B2(new_n792), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n990), .B1(new_n992), .B2(KEYINPUT113), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT113), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n983), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT47), .Z(new_n997));
  OAI221_X1 g0797(.A(new_n971), .B1(new_n813), .B2(new_n974), .C1(new_n997), .C2(new_n835), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT114), .Z(new_n999));
  OAI211_X1 g0799(.A(new_n549), .B(new_n555), .C1(new_n545), .C2(new_n692), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n555), .B2(new_n692), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n703), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1002), .A2(KEYINPUT44), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT44), .ZN(new_n1004));
  NOR3_X1   g0804(.A1(new_n703), .A2(new_n1004), .A3(new_n1001), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n703), .A2(new_n1001), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT45), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(KEYINPUT45), .B1(new_n703), .B2(new_n1001), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n1003), .A2(new_n1005), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(new_n699), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n691), .A2(new_n702), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n694), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1012), .B1(new_n1013), .B2(new_n702), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(new_n698), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n746), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n706), .B(KEYINPUT41), .Z(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n749), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1001), .B(KEYINPUT112), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n322), .A2(new_n328), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n688), .B1(new_n1024), .B2(new_n555), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n691), .A2(new_n702), .A3(new_n1001), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT42), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1020), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n700), .A2(new_n1022), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1030), .B(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n999), .B1(new_n1019), .B2(new_n1033), .ZN(G387));
  INV_X1    g0834(.A(new_n1015), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n746), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT116), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1036), .A2(new_n1037), .A3(new_n706), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n745), .A2(new_n1015), .ZN(new_n1039));
  OAI21_X1  g0839(.A(KEYINPUT116), .B1(new_n1039), .B2(new_n707), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1038), .B(new_n1040), .C1(new_n746), .C2(new_n1035), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n752), .B1(new_n238), .B2(new_n334), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n758), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1042), .B1(new_n708), .B2(new_n1043), .ZN(new_n1044));
  OR3_X1    g0844(.A1(new_n405), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1045));
  OAI21_X1  g0845(.A(KEYINPUT50), .B1(new_n405), .B2(G50), .ZN(new_n1046));
  AOI21_X1  g0846(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1045), .A2(new_n708), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1044), .A2(new_n1048), .B1(new_n205), .B2(new_n705), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n750), .B1(new_n1049), .B2(new_n969), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n575), .A2(new_n791), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n770), .A2(new_n363), .B1(new_n772), .B2(new_n202), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n782), .A2(new_n219), .B1(new_n779), .B2(new_n837), .ZN(new_n1053));
  NOR3_X1   g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n298), .B(new_n987), .C1(G159), .C2(new_n788), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(new_n405), .C2(new_n836), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n434), .B1(new_n797), .B2(G326), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n772), .A2(new_n303), .B1(new_n791), .B2(new_n799), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n796), .A2(G317), .B1(G311), .B2(new_n789), .ZN(new_n1059));
  INV_X1    g0859(.A(G322), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1059), .B1(new_n1060), .B2(new_n840), .C1(new_n785), .C2(new_n603), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT48), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1058), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n1062), .B2(new_n1061), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT49), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1057), .B1(new_n559), .B2(new_n775), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1056), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1050), .B1(new_n1068), .B2(new_n764), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1013), .B2(new_n813), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT115), .Z(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n1035), .B2(new_n749), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1041), .A2(new_n1072), .ZN(G393));
  XNOR2_X1  g0873(.A(new_n1010), .B(new_n700), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n707), .B1(new_n1039), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1036), .A2(new_n1011), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n969), .B1(G97), .B2(new_n705), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n242), .A2(new_n752), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n751), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n796), .A2(G159), .B1(G150), .B2(new_n788), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT51), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n791), .A2(new_n202), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n434), .B1(new_n775), .B2(new_n268), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n772), .A2(new_n219), .B1(new_n779), .B2(new_n841), .ZN(new_n1085));
  NOR4_X1   g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n785), .A2(new_n405), .B1(new_n363), .B2(new_n836), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT117), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n757), .B1(new_n559), .B2(new_n791), .C1(new_n836), .C2(new_n603), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n772), .A2(new_n799), .B1(new_n775), .B2(new_n205), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n782), .A2(new_n303), .B1(new_n779), .B2(new_n1060), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n801), .A2(new_n840), .B1(new_n770), .B2(new_n807), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT118), .B(KEYINPUT52), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1093), .B(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1086), .A2(new_n1088), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1080), .B1(new_n835), .B2(new_n1096), .C1(new_n1021), .C2(new_n813), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n1074), .B2(new_n749), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1077), .A2(new_n1099), .ZN(G390));
  NAND2_X1  g0900(.A1(new_n952), .A2(new_n955), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n831), .A2(new_n949), .B1(new_n929), .B2(new_n937), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1101), .B1(new_n1102), .B2(new_n953), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n692), .B(new_n828), .C1(new_n719), .C2(new_n720), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n949), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n929), .A2(new_n937), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n953), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n903), .B2(new_n912), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n738), .A2(G330), .A3(new_n828), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n1106), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1103), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1109), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n671), .A2(new_n663), .A3(new_n672), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n659), .A2(new_n660), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1117), .B1(new_n1118), .B2(new_n644), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n688), .B1(new_n1119), .B2(new_n661), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n948), .B1(new_n1120), .B2(new_n828), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n929), .A2(new_n937), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1108), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1116), .B1(new_n1123), .B2(new_n1101), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n886), .A2(G330), .A3(new_n938), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1115), .B(new_n749), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1101), .A2(new_n761), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n751), .B1(new_n405), .B2(new_n861), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n379), .A2(new_n1083), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n843), .A2(G97), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(G107), .A2(new_n789), .B1(new_n788), .B2(G283), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n770), .A2(new_n559), .B1(new_n779), .B2(new_n303), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n772), .A2(new_n268), .B1(new_n775), .B2(new_n219), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AND4_X1   g0934(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .A4(new_n1134), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n792), .A2(G159), .B1(G137), .B2(new_n789), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT54), .B(G143), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1136), .B1(new_n785), .B2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT119), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n977), .A2(G150), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT53), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n776), .A2(G50), .B1(new_n797), .B2(G125), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n847), .B2(new_n770), .ZN(new_n1143));
  INV_X1    g0943(.A(G128), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n379), .B1(new_n840), .B2(new_n1144), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n1141), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1135), .B1(new_n1139), .B2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1127), .B(new_n1128), .C1(new_n835), .C2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1126), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1115), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n886), .A2(G330), .A3(new_n516), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1151), .A2(new_n679), .A3(new_n960), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n949), .B(new_n1104), .C1(new_n1122), .C2(new_n1112), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n886), .A2(G330), .A3(new_n828), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1153), .B1(new_n1122), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1122), .A2(new_n1112), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1121), .B1(new_n1125), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1152), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1150), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n707), .B1(new_n1150), .B2(new_n1158), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1149), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(G378));
  NAND2_X1  g0962(.A1(new_n408), .A2(new_n893), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n423), .A2(new_n487), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1163), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n413), .A2(new_n418), .B1(KEYINPUT10), .B2(new_n421), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n486), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1164), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n1164), .B2(new_n1167), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n761), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n750), .B1(G50), .B2(new_n862), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n836), .A2(new_n847), .B1(new_n791), .B2(new_n837), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1137), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n796), .A2(G128), .B1(new_n977), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n839), .B2(new_n782), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1174), .B(new_n1177), .C1(G125), .C2(new_n788), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n253), .B(new_n308), .C1(new_n775), .C2(new_n428), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G124), .B2(new_n797), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n779), .A2(new_n799), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n775), .A2(new_n424), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(G107), .C2(new_n796), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n575), .B2(new_n782), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n308), .B(new_n298), .C1(new_n772), .C2(new_n202), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n836), .A2(new_n204), .B1(new_n840), .B2(new_n559), .ZN(new_n1190));
  NOR4_X1   g0990(.A1(new_n1188), .A2(new_n981), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1191), .A2(KEYINPUT58), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(KEYINPUT58), .ZN(new_n1193));
  AOI21_X1  g0993(.A(G50), .B1(new_n253), .B2(new_n308), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n434), .B2(G41), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1184), .A2(new_n1192), .A3(new_n1193), .A4(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1173), .B1(new_n1196), .B2(new_n764), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1172), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT121), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n877), .B1(new_n1171), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n945), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1199), .B1(new_n1171), .B2(KEYINPUT120), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n950), .B2(new_n958), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n956), .A2(new_n957), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n831), .A2(new_n949), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n942), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n1106), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1168), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1164), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1210), .A2(KEYINPUT120), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(KEYINPUT121), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1204), .A2(new_n1207), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1203), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1201), .A2(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n945), .A2(new_n1203), .A3(new_n1200), .A4(new_n1214), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1198), .B1(new_n1218), .B2(new_n748), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  AND4_X1   g1020(.A1(new_n945), .A2(new_n1203), .A3(new_n1200), .A4(new_n1214), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n945), .A2(new_n1200), .B1(new_n1203), .B2(new_n1214), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1152), .B1(new_n1150), .B2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1223), .A2(new_n1225), .A3(KEYINPUT57), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n706), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT57), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1220), .B1(new_n1227), .B2(new_n1228), .ZN(G375));
  NAND2_X1  g1029(.A1(new_n961), .A2(new_n1151), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1224), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1231), .A2(new_n1018), .A3(new_n1158), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n298), .B(new_n1186), .C1(new_n789), .C2(new_n1175), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n782), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1234), .A2(G150), .B1(new_n977), .B2(G159), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n796), .A2(G137), .B1(new_n797), .B2(G128), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n792), .A2(G50), .B1(G132), .B2(new_n788), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1233), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n843), .A2(G107), .B1(G116), .B2(new_n789), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1239), .A2(KEYINPUT122), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1051), .B1(G283), .B2(new_n796), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1240), .B1(KEYINPUT123), .B2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(KEYINPUT123), .B2(new_n1242), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1239), .A2(KEYINPUT122), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n977), .A2(G97), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n975), .B1(G303), .B2(new_n797), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n379), .B1(G294), .B2(new_n788), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1238), .B1(new_n1244), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n764), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n751), .B1(new_n219), .B2(new_n861), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1251), .B(new_n1252), .C1(new_n1106), .C2(new_n762), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n1224), .B2(new_n748), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1232), .A2(new_n1255), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(KEYINPUT124), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(G381));
  NOR3_X1   g1058(.A1(G387), .A2(G384), .A3(G390), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1041), .A2(new_n817), .A3(new_n1072), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1259), .A2(new_n1161), .A3(new_n1257), .A4(new_n1261), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1262), .A2(G375), .ZN(G407));
  NAND2_X1  g1063(.A1(new_n687), .A2(G213), .ZN(new_n1264));
  OR3_X1    g1064(.A1(G375), .A2(G378), .A3(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(G407), .A2(G213), .A3(new_n1265), .ZN(G409));
  AND3_X1   g1066(.A1(new_n1223), .A2(new_n1018), .A3(new_n1225), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1161), .B1(new_n1267), .B2(new_n1219), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT125), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(G378), .B(new_n1220), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1271));
  OAI211_X1 g1071(.A(KEYINPUT125), .B(new_n1161), .C1(new_n1267), .C2(new_n1219), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1157), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1153), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1154), .A2(new_n1122), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1230), .A2(new_n1274), .A3(new_n1277), .A4(KEYINPUT60), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n706), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1158), .A2(KEYINPUT60), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1279), .B1(new_n1231), .B2(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n866), .B1(new_n1281), .B2(new_n1254), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1280), .A2(new_n1231), .ZN(new_n1283));
  OAI211_X1 g1083(.A(G384), .B(new_n1255), .C1(new_n1283), .C2(new_n1279), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1273), .A2(new_n1264), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(KEYINPUT62), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1273), .A2(new_n1264), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n687), .A2(G213), .A3(G2897), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1290), .B(KEYINPUT126), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1285), .B(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1289), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT62), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1273), .A2(new_n1286), .A3(new_n1295), .A4(new_n1264), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1288), .A2(new_n1293), .A3(new_n1294), .A4(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(G390), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G387), .A2(new_n1298), .ZN(new_n1299));
  OAI211_X1 g1099(.A(G390), .B(new_n999), .C1(new_n1019), .C2(new_n1033), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(G393), .A2(G396), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1260), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1301), .A2(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1299), .A2(new_n1302), .A3(new_n1300), .A4(new_n1260), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1297), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1305), .ZN(new_n1308));
  AOI22_X1  g1108(.A1(new_n1300), .A2(new_n1299), .B1(new_n1302), .B2(new_n1260), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT61), .B1(new_n1289), .B2(new_n1292), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT63), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1287), .A2(new_n1312), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1273), .A2(new_n1286), .A3(KEYINPUT63), .A4(new_n1264), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1310), .A2(new_n1311), .A3(new_n1313), .A4(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1307), .A2(new_n1315), .ZN(G405));
  OAI21_X1  g1116(.A(KEYINPUT127), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(G375), .A2(new_n1161), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1271), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1319), .A2(new_n1286), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1319), .A2(new_n1286), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT127), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1304), .A2(new_n1323), .A3(new_n1305), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1317), .A2(new_n1321), .A3(new_n1322), .A4(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1322), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1306), .B(KEYINPUT127), .C1(new_n1320), .C2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(G402));
endmodule


