//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  AOI22_X1  g0006(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G50), .A2(G226), .ZN(new_n208));
  INV_X1    g0008(.A(G77), .ZN(new_n209));
  INV_X1    g0009(.A(G244), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n207), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G97), .B2(G257), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT64), .B(G68), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n212), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n203), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(G58), .A2(G68), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n206), .B(new_n222), .C1(new_n225), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(G264), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n232), .B(new_n233), .Z(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XOR2_X1   g0036(.A(G238), .B(G244), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n234), .B(new_n238), .Z(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n223), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT16), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n226), .B1(new_n213), .B2(G58), .ZN(new_n251));
  INV_X1    g0051(.A(G159), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  OAI22_X1  g0054(.A1(new_n251), .A2(new_n224), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n213), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT7), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n257), .B1(new_n258), .B2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n256), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n250), .B1(new_n255), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT79), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g0069(.A(KEYINPUT79), .B(new_n250), .C1(new_n255), .C2(new_n266), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n249), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT77), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n264), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n261), .A2(new_n263), .A3(KEYINPUT77), .ZN(new_n274));
  AOI21_X1  g0074(.A(G20), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n265), .B1(new_n275), .B2(KEYINPUT7), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n255), .B1(new_n276), .B2(G68), .ZN(new_n277));
  AOI21_X1  g0077(.A(KEYINPUT78), .B1(new_n277), .B2(KEYINPUT16), .ZN(new_n278));
  INV_X1    g0078(.A(new_n255), .ZN(new_n279));
  AOI211_X1 g0079(.A(new_n257), .B(G20), .C1(new_n261), .C2(new_n263), .ZN(new_n280));
  AND3_X1   g0080(.A1(new_n261), .A2(new_n263), .A3(KEYINPUT77), .ZN(new_n281));
  AOI21_X1  g0081(.A(KEYINPUT77), .B1(new_n261), .B2(new_n263), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n224), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n280), .B1(new_n283), .B2(new_n257), .ZN(new_n284));
  INV_X1    g0084(.A(G68), .ZN(new_n285));
  OAI211_X1 g0085(.A(KEYINPUT16), .B(new_n279), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT78), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n271), .B1(new_n278), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT80), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT67), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G41), .A2(G45), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(G1), .ZN(new_n294));
  INV_X1    g0094(.A(G1), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n295), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n291), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n297), .A2(G232), .ZN(new_n298));
  INV_X1    g0098(.A(G41), .ZN(new_n299));
  OAI211_X1 g0099(.A(G1), .B(G13), .C1(new_n260), .C2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G223), .ZN(new_n301));
  INV_X1    g0101(.A(G1698), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n258), .B(new_n303), .C1(G226), .C2(new_n302), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G87), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n300), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n295), .B1(G41), .B2(G45), .ZN(new_n307));
  INV_X1    g0107(.A(G274), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NOR4_X1   g0109(.A1(new_n298), .A2(new_n306), .A3(G190), .A4(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n304), .A2(new_n305), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n311), .A2(new_n291), .B1(G232), .B2(new_n297), .ZN(new_n312));
  INV_X1    g0112(.A(new_n309), .ZN(new_n313));
  AOI21_X1  g0113(.A(G200), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n290), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G190), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n312), .A2(new_n316), .A3(new_n313), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n298), .A2(new_n306), .A3(new_n309), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n317), .B(KEYINPUT80), .C1(new_n318), .C2(G200), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT8), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT69), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n321), .B1(new_n322), .B2(new_n215), .ZN(new_n323));
  NAND3_X1  g0123(.A1(KEYINPUT69), .A2(KEYINPUT8), .A3(G58), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n295), .A2(G13), .A3(G20), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n249), .B1(G1), .B2(new_n224), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n327), .B1(new_n329), .B2(new_n325), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n289), .A2(new_n320), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT17), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n289), .A2(new_n330), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT18), .ZN(new_n335));
  INV_X1    g0135(.A(G169), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n318), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(G179), .B2(new_n318), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n334), .A2(new_n335), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n330), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n286), .A2(new_n287), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n276), .A2(G68), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n343), .A2(KEYINPUT78), .A3(KEYINPUT16), .A4(new_n279), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n341), .B1(new_n345), .B2(new_n271), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n346), .A2(KEYINPUT17), .A3(new_n320), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT18), .B1(new_n346), .B2(new_n338), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n333), .A2(new_n340), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n326), .A2(G77), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n328), .A2(new_n209), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G20), .A2(G77), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT15), .B(G87), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n224), .A2(G33), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT8), .B(G58), .ZN(new_n356));
  OAI221_X1 g0156(.A(new_n353), .B1(new_n354), .B2(new_n355), .C1(new_n254), .C2(new_n356), .ZN(new_n357));
  AOI211_X1 g0157(.A(new_n351), .B(new_n352), .C1(new_n248), .C2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n302), .A2(G232), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G238), .A2(G1698), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n258), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n258), .A2(G107), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT71), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT71), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n361), .B(new_n365), .C1(G107), .C2(new_n258), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(new_n291), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n294), .A2(new_n296), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT68), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n368), .A2(new_n369), .A3(new_n300), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n369), .B1(new_n368), .B2(new_n300), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n367), .B(new_n313), .C1(new_n372), .C2(new_n210), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n358), .B1(new_n373), .B2(new_n336), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT72), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n297), .B(new_n369), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n309), .B1(new_n377), .B2(G244), .ZN(new_n378));
  AOI21_X1  g0178(.A(G169), .B1(new_n378), .B2(new_n367), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT72), .B1(new_n379), .B2(new_n358), .ZN(new_n380));
  INV_X1    g0180(.A(G179), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n378), .A2(new_n381), .A3(new_n367), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n376), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n373), .A2(G200), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n384), .B(new_n358), .C1(new_n316), .C2(new_n373), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT73), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT12), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n213), .A2(new_n389), .A3(new_n326), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n285), .B1(new_n328), .B2(KEYINPUT12), .ZN(new_n391));
  AOI211_X1 g0191(.A(new_n390), .B(new_n391), .C1(new_n389), .C2(new_n326), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n213), .A2(new_n224), .ZN(new_n393));
  INV_X1    g0193(.A(G50), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n254), .A2(new_n394), .B1(new_n355), .B2(new_n209), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n248), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  XOR2_X1   g0196(.A(KEYINPUT76), .B(KEYINPUT11), .Z(new_n397));
  XNOR2_X1  g0197(.A(new_n396), .B(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n392), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(G238), .B1(new_n370), .B2(new_n371), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G97), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n216), .A2(G1698), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(G226), .B2(G1698), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n402), .B1(new_n404), .B2(new_n264), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n291), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n401), .A2(new_n313), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT13), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT13), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n401), .A2(new_n409), .A3(new_n313), .A4(new_n406), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n400), .B1(new_n411), .B2(new_n316), .ZN(new_n412));
  INV_X1    g0212(.A(G200), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n408), .B2(new_n410), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT14), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n411), .B2(G169), .ZN(new_n417));
  AOI211_X1 g0217(.A(KEYINPUT14), .B(new_n336), .C1(new_n408), .C2(new_n410), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n411), .A2(new_n381), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n415), .B1(new_n422), .B2(new_n399), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n350), .A2(new_n388), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT10), .ZN(new_n425));
  OAI21_X1  g0225(.A(G20), .B1(new_n227), .B2(G50), .ZN(new_n426));
  INV_X1    g0226(.A(G150), .ZN(new_n427));
  OAI221_X1 g0227(.A(new_n426), .B1(new_n427), .B2(new_n254), .C1(new_n325), .C2(new_n355), .ZN(new_n428));
  INV_X1    g0228(.A(new_n326), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n428), .A2(new_n248), .B1(new_n394), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n329), .A2(G50), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT9), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  XOR2_X1   g0234(.A(KEYINPUT66), .B(G226), .Z(new_n435));
  NAND2_X1  g0235(.A1(new_n377), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n300), .B1(new_n264), .B2(new_n209), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n302), .A2(G222), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n258), .B(new_n438), .C1(new_n301), .C2(new_n302), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n309), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n436), .A2(G190), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n430), .A2(KEYINPUT9), .A3(new_n431), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n434), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n436), .A2(new_n440), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G200), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n425), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(KEYINPUT74), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT74), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n444), .A2(new_n449), .A3(G200), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n443), .A2(new_n448), .A3(new_n425), .A4(new_n450), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n451), .A2(KEYINPUT75), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n451), .A2(KEYINPUT75), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n447), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n444), .A2(new_n336), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n436), .A2(new_n381), .A3(new_n440), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n432), .A3(new_n456), .ZN(new_n457));
  XNOR2_X1  g0257(.A(new_n457), .B(KEYINPUT70), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n387), .A2(KEYINPUT73), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n424), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G45), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(G1), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n308), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n219), .B1(new_n462), .B2(G1), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n300), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT83), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n464), .A2(new_n300), .A3(KEYINPUT83), .A4(new_n465), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n210), .A2(G1698), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n470), .B1(G238), .B2(G1698), .ZN(new_n471));
  INV_X1    g0271(.A(G116), .ZN(new_n472));
  OAI22_X1  g0272(.A1(new_n471), .A2(new_n264), .B1(new_n260), .B2(new_n472), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n468), .A2(new_n469), .B1(new_n473), .B2(new_n291), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G200), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT19), .ZN(new_n477));
  INV_X1    g0277(.A(G97), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n477), .B1(new_n355), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT84), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n258), .A2(new_n224), .A3(G68), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n224), .B1(new_n402), .B2(new_n477), .ZN(new_n482));
  NOR2_X1   g0282(.A1(G97), .A2(G107), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n218), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT84), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n486), .B(new_n477), .C1(new_n355), .C2(new_n478), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n480), .A2(new_n481), .A3(new_n485), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n248), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n249), .B(new_n326), .C1(G1), .C2(new_n260), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G87), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n354), .A2(new_n429), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n489), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n474), .A2(G190), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n476), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n475), .A2(new_n336), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n474), .A2(new_n381), .ZN(new_n498));
  XOR2_X1   g0298(.A(new_n354), .B(KEYINPUT85), .Z(new_n499));
  OAI211_X1 g0299(.A(new_n489), .B(new_n493), .C1(new_n490), .C2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g0302(.A1(KEYINPUT5), .A2(G41), .ZN(new_n503));
  NOR2_X1   g0303(.A1(KEYINPUT5), .A2(G41), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n463), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n300), .ZN(new_n506));
  INV_X1    g0306(.A(G257), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n210), .A2(G1698), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT82), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT4), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n509), .A2(new_n512), .A3(new_n261), .A4(new_n263), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n510), .B2(new_n511), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G283), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n258), .A2(G250), .A3(G1698), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n258), .A2(KEYINPUT82), .A3(KEYINPUT4), .A4(new_n509), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n514), .A2(new_n515), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n508), .B1(new_n518), .B2(new_n291), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n463), .B(G274), .C1(new_n504), .C2(new_n503), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G200), .ZN(new_n522));
  INV_X1    g0322(.A(new_n520), .ZN(new_n523));
  AOI211_X1 g0323(.A(new_n523), .B(new_n508), .C1(new_n518), .C2(new_n291), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G190), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT81), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n326), .A2(G97), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT7), .B1(new_n264), .B2(new_n224), .ZN(new_n528));
  OAI21_X1  g0328(.A(G107), .B1(new_n528), .B2(new_n280), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT6), .ZN(new_n530));
  AND2_X1   g0330(.A1(G97), .A2(G107), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(new_n483), .ZN(new_n532));
  INV_X1    g0332(.A(G107), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(KEYINPUT6), .A3(G97), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n535), .A2(G20), .B1(G77), .B2(new_n253), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n529), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n527), .B1(new_n537), .B2(new_n248), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n491), .A2(G97), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n526), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n535), .A2(G20), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n253), .A2(G77), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n533), .B1(new_n259), .B2(new_n265), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n248), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n527), .ZN(new_n546));
  AND4_X1   g0346(.A1(new_n526), .A2(new_n545), .A3(new_n539), .A4(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n522), .B(new_n525), .C1(new_n540), .C2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n518), .A2(new_n291), .ZN(new_n549));
  INV_X1    g0349(.A(new_n508), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n549), .A2(G179), .A3(new_n520), .A4(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n524), .B2(new_n336), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n545), .A2(new_n539), .A3(new_n546), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n548), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n515), .B(new_n224), .C1(G33), .C2(new_n478), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT87), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n247), .A2(new_n223), .B1(G20), .B2(new_n472), .ZN(new_n558));
  AOI21_X1  g0358(.A(G20), .B1(new_n260), .B2(G97), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT87), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n560), .A3(new_n515), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n557), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT20), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n557), .A2(new_n561), .A3(KEYINPUT20), .A4(new_n558), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(KEYINPUT88), .A3(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n326), .A2(G116), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(new_n491), .B2(G116), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT88), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n562), .A2(new_n569), .A3(new_n563), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n566), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G264), .A2(G1698), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n258), .B(new_n573), .C1(new_n507), .C2(G1698), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n574), .B(new_n291), .C1(G303), .C2(new_n258), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n505), .A2(G270), .A3(new_n300), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(KEYINPUT86), .A3(new_n520), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT86), .B1(new_n576), .B2(new_n520), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G200), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n572), .B(new_n581), .C1(new_n316), .C2(new_n580), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n576), .A2(new_n520), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT86), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n577), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n571), .A2(G179), .A3(new_n575), .A4(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n336), .B1(new_n586), .B2(new_n575), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT21), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n588), .A2(new_n589), .A3(new_n571), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n589), .B1(new_n588), .B2(new_n571), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n582), .B(new_n587), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n555), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n429), .A2(KEYINPUT25), .A3(new_n533), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(KEYINPUT25), .B1(new_n429), .B2(new_n533), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n490), .A2(new_n533), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(G264), .ZN(new_n598));
  OAI21_X1  g0398(.A(KEYINPUT90), .B1(new_n506), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT90), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n505), .A2(new_n600), .A3(G264), .A4(new_n300), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n258), .B1(G257), .B2(new_n302), .ZN(new_n602));
  NOR2_X1   g0402(.A1(G250), .A2(G1698), .ZN(new_n603));
  INV_X1    g0403(.A(G294), .ZN(new_n604));
  OAI22_X1  g0404(.A1(new_n602), .A2(new_n603), .B1(new_n260), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n599), .A2(new_n601), .B1(new_n605), .B2(new_n291), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n413), .B1(new_n606), .B2(new_n520), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT24), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n261), .A2(new_n263), .A3(new_n224), .A4(G87), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT22), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT22), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n258), .A2(new_n611), .A3(new_n224), .A4(G87), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n224), .A2(G107), .ZN(new_n614));
  XNOR2_X1  g0414(.A(new_n614), .B(KEYINPUT23), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n260), .A2(new_n472), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n224), .ZN(new_n617));
  AND4_X1   g0417(.A1(new_n608), .A2(new_n613), .A3(new_n615), .A4(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n610), .A2(new_n612), .B1(new_n224), .B2(new_n616), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n608), .B1(new_n619), .B2(new_n615), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n248), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT89), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT89), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n623), .B(new_n248), .C1(new_n618), .C2(new_n620), .ZN(new_n624));
  AOI211_X1 g0424(.A(new_n597), .B(new_n607), .C1(new_n622), .C2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n606), .A2(new_n520), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(G190), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n622), .A2(new_n624), .ZN(new_n629));
  INV_X1    g0429(.A(new_n597), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n626), .A2(new_n336), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(G179), .B2(new_n626), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n625), .A2(new_n628), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  AND4_X1   g0435(.A1(new_n461), .A2(new_n502), .A3(new_n593), .A4(new_n635), .ZN(G372));
  NAND2_X1  g0436(.A1(new_n422), .A2(new_n399), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n415), .B1(new_n637), .B2(new_n383), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n638), .A2(new_n333), .A3(new_n347), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT92), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n335), .B1(new_n334), .B2(new_n339), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n346), .A2(KEYINPUT18), .A3(new_n338), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n340), .A2(new_n348), .A3(KEYINPUT92), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n454), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n458), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  OR3_X1    g0449(.A1(new_n424), .A2(new_n459), .A3(new_n460), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n571), .A2(G169), .A3(new_n580), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT21), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n588), .A2(new_n589), .A3(new_n571), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n597), .B1(new_n622), .B2(new_n624), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n654), .B(new_n587), .C1(new_n655), .C2(new_n633), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n655), .B(new_n628), .C1(new_n413), .C2(new_n627), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n553), .A2(KEYINPUT81), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n538), .A2(new_n526), .A3(new_n539), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n658), .A2(new_n659), .B1(G190), .B2(new_n524), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n660), .A2(new_n522), .B1(new_n552), .B2(new_n553), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT91), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n494), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n494), .A2(new_n662), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n476), .B(new_n495), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n656), .A2(new_n657), .A3(new_n661), .A4(new_n665), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n552), .A2(new_n658), .A3(new_n659), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n501), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n552), .A2(new_n496), .A3(new_n501), .A4(new_n553), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(KEYINPUT26), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n649), .B1(new_n650), .B2(new_n674), .ZN(G369));
  NAND2_X1  g0475(.A1(new_n654), .A2(new_n587), .ZN(new_n676));
  INV_X1    g0476(.A(G13), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(G20), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n295), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n680), .A2(G213), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G343), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT93), .Z(new_n684));
  NAND2_X1  g0484(.A1(new_n676), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT94), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n631), .A2(new_n634), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n657), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n655), .A2(new_n684), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n686), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n689), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n635), .A2(KEYINPUT94), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n685), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n684), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n687), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n631), .A2(new_n634), .A3(new_n694), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n690), .A2(new_n692), .A3(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n684), .A2(new_n572), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n676), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n592), .B2(new_n699), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G330), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n696), .A2(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n204), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n484), .A2(G116), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n228), .B2(new_n708), .ZN(new_n711));
  XOR2_X1   g0511(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n712));
  XNOR2_X1  g0512(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n635), .A2(new_n593), .A3(new_n502), .A4(new_n684), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n519), .A2(G179), .A3(new_n474), .A4(new_n520), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n606), .A2(new_n586), .A3(new_n575), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n716), .A2(KEYINPUT30), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n715), .B2(new_n717), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n474), .A2(G179), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n521), .A2(new_n626), .A3(new_n580), .A4(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n719), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n694), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT31), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT31), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n724), .A2(new_n727), .A3(new_n694), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n714), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G330), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n668), .B1(new_n667), .B2(new_n665), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n501), .B1(new_n671), .B2(KEYINPUT26), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n694), .B1(new_n666), .B2(new_n735), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n736), .A2(KEYINPUT96), .A3(KEYINPUT29), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT96), .B1(new_n736), .B2(KEYINPUT29), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n694), .B1(new_n666), .B2(new_n673), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n740), .A2(KEYINPUT29), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n732), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n713), .B1(new_n742), .B2(G1), .ZN(G364));
  AOI21_X1  g0543(.A(new_n223), .B1(G20), .B2(new_n336), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n224), .A2(new_n316), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n381), .A2(G200), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n215), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n413), .A2(G179), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n751), .A2(KEYINPUT100), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(KEYINPUT100), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n224), .A2(G190), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G179), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n252), .ZN(new_n758));
  XNOR2_X1  g0558(.A(KEYINPUT99), .B(KEYINPUT32), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n754), .A2(new_n218), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n224), .B1(new_n756), .B2(G190), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n478), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n755), .A2(new_n750), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G107), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n755), .A2(new_n747), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n765), .B1(new_n209), .B2(new_n766), .ZN(new_n767));
  OR4_X1    g0567(.A1(new_n749), .A2(new_n760), .A3(new_n762), .A4(new_n767), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n264), .B(new_n768), .C1(new_n758), .C2(new_n759), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n381), .A2(new_n413), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n770), .A2(new_n746), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n770), .A2(new_n755), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n769), .B1(new_n394), .B2(new_n772), .C1(new_n285), .C2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n766), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G283), .A2(new_n764), .B1(new_n776), .B2(G311), .ZN(new_n777));
  INV_X1    g0577(.A(G326), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n777), .B(new_n264), .C1(new_n778), .C2(new_n772), .ZN(new_n779));
  INV_X1    g0579(.A(new_n754), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n779), .B1(G303), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n761), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G294), .ZN(new_n783));
  INV_X1    g0583(.A(new_n748), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G322), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT33), .B(G317), .ZN(new_n786));
  INV_X1    g0586(.A(new_n757), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n773), .A2(new_n786), .B1(new_n787), .B2(G329), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n781), .A2(new_n783), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n745), .B1(new_n775), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n701), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n790), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n273), .A2(new_n274), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n204), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT97), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n229), .A2(new_n462), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n799), .B(new_n800), .C1(new_n462), .C2(new_n242), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n706), .A2(new_n264), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G355), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n801), .B(new_n803), .C1(G116), .C2(new_n204), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n793), .A2(new_n744), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT98), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n678), .A2(G45), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n708), .A2(G1), .A3(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n796), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n701), .A2(G330), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n812), .A2(new_n702), .A3(new_n809), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n811), .A2(new_n813), .ZN(G396));
  NAND2_X1  g0614(.A1(new_n386), .A2(KEYINPUT102), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT102), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n383), .A2(new_n816), .A3(new_n385), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n740), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n684), .A2(new_n358), .ZN(new_n820));
  AND3_X1   g0620(.A1(new_n383), .A2(new_n816), .A3(new_n385), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n816), .B1(new_n383), .B2(new_n385), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n820), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n815), .A2(new_n824), .A3(new_n817), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n819), .B1(new_n826), .B2(new_n740), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(new_n732), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n809), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n826), .A2(new_n792), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n363), .B1(new_n754), .B2(new_n264), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT101), .Z(new_n832));
  AOI21_X1  g0632(.A(new_n762), .B1(G311), .B2(new_n787), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n472), .B2(new_n766), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n771), .A2(G303), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n763), .A2(new_n218), .ZN(new_n836));
  NOR4_X1   g0636(.A1(new_n832), .A2(new_n834), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G283), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n837), .B1(new_n838), .B2(new_n774), .C1(new_n604), .C2(new_n748), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G143), .A2(new_n784), .B1(new_n776), .B2(G159), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n771), .A2(G137), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n840), .B(new_n841), .C1(new_n427), .C2(new_n774), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT34), .Z(new_n843));
  INV_X1    g0643(.A(G132), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n754), .A2(new_n394), .B1(new_n844), .B2(new_n757), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n843), .A2(new_n797), .A3(new_n845), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n846), .B1(new_n215), .B2(new_n761), .C1(new_n285), .C2(new_n763), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n745), .B1(new_n839), .B2(new_n847), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n830), .A2(new_n809), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n744), .A2(new_n791), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n849), .B1(G77), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n829), .A2(new_n852), .ZN(G384));
  OR2_X1    g0653(.A1(new_n412), .A2(new_n414), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n694), .A2(new_n399), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n417), .A2(new_n418), .A3(new_n420), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n854), .B(new_n855), .C1(new_n856), .C2(new_n400), .ZN(new_n857));
  INV_X1    g0657(.A(new_n855), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n422), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  AND4_X1   g0660(.A1(new_n730), .A2(new_n860), .A3(new_n825), .A4(new_n823), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT105), .ZN(new_n862));
  INV_X1    g0662(.A(new_n682), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n346), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n862), .B1(new_n346), .B2(new_n863), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n340), .A2(KEYINPUT92), .A3(new_n348), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT92), .B1(new_n340), .B2(new_n348), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n331), .A2(new_n332), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT17), .B1(new_n346), .B2(new_n320), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT106), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT106), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n333), .A2(new_n875), .A3(new_n347), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n868), .B1(new_n871), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT105), .B1(new_n334), .B2(new_n682), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n331), .B1(new_n879), .B2(new_n864), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n334), .A2(KEYINPUT92), .A3(new_n339), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n640), .B1(new_n346), .B2(new_n338), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT37), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT37), .B1(new_n334), .B2(new_n339), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n331), .B(new_n885), .C1(new_n879), .C2(new_n864), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT38), .B1(new_n878), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n343), .A2(new_n279), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n342), .A2(new_n344), .B1(new_n250), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n341), .B1(new_n890), .B2(new_n248), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n331), .B1(new_n891), .B2(new_n863), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n338), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT37), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n886), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n891), .A2(new_n863), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n349), .A2(new_n896), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n895), .A2(KEYINPUT38), .A3(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(KEYINPUT40), .B(new_n861), .C1(new_n888), .C2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n895), .B2(new_n897), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n861), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n899), .A2(G330), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n461), .A2(new_n732), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT109), .Z(new_n907));
  NAND3_X1  g0707(.A1(new_n899), .A2(new_n730), .A3(new_n903), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n907), .B1(new_n650), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n888), .B2(new_n898), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n898), .A2(new_n900), .A3(new_n910), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n422), .A2(new_n399), .A3(new_n684), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n911), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n898), .A2(new_n900), .ZN(new_n917));
  INV_X1    g0717(.A(new_n860), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n383), .A2(new_n694), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n918), .B1(new_n819), .B2(new_n919), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n917), .A2(new_n920), .B1(new_n871), .B2(new_n863), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n916), .A2(KEYINPUT107), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT107), .B1(new_n916), .B2(new_n921), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n666), .A2(new_n735), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(KEYINPUT29), .A3(new_n684), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT96), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n736), .A2(KEYINPUT96), .A3(KEYINPUT29), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(new_n741), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT108), .B1(new_n930), .B2(new_n650), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT108), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n739), .A2(new_n932), .A3(new_n461), .A4(new_n741), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n648), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n924), .B(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n909), .B(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n295), .B2(new_n678), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n209), .B(new_n228), .C1(new_n213), .C2(G58), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n285), .A2(G50), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT104), .ZN(new_n940));
  OAI211_X1 g0740(.A(G1), .B(new_n677), .C1(new_n938), .C2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n472), .B1(new_n535), .B2(KEYINPUT35), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n942), .B(new_n225), .C1(KEYINPUT35), .C2(new_n535), .ZN(new_n943));
  XOR2_X1   g0743(.A(KEYINPUT103), .B(KEYINPUT36), .Z(new_n944));
  XNOR2_X1  g0744(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n937), .A2(new_n941), .A3(new_n945), .ZN(G367));
  NAND3_X1  g0746(.A1(new_n694), .A2(new_n658), .A3(new_n659), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n661), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n667), .A2(new_n694), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n704), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n663), .A2(new_n664), .ZN(new_n953));
  OR3_X1    g0753(.A1(new_n953), .A2(new_n670), .A3(new_n684), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n670), .B1(new_n953), .B2(new_n684), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n954), .A2(new_n665), .A3(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT110), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(KEYINPUT111), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n958), .A2(KEYINPUT111), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT112), .ZN(new_n963));
  INV_X1    g0763(.A(new_n957), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n963), .B1(new_n964), .B2(new_n958), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n957), .A2(KEYINPUT112), .A3(KEYINPUT43), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n693), .ZN(new_n968));
  OAI21_X1  g0768(.A(KEYINPUT42), .B1(new_n968), .B2(new_n555), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n554), .B1(new_n951), .B2(new_n687), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n684), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT42), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n693), .A2(new_n972), .A3(new_n661), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n969), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n962), .B1(new_n967), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n967), .A2(new_n974), .A3(new_n962), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n952), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n977), .ZN(new_n979));
  INV_X1    g0779(.A(new_n952), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n979), .A2(new_n980), .A3(new_n975), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n707), .B(KEYINPUT41), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n704), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n951), .B1(new_n693), .B2(new_n695), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n986), .A2(KEYINPUT44), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(KEYINPUT44), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT45), .B1(new_n696), .B2(new_n950), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT45), .ZN(new_n991));
  NOR4_X1   g0791(.A1(new_n693), .A2(new_n991), .A3(new_n695), .A4(new_n951), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n985), .B1(new_n989), .B2(new_n993), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n690), .A2(new_n692), .A3(new_n697), .A4(new_n685), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n995), .A2(KEYINPUT113), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(KEYINPUT113), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n968), .A2(new_n702), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n998), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n702), .B1(new_n1001), .B2(new_n996), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n742), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n696), .A2(new_n950), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n991), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n992), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1008), .A2(new_n704), .A3(new_n988), .A4(new_n987), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n994), .A2(new_n1004), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n984), .B1(new_n1010), .B2(new_n742), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n808), .A2(G1), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n982), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n809), .B1(new_n964), .B2(new_n793), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n799), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n806), .B1(new_n204), .B2(new_n354), .C1(new_n1015), .C2(new_n234), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n774), .A2(new_n252), .B1(new_n766), .B2(new_n394), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G150), .A2(new_n784), .B1(new_n787), .B2(G137), .ZN(new_n1018));
  INV_X1    g0818(.A(G143), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1018), .B1(new_n1019), .B2(new_n772), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1017), .B(new_n1020), .C1(G77), .C2(new_n764), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n782), .A2(G68), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n780), .A2(G58), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1021), .A2(new_n258), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n780), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT46), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n754), .B2(new_n472), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1025), .B(new_n1027), .C1(new_n604), .C2(new_n774), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT114), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G303), .A2(new_n784), .B1(new_n776), .B2(G283), .ZN(new_n1031));
  INV_X1    g0831(.A(G311), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1031), .B1(new_n1032), .B2(new_n772), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n787), .A2(G317), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n797), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G97), .B2(new_n764), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1030), .A2(new_n1034), .A3(new_n1035), .A4(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n761), .A2(new_n533), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1024), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT47), .Z(new_n1041));
  OAI211_X1 g0841(.A(new_n1014), .B(new_n1016), .C1(new_n745), .C2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1013), .A2(new_n1042), .ZN(G387));
  AOI21_X1  g0843(.A(new_n742), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1044));
  OR3_X1    g0844(.A1(new_n1004), .A2(new_n1044), .A3(new_n708), .ZN(new_n1045));
  AND3_X1   g0845(.A1(new_n1002), .A2(new_n1000), .A3(new_n1012), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G322), .A2(new_n771), .B1(new_n773), .B2(G311), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n776), .A2(G303), .ZN(new_n1048));
  INV_X1    g0848(.A(G317), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1047), .B(new_n1048), .C1(new_n1049), .C2(new_n748), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT48), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n838), .B2(new_n761), .C1(new_n604), .C2(new_n754), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT49), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1036), .B1(G116), .B2(new_n764), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1053), .B(new_n1054), .C1(new_n778), .C2(new_n757), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n499), .A2(new_n761), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n766), .A2(new_n285), .B1(new_n757), .B2(new_n427), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n774), .A2(new_n325), .B1(new_n478), .B2(new_n763), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n780), .A2(G77), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n771), .A2(G159), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n797), .B1(G50), .B2(new_n784), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n745), .B1(new_n1055), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n709), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1065), .A2(new_n802), .B1(new_n533), .B2(new_n706), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n238), .A2(G45), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT115), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n356), .A2(G50), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT50), .ZN(new_n1070));
  AOI21_X1  g0870(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1070), .A2(new_n709), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n799), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1066), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n809), .B(new_n1064), .C1(new_n806), .C2(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT116), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n698), .A2(new_n794), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1046), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1045), .A2(new_n1078), .ZN(G393));
  OAI221_X1 g0879(.A(new_n806), .B1(new_n478), .B2(new_n204), .C1(new_n1015), .C2(new_n245), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n784), .A2(G159), .B1(new_n771), .B2(G150), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT51), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n1019), .A2(new_n757), .B1(new_n761), .B2(new_n209), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n766), .A2(new_n356), .ZN(new_n1084));
  OR3_X1    g0884(.A1(new_n797), .A2(new_n836), .A3(new_n1084), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1086), .B1(new_n394), .B2(new_n774), .C1(new_n256), .C2(new_n754), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n772), .A2(new_n1049), .B1(new_n748), .B2(new_n1032), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT52), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n780), .A2(G283), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n258), .B1(new_n787), .B2(G322), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1089), .A2(new_n765), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n766), .A2(new_n604), .B1(new_n761), .B2(new_n472), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G303), .B2(new_n773), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT117), .Z(new_n1095));
  OAI21_X1  g0895(.A(new_n1087), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n809), .B1(new_n1096), .B2(new_n744), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1080), .B(new_n1097), .C1(new_n950), .C2(new_n794), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n994), .A2(new_n1009), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1012), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n708), .B1(new_n1099), .B2(new_n1003), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1101), .B1(new_n1010), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(G390));
  NAND4_X1  g0904(.A1(new_n826), .A2(G330), .A3(new_n730), .A4(new_n860), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n920), .A2(new_n915), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n911), .B2(new_n913), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n898), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n645), .A2(new_n874), .A3(new_n876), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1110), .A2(new_n868), .B1(new_n886), .B2(new_n884), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1109), .B1(new_n1111), .B2(KEYINPUT38), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n736), .A2(new_n818), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n919), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n860), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n914), .B(KEYINPUT118), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1112), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1106), .B1(new_n1108), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1112), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n912), .B1(new_n1112), .B2(new_n910), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1105), .B(new_n1119), .C1(new_n1120), .C2(new_n1107), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n931), .A2(new_n933), .ZN(new_n1123));
  AND3_X1   g0923(.A1(new_n1123), .A2(new_n649), .A3(new_n905), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n730), .A2(G330), .A3(new_n825), .A4(new_n823), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n918), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1105), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n819), .A2(new_n919), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(KEYINPUT119), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n1127), .A2(new_n1114), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT119), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1127), .A2(new_n1132), .A3(new_n1128), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1130), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1124), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1122), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1118), .A2(new_n1124), .A3(new_n1121), .A4(new_n1134), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1136), .A2(new_n707), .A3(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1118), .A2(new_n1012), .A3(new_n1121), .ZN(new_n1139));
  OR2_X1    g0939(.A1(new_n1120), .A2(new_n792), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n850), .A2(new_n325), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n264), .B1(new_n604), .B2(new_n757), .C1(new_n754), .C2(new_n218), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n748), .A2(new_n472), .B1(new_n761), .B2(new_n209), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT121), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n774), .A2(new_n533), .B1(new_n763), .B2(new_n285), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n1142), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n838), .B2(new_n772), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(G97), .B2(new_n776), .ZN(new_n1148));
  OR3_X1    g0948(.A1(new_n754), .A2(KEYINPUT53), .A3(new_n427), .ZN(new_n1149));
  OAI21_X1  g0949(.A(KEYINPUT53), .B1(new_n754), .B2(new_n427), .ZN(new_n1150));
  INV_X1    g0950(.A(G125), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1149), .B(new_n1150), .C1(new_n1151), .C2(new_n757), .ZN(new_n1152));
  XOR2_X1   g0952(.A(KEYINPUT54), .B(G143), .Z(new_n1153));
  AOI22_X1  g0953(.A1(new_n776), .A2(new_n1153), .B1(new_n773), .B2(G137), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT120), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G50), .A2(new_n764), .B1(new_n771), .B2(G128), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(new_n258), .A3(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n748), .A2(new_n844), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n761), .A2(new_n252), .ZN(new_n1159));
  NOR4_X1   g0959(.A1(new_n1152), .A2(new_n1157), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n744), .B1(new_n1148), .B2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1140), .A2(new_n810), .A3(new_n1141), .A4(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT122), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1139), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1163), .B1(new_n1139), .B2(new_n1162), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1138), .B1(new_n1164), .B2(new_n1165), .ZN(G378));
  AND4_X1   g0966(.A1(KEYINPUT125), .A2(new_n1123), .A3(new_n649), .A4(new_n905), .ZN(new_n1167));
  AOI21_X1  g0967(.A(KEYINPUT125), .B1(new_n934), .B2(new_n905), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1137), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n916), .A2(new_n921), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT107), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n916), .A2(KEYINPUT107), .A3(new_n921), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT124), .B(KEYINPUT56), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n432), .A2(new_n682), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT55), .Z(new_n1178));
  INV_X1    g0978(.A(new_n454), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n457), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1179), .A2(new_n1180), .A3(new_n1178), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1176), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1183), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1185), .A2(new_n1175), .A3(new_n1181), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1187), .A2(new_n899), .A3(G330), .A4(new_n903), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1187), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n904), .A2(new_n1189), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1173), .A2(new_n1174), .A3(new_n1188), .A4(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1188), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n923), .B2(new_n922), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1170), .A2(KEYINPUT57), .A3(new_n1191), .A4(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n707), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1192), .A2(new_n922), .A3(new_n923), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n1173), .A2(new_n1174), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT57), .B1(new_n1198), .B2(new_n1170), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1193), .A2(new_n1191), .A3(new_n1012), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1060), .B1(new_n838), .B2(new_n757), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1022), .B1(new_n774), .B2(new_n478), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n797), .B1(new_n499), .B2(new_n766), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n772), .A2(new_n472), .B1(new_n763), .B2(new_n215), .ZN(new_n1205));
  NOR4_X1   g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1206), .B(new_n299), .C1(new_n533), .C2(new_n748), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT58), .ZN(new_n1208));
  AOI21_X1  g1008(.A(G41), .B1(new_n1036), .B2(G33), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n761), .A2(new_n427), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n776), .A2(G137), .B1(new_n773), .B2(G132), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT123), .ZN(new_n1212));
  INV_X1    g1012(.A(G128), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1212), .B1(new_n1151), .B2(new_n772), .C1(new_n1213), .C2(new_n748), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1210), .B(new_n1214), .C1(new_n780), .C2(new_n1153), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT59), .ZN(new_n1216));
  AOI21_X1  g1016(.A(G33), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(G41), .B1(new_n787), .B2(G124), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1217), .B(new_n1218), .C1(new_n252), .C2(new_n763), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1208), .B1(G50), .B2(new_n1209), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n809), .B1(new_n1221), .B2(new_n744), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1222), .B1(G50), .B2(new_n851), .C1(new_n1187), .C2(new_n792), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1201), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1200), .A2(new_n1225), .ZN(G375));
  AND3_X1   g1026(.A1(new_n1130), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n934), .A2(new_n905), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1229), .A2(new_n1135), .A3(new_n983), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1056), .B1(G303), .B2(new_n787), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n258), .B1(new_n771), .B2(G294), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1231), .B(new_n1232), .C1(new_n478), .C2(new_n754), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n766), .A2(new_n533), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n748), .A2(new_n838), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n774), .A2(new_n472), .B1(new_n763), .B2(new_n209), .ZN(new_n1236));
  NOR4_X1   g1036(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n772), .A2(new_n844), .B1(new_n763), .B2(new_n215), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(G137), .B2(new_n784), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1239), .B1(new_n394), .B2(new_n761), .C1(new_n252), .C2(new_n754), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n757), .A2(new_n1213), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n766), .A2(new_n427), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1153), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1036), .B1(new_n774), .B2(new_n1243), .ZN(new_n1244));
  NOR4_X1   g1044(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .A4(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n744), .B1(new_n1237), .B2(new_n1245), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n810), .B(new_n1246), .C1(new_n860), .C2(new_n792), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n285), .B2(new_n850), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n1134), .B2(new_n1012), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1230), .A2(new_n1249), .ZN(G381));
  AND2_X1   g1050(.A1(new_n1139), .A2(new_n1162), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1138), .A2(new_n1251), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(G375), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(G384), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1230), .A2(new_n1254), .A3(new_n1249), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1013), .A2(new_n1103), .A3(new_n1042), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1045), .A2(new_n811), .A3(new_n813), .A4(new_n1078), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1253), .A2(new_n1256), .A3(new_n1259), .ZN(G407));
  INV_X1    g1060(.A(KEYINPUT126), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1253), .A2(new_n1256), .A3(new_n1259), .ZN(new_n1262));
  INV_X1    g1062(.A(G343), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1252), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1200), .A2(new_n1263), .A3(new_n1225), .A4(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(G213), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1261), .B1(new_n1262), .B2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(G407), .A2(KEYINPUT126), .A3(G213), .A4(new_n1265), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(G409));
  INV_X1    g1069(.A(KEYINPUT61), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(G393), .A2(G396), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1258), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n1013), .A2(new_n1103), .A3(new_n1042), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1103), .B1(new_n1013), .B2(new_n1042), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1273), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G387), .A2(G390), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(new_n1257), .A3(new_n1272), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1263), .A2(G213), .ZN(new_n1280));
  OAI211_X1 g1080(.A(G378), .B(new_n1225), .C1(new_n1195), .C2(new_n1199), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1198), .A2(new_n983), .A3(new_n1170), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1264), .B1(new_n1282), .B2(new_n1224), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1280), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1227), .A2(KEYINPUT60), .A3(new_n1228), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(new_n707), .A3(new_n1135), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT60), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1249), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1254), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT60), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1229), .A2(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1291), .A2(new_n707), .A3(new_n1135), .A4(new_n1285), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(G384), .A3(new_n1249), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1289), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1280), .A2(G2897), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1289), .A2(new_n1293), .A3(new_n1295), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1270), .B(new_n1279), .C1(new_n1284), .C2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  AOI211_X1 g1101(.A(new_n1280), .B(new_n1294), .C1(new_n1281), .C2(new_n1283), .ZN(new_n1302));
  OAI21_X1  g1102(.A(KEYINPUT63), .B1(new_n1302), .B2(KEYINPUT127), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1294), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1284), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT127), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT63), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1305), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1301), .A2(new_n1303), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT62), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1284), .A2(new_n1310), .A3(new_n1304), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1270), .B1(new_n1284), .B2(new_n1299), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1310), .B1(new_n1284), .B2(new_n1304), .ZN(new_n1313));
  NOR3_X1   g1113(.A1(new_n1311), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1309), .B1(new_n1314), .B2(new_n1279), .ZN(G405));
  INV_X1    g1115(.A(new_n1279), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(G375), .A2(new_n1264), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1317), .A2(new_n1281), .A3(new_n1294), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1294), .B1(new_n1317), .B2(new_n1281), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1316), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1320), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1322), .A2(new_n1318), .A3(new_n1279), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1321), .A2(new_n1323), .ZN(G402));
endmodule


