//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1199, new_n1200, new_n1201,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  XOR2_X1   g0005(.A(KEYINPUT65), .B(G244), .Z(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(new_n202), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G107), .A2(G264), .ZN(new_n211));
  NAND4_X1  g0011(.A1(new_n208), .A2(new_n209), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n205), .B1(new_n207), .B2(new_n212), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n217), .A2(G20), .A3(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n205), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XOR2_X1   g0022(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n223));
  XNOR2_X1  g0023(.A(new_n222), .B(new_n223), .ZN(new_n224));
  AND4_X1   g0024(.A1(new_n214), .A2(new_n215), .A3(new_n220), .A4(new_n224), .ZN(G361));
  XNOR2_X1  g0025(.A(G250), .B(G257), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT66), .ZN(new_n227));
  XOR2_X1   g0027(.A(G264), .B(G270), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n229), .B(new_n234), .Z(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(G50), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n239), .A2(G68), .ZN(new_n240));
  INV_X1    g0040(.A(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n238), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT16), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT78), .B(KEYINPUT7), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT3), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n248), .B1(new_n253), .B2(G20), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G20), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n241), .B1(new_n254), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G58), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(new_n241), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G58), .A2(G68), .ZN(new_n263));
  OAI21_X1  g0063(.A(G20), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G159), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n247), .B1(new_n260), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n218), .B1(new_n205), .B2(new_n250), .ZN(new_n269));
  OAI21_X1  g0069(.A(KEYINPUT77), .B1(new_n255), .B2(new_n256), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT77), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n251), .A2(new_n271), .A3(new_n252), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(new_n272), .A3(new_n258), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT7), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OR3_X1    g0075(.A1(new_n253), .A2(new_n248), .A3(G20), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n241), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n267), .A2(new_n247), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n268), .B(new_n269), .C1(new_n277), .C2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n261), .A2(KEYINPUT8), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT8), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G58), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(KEYINPUT69), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT69), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n286), .B1(new_n281), .B2(new_n283), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G1), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G20), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(G13), .A3(G20), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT70), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT70), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n294), .A2(new_n289), .A3(G13), .A4(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n269), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n291), .A2(new_n298), .B1(new_n296), .B2(new_n288), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n280), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n289), .B1(G41), .B2(G45), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G41), .ZN(new_n304));
  OAI211_X1 g0104(.A(G1), .B(G13), .C1(new_n250), .C2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n305), .A3(G274), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n302), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n306), .B1(new_n307), .B2(new_n231), .ZN(new_n308));
  INV_X1    g0108(.A(G226), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G1698), .ZN(new_n310));
  OAI221_X1 g0110(.A(new_n310), .B1(G223), .B2(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G87), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n305), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G179), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(new_n314), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n301), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT18), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT18), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n301), .A2(new_n320), .A3(new_n317), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G200), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n314), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G190), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n308), .A2(new_n313), .A3(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n327), .A2(new_n280), .A3(new_n300), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT17), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n327), .A2(new_n280), .A3(KEYINPUT17), .A4(new_n300), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n322), .A2(new_n332), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n284), .A2(new_n265), .B1(G20), .B2(G77), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n258), .A2(G33), .ZN(new_n335));
  XOR2_X1   g0135(.A(KEYINPUT15), .B(G87), .Z(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n334), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n296), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n338), .A2(new_n269), .B1(new_n202), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n298), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n341), .A2(G77), .A3(new_n290), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n231), .A2(G1698), .ZN(new_n344));
  INV_X1    g0144(.A(G238), .ZN(new_n345));
  INV_X1    g0145(.A(G1698), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n253), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G107), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n349), .B2(new_n253), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT72), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n305), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n351), .B2(new_n350), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n307), .A2(new_n206), .ZN(new_n354));
  INV_X1    g0154(.A(new_n306), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n343), .B1(new_n358), .B2(G190), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n323), .B2(new_n358), .ZN(new_n360));
  INV_X1    g0160(.A(G179), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n357), .A2(new_n316), .B1(new_n342), .B2(new_n340), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT73), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n306), .B1(new_n307), .B2(new_n309), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n253), .A2(G1698), .ZN(new_n370));
  INV_X1    g0170(.A(G223), .ZN(new_n371));
  OAI22_X1  g0171(.A1(new_n370), .A2(new_n371), .B1(new_n202), .B2(new_n253), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n257), .A2(G1698), .ZN(new_n373));
  AOI21_X1  g0173(.A(KEYINPUT67), .B1(new_n373), .B2(G222), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(KEYINPUT67), .A3(G222), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n372), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT68), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n369), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI211_X1 g0179(.A(KEYINPUT68), .B(new_n372), .C1(new_n375), .C2(new_n376), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n368), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n381), .A2(G179), .ZN(new_n382));
  INV_X1    g0182(.A(G150), .ZN(new_n383));
  INV_X1    g0183(.A(new_n265), .ZN(new_n384));
  OAI22_X1  g0184(.A1(new_n383), .A2(new_n384), .B1(new_n201), .B2(new_n258), .ZN(new_n385));
  INV_X1    g0185(.A(new_n335), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n385), .B1(new_n288), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n387), .A2(new_n297), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n290), .A2(G50), .ZN(new_n389));
  XOR2_X1   g0189(.A(new_n389), .B(KEYINPUT71), .Z(new_n390));
  OAI22_X1  g0190(.A1(new_n390), .A2(new_n298), .B1(G50), .B2(new_n296), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(new_n381), .B2(new_n316), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n382), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n366), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT9), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n392), .B(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n381), .A2(G200), .ZN(new_n398));
  OAI211_X1 g0198(.A(G190), .B(new_n368), .C1(new_n379), .C2(new_n380), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  OR2_X1    g0200(.A1(new_n400), .A2(KEYINPUT10), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(KEYINPUT10), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n335), .A2(new_n202), .B1(new_n258), .B2(G68), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT76), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n404), .A2(new_n405), .B1(new_n239), .B2(new_n384), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n404), .A2(new_n405), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n269), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT11), .ZN(new_n409));
  OR2_X1    g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n409), .ZN(new_n411));
  OR3_X1    g0211(.A1(new_n296), .A2(KEYINPUT12), .A3(G68), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT12), .B1(new_n296), .B2(G68), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n341), .A2(G68), .A3(new_n290), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n410), .A2(new_n411), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n231), .A2(G1698), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(G226), .B2(G1698), .ZN(new_n418));
  INV_X1    g0218(.A(G97), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n418), .A2(new_n257), .B1(new_n250), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n355), .B1(new_n420), .B2(new_n369), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT74), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n345), .B1(new_n307), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n422), .B2(new_n307), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT13), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT13), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n421), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT14), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(G169), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n361), .B2(new_n429), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n430), .B1(new_n429), .B2(G169), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n416), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n426), .A2(G190), .A3(new_n428), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT75), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n435), .B(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n416), .B1(new_n429), .B2(G200), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  AND4_X1   g0241(.A1(new_n333), .A2(new_n395), .A3(new_n403), .A4(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n305), .A2(G274), .ZN(new_n443));
  INV_X1    g0243(.A(G45), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(G1), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT5), .B(G41), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G257), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(new_n445), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n305), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n447), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT81), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n253), .A2(new_n346), .ZN(new_n453));
  INV_X1    g0253(.A(G244), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT4), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT4), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n452), .B(new_n457), .C1(new_n453), .C2(new_n454), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n257), .A2(new_n346), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n459), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n456), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n369), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT82), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT82), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n461), .A2(new_n464), .A3(new_n369), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n451), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n451), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n466), .A2(new_n361), .B1(new_n316), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n349), .A2(KEYINPUT6), .A3(G97), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n470), .A2(KEYINPUT79), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(KEYINPUT79), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n419), .A2(new_n349), .ZN(new_n473));
  NOR2_X1   g0273(.A1(G97), .A2(G107), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n471), .B(new_n472), .C1(new_n475), .C2(KEYINPUT6), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n476), .A2(G20), .B1(G77), .B2(new_n265), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n254), .A2(new_n259), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G107), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n297), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n296), .A2(G97), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n298), .B1(new_n289), .B2(G33), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n482), .B1(new_n483), .B2(G97), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT80), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n481), .A2(new_n486), .A3(new_n484), .ZN(new_n487));
  INV_X1    g0287(.A(new_n484), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT80), .B1(new_n488), .B2(new_n480), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n462), .A2(G190), .A3(new_n467), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n465), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n464), .B1(new_n461), .B2(new_n369), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n467), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G200), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n469), .A2(new_n485), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n253), .A2(new_n258), .A3(G87), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n497), .B(KEYINPUT22), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT24), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT23), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n258), .B2(G107), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n349), .A2(KEYINPUT23), .A3(G20), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n386), .A2(G116), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n498), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n499), .B1(new_n498), .B2(new_n503), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n269), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT25), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n296), .B2(G107), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n339), .A2(KEYINPUT25), .A3(new_n349), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n483), .A2(G107), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n448), .A2(G1698), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n253), .B(new_n512), .C1(G250), .C2(G1698), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G294), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n305), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n449), .A2(G264), .A3(new_n305), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(new_n447), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G169), .ZN(new_n519));
  OR2_X1    g0319(.A1(new_n517), .A2(KEYINPUT83), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n517), .A2(KEYINPUT83), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n515), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n447), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n519), .B1(new_n523), .B2(new_n361), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n511), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n525), .A2(KEYINPUT84), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT84), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n527), .B1(new_n511), .B2(new_n524), .ZN(new_n528));
  AOI21_X1  g0328(.A(G200), .B1(new_n522), .B2(new_n447), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n518), .A2(G190), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n506), .B(new_n510), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n526), .A2(new_n528), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(G270), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n447), .B1(new_n534), .B2(new_n450), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n459), .A2(G264), .B1(G303), .B2(new_n257), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n448), .B2(new_n453), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n535), .B1(new_n537), .B2(new_n369), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(new_n316), .ZN(new_n539));
  AOI21_X1  g0339(.A(G20), .B1(G33), .B2(G283), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(G33), .B2(new_n419), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n541), .B(new_n269), .C1(new_n258), .C2(G116), .ZN(new_n542));
  XOR2_X1   g0342(.A(new_n542), .B(KEYINPUT20), .Z(new_n543));
  NAND2_X1  g0343(.A1(new_n483), .A2(G116), .ZN(new_n544));
  INV_X1    g0344(.A(G116), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n339), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT21), .B1(new_n539), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n547), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n538), .A2(G190), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n550), .B(new_n551), .C1(new_n323), .C2(new_n538), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n547), .A2(G179), .A3(new_n538), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n539), .A2(new_n547), .A3(KEYINPUT21), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n549), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n253), .A2(new_n258), .A3(G68), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n335), .A2(new_n419), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n250), .A2(new_n419), .ZN(new_n558));
  AOI21_X1  g0358(.A(G20), .B1(new_n558), .B2(KEYINPUT19), .ZN(new_n559));
  NOR3_X1   g0359(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n560));
  OAI221_X1 g0360(.A(new_n556), .B1(KEYINPUT19), .B2(new_n557), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n561), .A2(new_n269), .B1(new_n339), .B2(new_n337), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n483), .A2(G87), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n443), .A2(new_n445), .ZN(new_n565));
  INV_X1    g0365(.A(new_n445), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n566), .A2(G250), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n305), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G116), .ZN(new_n570));
  OAI221_X1 g0370(.A(new_n570), .B1(new_n453), .B2(new_n345), .C1(new_n454), .C2(new_n370), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n569), .B1(new_n571), .B2(new_n369), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n564), .B1(G190), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n323), .B2(new_n572), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n483), .A2(new_n336), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n572), .A2(new_n361), .B1(new_n562), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(G169), .B2(new_n572), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n555), .A2(new_n578), .ZN(new_n579));
  AND4_X1   g0379(.A1(new_n442), .A2(new_n496), .A3(new_n533), .A4(new_n579), .ZN(G372));
  INV_X1    g0380(.A(KEYINPUT85), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n571), .A2(new_n581), .A3(new_n369), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n581), .B1(new_n571), .B2(new_n369), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n565), .B(new_n568), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n316), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n576), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(G200), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n573), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n587), .A2(new_n589), .A3(new_n531), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n496), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n525), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n554), .A2(new_n553), .ZN(new_n593));
  OAI21_X1  g0393(.A(KEYINPUT86), .B1(new_n593), .B2(new_n548), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT86), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n549), .A2(new_n595), .A3(new_n553), .A4(new_n554), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n592), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n469), .A2(new_n485), .A3(new_n577), .A4(new_n574), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT26), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n576), .A2(new_n586), .B1(new_n588), .B2(new_n573), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT26), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n487), .A2(new_n489), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n469), .A4(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n600), .A2(new_n604), .A3(new_n587), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n598), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n442), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g0408(.A(new_n608), .B(KEYINPUT87), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT89), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n439), .A2(new_n362), .A3(new_n363), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n434), .ZN(new_n612));
  INV_X1    g0412(.A(new_n332), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n322), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT88), .ZN(new_n616));
  INV_X1    g0416(.A(new_n402), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n400), .A2(KEYINPUT10), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n401), .A2(KEYINPUT88), .A3(new_n402), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n614), .A2(new_n615), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n394), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n610), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n619), .A2(new_n620), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n322), .B1(new_n612), .B2(new_n613), .ZN(new_n626));
  OAI211_X1 g0426(.A(KEYINPUT89), .B(new_n394), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n609), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  XNOR2_X1  g0428(.A(new_n628), .B(KEYINPUT90), .ZN(G369));
  NAND3_X1  g0429(.A1(new_n289), .A2(new_n258), .A3(G13), .ZN(new_n630));
  OR2_X1    g0430(.A1(new_n630), .A2(KEYINPUT27), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(KEYINPUT27), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(G213), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(G343), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n550), .A2(new_n636), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n555), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n594), .A2(new_n596), .A3(new_n637), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(G330), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n511), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n533), .B1(new_n643), .B2(new_n636), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n644), .B1(new_n525), .B2(new_n636), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n549), .A2(new_n553), .A3(new_n554), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n636), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n533), .A2(new_n649), .B1(new_n592), .B2(new_n636), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n646), .A2(new_n650), .ZN(G399));
  INV_X1    g0451(.A(new_n221), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(G41), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n560), .A2(new_n545), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n653), .A2(new_n654), .A3(new_n289), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n217), .B2(new_n653), .ZN(new_n656));
  XOR2_X1   g0456(.A(new_n656), .B(KEYINPUT28), .Z(new_n657));
  INV_X1    g0457(.A(KEYINPUT29), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n526), .A2(new_n528), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n496), .B(new_n590), .C1(new_n659), .C2(new_n647), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT93), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n599), .A2(new_n661), .A3(new_n602), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n601), .A2(new_n469), .A3(new_n603), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n662), .B1(new_n602), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n661), .B1(new_n599), .B2(new_n602), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n660), .B(new_n587), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n658), .B1(new_n666), .B2(new_n636), .ZN(new_n667));
  INV_X1    g0467(.A(G330), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT91), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n538), .A2(new_n522), .A3(new_n572), .A4(G179), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n669), .B1(new_n670), .B2(new_n468), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT30), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n538), .A2(G179), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n494), .A2(new_n523), .A3(new_n585), .A4(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT30), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n669), .B(new_n675), .C1(new_n670), .C2(new_n468), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n672), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n635), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT31), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT92), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n533), .A2(new_n579), .A3(new_n496), .A4(new_n636), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n677), .A2(KEYINPUT31), .A3(new_n635), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT92), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n668), .B1(new_n684), .B2(new_n687), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n606), .A2(KEYINPUT29), .A3(new_n635), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n667), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n657), .B1(new_n690), .B2(G1), .ZN(G364));
  AND2_X1   g0491(.A1(new_n258), .A2(G13), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n289), .B1(new_n692), .B2(G45), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(new_n653), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(G13), .A2(G33), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G20), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT94), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n638), .A2(new_n639), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n218), .B1(G20), .B2(new_n316), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n270), .A2(new_n272), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n221), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(new_n444), .B2(new_n217), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n444), .B2(new_n245), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n652), .A2(new_n257), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n711), .A2(G355), .B1(new_n545), .B2(new_n652), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n705), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n325), .A2(G179), .A3(G200), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(new_n258), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G97), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n258), .A2(new_n361), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G200), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G190), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n719), .A2(new_n325), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI221_X1 g0523(.A(new_n717), .B1(new_n721), .B2(new_n241), .C1(new_n239), .C2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT95), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(new_n258), .B2(G190), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n323), .A2(G179), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n325), .A2(KEYINPUT95), .A3(G20), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n349), .ZN(new_n730));
  INV_X1    g0530(.A(new_n718), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n731), .A2(new_n325), .A3(G200), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n253), .B1(new_n733), .B2(new_n261), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n727), .A2(G20), .A3(G190), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G87), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n731), .A2(G190), .A3(G200), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n737), .B1(new_n739), .B2(new_n202), .ZN(new_n740));
  OR4_X1    g0540(.A1(new_n724), .A2(new_n730), .A3(new_n734), .A4(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G179), .A2(G200), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n726), .A2(new_n728), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G159), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g0545(.A(KEYINPUT96), .B(KEYINPUT32), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n745), .B(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(G322), .ZN(new_n748));
  INV_X1    g0548(.A(G311), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n733), .A2(new_n748), .B1(new_n739), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n750), .B1(G294), .B2(new_n716), .ZN(new_n751));
  XNOR2_X1  g0551(.A(KEYINPUT33), .B(G317), .ZN(new_n752));
  AOI22_X1  g0552(.A1(G326), .A2(new_n722), .B1(new_n720), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n729), .ZN(new_n754));
  INV_X1    g0554(.A(new_n743), .ZN(new_n755));
  AOI22_X1  g0555(.A1(G283), .A2(new_n754), .B1(new_n755), .B2(G329), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n751), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G303), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n257), .B1(new_n735), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT97), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n741), .A2(new_n747), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n713), .B1(new_n761), .B2(new_n703), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n696), .B1(new_n702), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n640), .B(G330), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n763), .B1(new_n764), .B2(new_n696), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT98), .ZN(G396));
  NAND2_X1  g0566(.A1(new_n343), .A2(new_n635), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n360), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n364), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n362), .A2(new_n363), .A3(new_n636), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(new_n606), .B2(new_n635), .ZN(new_n772));
  INV_X1    g0572(.A(new_n771), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n636), .B(new_n773), .C1(new_n598), .C2(new_n605), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n688), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n695), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n688), .A2(new_n772), .A3(new_n774), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n703), .A2(new_n697), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n696), .B1(new_n202), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n717), .B1(new_n723), .B2(new_n758), .ZN(new_n781));
  INV_X1    g0581(.A(G294), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n733), .A2(new_n782), .B1(new_n349), .B2(new_n735), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n253), .B(new_n783), .C1(G116), .C2(new_n738), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n754), .A2(G87), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n784), .B(new_n785), .C1(new_n749), .C2(new_n743), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n781), .B(new_n786), .C1(G283), .C2(new_n720), .ZN(new_n787));
  XNOR2_X1  g0587(.A(KEYINPUT100), .B(G143), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n733), .A2(new_n788), .B1(new_n739), .B2(new_n744), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G137), .A2(new_n722), .B1(new_n720), .B2(G150), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(KEYINPUT99), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n790), .A2(KEYINPUT99), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n789), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(KEYINPUT34), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(KEYINPUT34), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n707), .B1(G50), .B2(new_n736), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n729), .A2(new_n241), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(G132), .B2(new_n755), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n797), .B(new_n799), .C1(new_n261), .C2(new_n715), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n787), .B1(new_n795), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n703), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n780), .B1(new_n802), .B2(new_n803), .C1(new_n773), .C2(new_n698), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n778), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G384));
  INV_X1    g0606(.A(KEYINPUT38), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT102), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n275), .A2(new_n276), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G68), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n297), .B1(new_n810), .B2(new_n278), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n247), .B1(new_n277), .B2(new_n267), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n299), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n808), .B1(new_n813), .B2(new_n633), .ZN(new_n814));
  INV_X1    g0614(.A(new_n267), .ZN(new_n815));
  AOI21_X1  g0615(.A(KEYINPUT16), .B1(new_n810), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n269), .B1(new_n277), .B2(new_n279), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n300), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n633), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n818), .A2(KEYINPUT102), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(new_n317), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n814), .A2(new_n820), .A3(new_n328), .A4(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT103), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n822), .A2(new_n823), .A3(KEYINPUT37), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n814), .A2(new_n820), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n322), .B2(new_n332), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n301), .A2(new_n819), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT37), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n318), .A2(new_n828), .A3(new_n829), .A4(new_n328), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT103), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(KEYINPUT37), .B2(new_n822), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n807), .B1(new_n827), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n822), .A2(KEYINPUT37), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n830), .A2(KEYINPUT103), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n836), .A2(KEYINPUT38), .A3(new_n824), .A4(new_n826), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n833), .A2(KEYINPUT104), .A3(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT104), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n839), .B(new_n807), .C1(new_n827), .C2(new_n832), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT105), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n333), .A2(new_n828), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n318), .A2(new_n828), .A3(new_n328), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(new_n829), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n807), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT39), .B1(new_n837), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n842), .A2(new_n843), .A3(new_n849), .ZN(new_n850));
  OR2_X1    g0650(.A1(new_n434), .A2(new_n635), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT39), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n838), .B2(new_n840), .ZN(new_n854));
  OAI21_X1  g0654(.A(KEYINPUT105), .B1(new_n854), .B2(new_n848), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n850), .A2(new_n852), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n440), .A2(new_n416), .A3(new_n635), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n416), .A2(new_n635), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n434), .A2(new_n439), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n774), .B2(new_n770), .ZN(new_n862));
  INV_X1    g0662(.A(new_n841), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n862), .A2(new_n863), .B1(new_n322), .B2(new_n633), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n856), .A2(KEYINPUT106), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT106), .B1(new_n856), .B2(new_n864), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n442), .B1(new_n667), .B2(new_n689), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n623), .A2(new_n627), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT107), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n867), .B(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n683), .A2(new_n680), .A3(new_n685), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n771), .B1(new_n857), .B2(new_n859), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT40), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(new_n840), .A4(new_n838), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n837), .A2(new_n847), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT40), .B1(new_n880), .B2(new_n875), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n442), .A2(new_n873), .ZN(new_n884));
  OAI21_X1  g0684(.A(G330), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n884), .B2(new_n883), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n872), .A2(new_n886), .B1(new_n289), .B2(new_n692), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n872), .B2(new_n886), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n218), .A2(new_n258), .A3(new_n545), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n476), .B(KEYINPUT101), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT35), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n892), .B2(new_n891), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT36), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n217), .B(G77), .C1(new_n261), .C2(new_n241), .ZN(new_n896));
  AOI211_X1 g0696(.A(new_n289), .B(G13), .C1(new_n896), .C2(new_n240), .ZN(new_n897));
  OR3_X1    g0697(.A1(new_n888), .A2(new_n895), .A3(new_n897), .ZN(G367));
  AOI21_X1  g0698(.A(new_n636), .B1(new_n562), .B2(new_n563), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n601), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n587), .B2(new_n900), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n902), .A2(new_n700), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n704), .B1(new_n221), .B2(new_n337), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n229), .A2(new_n708), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n695), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT112), .Z(new_n907));
  OAI22_X1  g0707(.A1(new_n733), .A2(new_n383), .B1(new_n739), .B2(new_n239), .ZN(new_n908));
  AOI211_X1 g0708(.A(new_n257), .B(new_n908), .C1(G58), .C2(new_n736), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n715), .A2(new_n241), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n723), .A2(new_n788), .ZN(new_n911));
  AOI211_X1 g0711(.A(new_n910), .B(new_n911), .C1(G159), .C2(new_n720), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n729), .A2(new_n202), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n755), .A2(G137), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n909), .A2(new_n912), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n736), .A2(KEYINPUT46), .A3(G116), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT46), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n735), .B2(new_n545), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n917), .B(new_n919), .C1(new_n721), .C2(new_n782), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT113), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(G283), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n733), .A2(new_n758), .B1(new_n739), .B2(new_n923), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n723), .A2(new_n749), .B1(new_n349), .B2(new_n715), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n924), .A2(new_n706), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n920), .A2(new_n921), .ZN(new_n927));
  AOI22_X1  g0727(.A1(G97), .A2(new_n754), .B1(new_n755), .B2(G317), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n916), .B1(new_n922), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT47), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n803), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n907), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n903), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n496), .B1(new_n603), .B2(new_n635), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n636), .B(new_n469), .C1(new_n489), .C2(new_n487), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT108), .ZN(new_n939));
  INV_X1    g0739(.A(new_n646), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT109), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n902), .A2(KEYINPUT43), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n941), .A2(new_n942), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n943), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n945), .B1(new_n943), .B2(new_n946), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n938), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n649), .A2(new_n533), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT42), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n939), .A2(new_n659), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n469), .A2(new_n485), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n635), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(KEYINPUT43), .B2(new_n902), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n949), .B(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT110), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT44), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n650), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n950), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n961), .A2(new_n962), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n938), .A2(new_n650), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT45), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n966), .A2(new_n940), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n940), .B1(new_n966), .B2(new_n968), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n951), .A2(KEYINPUT111), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n645), .A2(new_n649), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n951), .A2(KEYINPUT111), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(new_n642), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n690), .B1(new_n971), .B2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n653), .B(KEYINPUT41), .Z(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n694), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n935), .B1(new_n960), .B2(new_n980), .ZN(G387));
  XNOR2_X1  g0781(.A(new_n975), .B(new_n641), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n645), .A2(new_n700), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n711), .A2(new_n654), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(G107), .B2(new_n221), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n708), .B1(new_n234), .B2(G45), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n444), .B1(new_n241), .B2(new_n202), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(new_n654), .B2(KEYINPUT114), .ZN(new_n988));
  AND3_X1   g0788(.A1(new_n284), .A2(KEYINPUT50), .A3(new_n239), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT50), .B1(new_n284), .B2(new_n239), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n988), .B1(KEYINPUT114), .B2(new_n654), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n985), .B1(new_n986), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n695), .B1(new_n992), .B2(new_n705), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT115), .Z(new_n994));
  AOI21_X1  g0794(.A(new_n707), .B1(G77), .B2(new_n736), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n419), .B2(new_n729), .C1(new_n383), .C2(new_n743), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT116), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n288), .A2(new_n720), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n337), .A2(new_n715), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n733), .A2(new_n239), .B1(new_n739), .B2(new_n241), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(G159), .C2(new_n722), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n997), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n706), .B1(G326), .B2(new_n755), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n715), .A2(new_n923), .B1(new_n735), .B2(new_n782), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G303), .A2(new_n738), .B1(new_n732), .B2(G317), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n749), .B2(new_n721), .C1(new_n748), .C2(new_n723), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT48), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n1007), .B2(new_n1006), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT49), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1003), .B1(new_n545), .B2(new_n729), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1002), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n994), .B1(new_n703), .B2(new_n1013), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n982), .A2(new_n694), .B1(new_n983), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n690), .ZN(new_n1016));
  OAI211_X1 g0816(.A(KEYINPUT117), .B(new_n653), .C1(new_n976), .C2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n976), .A2(new_n1016), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n982), .A2(new_n690), .ZN(new_n1020));
  AOI21_X1  g0820(.A(KEYINPUT117), .B1(new_n1020), .B2(new_n653), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1015), .B1(new_n1019), .B2(new_n1021), .ZN(G393));
  NAND3_X1  g0822(.A1(new_n969), .A2(new_n694), .A3(new_n970), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n704), .B1(new_n419), .B2(new_n221), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n708), .A2(new_n238), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n695), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n732), .A2(G159), .B1(new_n722), .B2(G150), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT51), .Z(new_n1028));
  NOR2_X1   g0828(.A1(new_n735), .A2(new_n241), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1029), .B(new_n707), .C1(new_n284), .C2(new_n738), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n715), .A2(new_n202), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G50), .B2(new_n720), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n785), .B1(new_n743), .B2(new_n788), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1028), .A2(new_n1030), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n732), .A2(G311), .B1(new_n722), .B2(G317), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT52), .Z(new_n1037));
  AOI211_X1 g0837(.A(new_n253), .B(new_n730), .C1(G283), .C2(new_n736), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1037), .B(new_n1038), .C1(new_n748), .C2(new_n743), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G294), .A2(new_n738), .B1(new_n716), .B2(G116), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n758), .B2(new_n721), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT118), .Z(new_n1042));
  OAI21_X1  g0842(.A(new_n1035), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1026), .B1(new_n1043), .B2(new_n703), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n939), .B2(new_n700), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1023), .A2(new_n1045), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n971), .A2(new_n1020), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n653), .B1(new_n971), .B2(new_n1020), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1046), .B1(new_n1047), .B2(new_n1048), .ZN(G390));
  AOI21_X1  g0849(.A(new_n843), .B1(new_n842), .B2(new_n849), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n854), .A2(KEYINPUT105), .A3(new_n848), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1050), .A2(new_n1051), .B1(new_n852), .B2(new_n862), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n666), .A2(new_n636), .A3(new_n769), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n1053), .A2(new_n770), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n851), .B(new_n879), .C1(new_n1054), .C2(new_n861), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n688), .A2(new_n773), .A3(new_n860), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1052), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n873), .A2(G330), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n1058), .A2(new_n771), .A3(new_n861), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n862), .A2(new_n852), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n850), .B2(new_n855), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n861), .B1(new_n1053), .B2(new_n770), .ZN(new_n1062));
  NOR3_X1   g0862(.A1(new_n1062), .A2(new_n852), .A3(new_n880), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1059), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1057), .A2(new_n1064), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n873), .A2(G330), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n442), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n868), .A2(new_n869), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n774), .A2(new_n770), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n860), .B1(new_n688), .B2(new_n773), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1069), .B1(new_n1070), .B2(new_n1059), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n861), .B1(new_n1058), .B2(new_n771), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1054), .A2(new_n1056), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1068), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1065), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1057), .A2(new_n1064), .A3(new_n1074), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1076), .A2(new_n653), .A3(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1057), .A2(new_n1064), .A3(new_n694), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n779), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G97), .A2(new_n738), .B1(new_n732), .B2(G116), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(new_n257), .A3(new_n737), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n798), .B(new_n1082), .C1(G294), .C2(new_n755), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n723), .A2(new_n923), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1031), .B(new_n1084), .C1(G107), .C2(new_n720), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n722), .A2(G128), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n744), .B2(new_n715), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n736), .A2(G150), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1087), .B1(KEYINPUT53), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n257), .B1(new_n732), .B2(G132), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(KEYINPUT54), .B(G143), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1090), .B1(new_n739), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(G137), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n721), .A2(new_n1093), .B1(new_n1088), .B2(KEYINPUT53), .ZN(new_n1094));
  INV_X1    g0894(.A(G125), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n239), .A2(new_n729), .B1(new_n743), .B2(new_n1095), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n1092), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1083), .A2(new_n1085), .B1(new_n1089), .B2(new_n1097), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n695), .B1(new_n288), .B2(new_n1080), .C1(new_n1098), .C2(new_n803), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n850), .A2(new_n855), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1099), .B1(new_n1100), .B2(new_n697), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT119), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1078), .A2(new_n1079), .A3(new_n1102), .ZN(G378));
  INV_X1    g0903(.A(KEYINPUT57), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1068), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1077), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n856), .A2(new_n864), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT106), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n856), .A2(KEYINPUT106), .A3(new_n864), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n624), .A2(new_n394), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n392), .A2(new_n633), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n624), .B(new_n394), .C1(new_n392), .C2(new_n633), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1113), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1120), .A2(G330), .A3(new_n882), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n882), .A2(G330), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1109), .A2(new_n1110), .A3(new_n1121), .A4(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1121), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n865), .B2(new_n866), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1104), .B1(new_n1106), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT121), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1077), .A2(new_n1105), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1132), .A2(KEYINPUT57), .A3(new_n1125), .A4(new_n1127), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n1133), .A2(new_n653), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1132), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1135), .A2(KEYINPUT121), .A3(new_n1104), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1131), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1125), .A2(new_n1127), .A3(new_n694), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n696), .B1(new_n239), .B2(new_n779), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n707), .A2(new_n304), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(G77), .B2(new_n736), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n754), .A2(G58), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(new_n923), .C2(new_n743), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT120), .Z(new_n1144));
  OAI22_X1  g0944(.A1(new_n349), .A2(new_n733), .B1(new_n739), .B2(new_n337), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n721), .A2(new_n419), .B1(new_n723), .B2(new_n545), .ZN(new_n1146));
  OR4_X1    g0946(.A1(new_n910), .A2(new_n1144), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT58), .ZN(new_n1148));
  OR2_X1    g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1091), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n732), .A2(G128), .B1(new_n736), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n1093), .B2(new_n739), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G150), .A2(new_n716), .B1(new_n720), .B2(G132), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1153), .B(new_n1154), .C1(new_n1095), .C2(new_n723), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1155), .A2(KEYINPUT59), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(G33), .A2(G41), .ZN(new_n1157));
  INV_X1    g0957(.A(G124), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1157), .B1(new_n729), .B2(new_n744), .C1(new_n1158), .C2(new_n743), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n1155), .B2(KEYINPUT59), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1157), .A2(G50), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1156), .A2(new_n1160), .B1(new_n1140), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1149), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n1148), .B2(new_n1147), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1139), .B1(new_n803), .B2(new_n1164), .C1(new_n1120), .C2(new_n698), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1138), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1137), .A2(new_n1166), .ZN(G375));
  AOI22_X1  g0967(.A1(new_n732), .A2(G283), .B1(G97), .B2(new_n736), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1168), .B(new_n257), .C1(new_n349), .C2(new_n739), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n913), .B(new_n1169), .C1(G303), .C2(new_n755), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n721), .A2(new_n545), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n999), .B(new_n1171), .C1(G294), .C2(new_n722), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n721), .A2(new_n1091), .B1(new_n239), .B2(new_n715), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n707), .B(new_n1173), .C1(G132), .C2(new_n722), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n738), .A2(G150), .B1(G159), .B2(new_n736), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1175), .B(new_n1142), .C1(new_n1093), .C2(new_n733), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G128), .B2(new_n755), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1170), .A2(new_n1172), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n695), .B1(G68), .B2(new_n1080), .C1(new_n1178), .C2(new_n803), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n861), .B2(new_n697), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n693), .B(KEYINPUT122), .Z(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1180), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1075), .A2(new_n979), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1181), .A2(new_n1105), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(G381));
  AOI21_X1  g0987(.A(G378), .B1(G375), .B2(KEYINPUT124), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(KEYINPUT124), .B2(G375), .ZN(new_n1189));
  INV_X1    g0989(.A(G387), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1191));
  INV_X1    g0991(.A(G396), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1191), .A2(new_n1192), .A3(new_n1015), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(G390), .A2(G384), .A3(G381), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1190), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT123), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1189), .A2(new_n1197), .ZN(G407));
  NAND2_X1  g0998(.A1(new_n634), .A2(G213), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT125), .Z(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  OAI211_X1 g1001(.A(G407), .B(G213), .C1(new_n1189), .C2(new_n1201), .ZN(G409));
  INV_X1    g1002(.A(KEYINPUT61), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1137), .A2(G378), .A3(new_n1166), .ZN(new_n1204));
  INV_X1    g1004(.A(G378), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1135), .A2(new_n978), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1165), .B1(new_n1128), .B2(new_n1182), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1205), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1200), .B1(new_n1204), .B2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1075), .A2(new_n1186), .A3(KEYINPUT60), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n653), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1186), .B1(new_n1075), .B2(KEYINPUT60), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1184), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n805), .ZN(new_n1214));
  OAI211_X1 g1014(.A(G384), .B(new_n1184), .C1(new_n1211), .C2(new_n1212), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1214), .A2(new_n1215), .B1(G2897), .B2(new_n1200), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1199), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1219), .A2(G2897), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1216), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1203), .B1(new_n1209), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(KEYINPUT126), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1218), .A2(KEYINPUT62), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1209), .A2(new_n1224), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1219), .B(new_n1217), .C1(new_n1204), .C2(new_n1208), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1225), .B1(new_n1226), .B2(KEYINPUT62), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT126), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1228), .B(new_n1203), .C1(new_n1209), .C2(new_n1221), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1223), .A2(new_n1227), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(G393), .A2(G396), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1193), .A2(G390), .A3(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(G390), .B1(new_n1193), .B2(new_n1231), .ZN(new_n1234));
  OR3_X1    g1034(.A1(new_n1233), .A2(new_n1234), .A3(G387), .ZN(new_n1235));
  OAI21_X1  g1035(.A(G387), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1230), .A2(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1226), .A2(KEYINPUT63), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1219), .B1(new_n1204), .B2(new_n1208), .ZN(new_n1240));
  OR2_X1    g1040(.A1(new_n1240), .A2(new_n1221), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1209), .A2(KEYINPUT63), .A3(new_n1218), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1237), .A2(KEYINPUT61), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1239), .A2(new_n1241), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1238), .A2(new_n1244), .ZN(G405));
  AND3_X1   g1045(.A1(new_n1235), .A2(new_n1236), .A3(new_n1218), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1218), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1247));
  OAI21_X1  g1047(.A(KEYINPUT127), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1237), .A2(new_n1217), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT127), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1235), .A2(new_n1236), .A3(new_n1218), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1248), .A2(new_n1252), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(G375), .B(G378), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1253), .B(new_n1254), .ZN(G402));
endmodule


