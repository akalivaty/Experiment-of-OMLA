//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT2), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G113), .ZN(new_n193));
  INV_X1    g007(.A(G113), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(KEYINPUT2), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n189), .B(new_n191), .C1(new_n193), .C2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n189), .A2(new_n191), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT2), .B(G113), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n196), .A2(new_n199), .A3(KEYINPUT66), .ZN(new_n200));
  AOI21_X1  g014(.A(KEYINPUT66), .B1(new_n196), .B2(new_n199), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT11), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G137), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT11), .A3(G134), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n204), .A2(G137), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G131), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n205), .A2(new_n207), .A3(new_n212), .A4(new_n208), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n210), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n209), .A2(KEYINPUT65), .A3(G131), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT64), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n219), .A3(G143), .ZN(new_n220));
  AND2_X1   g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  INV_X1    g035(.A(G143), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G146), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n220), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n216), .A2(G143), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT64), .B(G146), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(G143), .ZN(new_n227));
  NOR2_X1   g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n221), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n214), .A2(new_n215), .A3(new_n224), .A4(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G128), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n220), .A2(new_n223), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n232), .B1(new_n220), .B2(KEYINPUT1), .ZN(new_n235));
  INV_X1    g049(.A(new_n225), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n217), .A2(new_n219), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n236), .B1(new_n237), .B2(new_n222), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n234), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n208), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n204), .A2(G137), .ZN(new_n241));
  OAI21_X1  g055(.A(G131), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n242), .A2(new_n213), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT30), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n231), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n245), .B1(new_n231), .B2(new_n244), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n202), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT31), .ZN(new_n249));
  NOR2_X1   g063(.A1(G237), .A2(G953), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G210), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n251), .B(KEYINPUT27), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(G101), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n252), .B(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n196), .A2(new_n199), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT66), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n196), .A2(new_n199), .A3(KEYINPUT66), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n231), .A2(new_n244), .A3(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n248), .A2(new_n249), .A3(new_n254), .A4(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n254), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT28), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n231), .A2(new_n244), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n202), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n264), .B1(new_n266), .B2(new_n260), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n260), .A2(new_n264), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n263), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n249), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n248), .A2(new_n254), .A3(new_n260), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n262), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(G472), .A2(G902), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n187), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n231), .A2(new_n244), .A3(new_n259), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n259), .B1(new_n231), .B2(new_n244), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT28), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n254), .B1(new_n279), .B2(new_n268), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n272), .B1(new_n280), .B2(KEYINPUT31), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n261), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(KEYINPUT32), .A3(new_n274), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n276), .A2(KEYINPUT67), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n275), .B1(new_n281), .B2(new_n261), .ZN(new_n285));
  OR3_X1    g099(.A1(new_n285), .A2(KEYINPUT67), .A3(KEYINPUT32), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n279), .A2(new_n254), .A3(new_n268), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT29), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n248), .A2(new_n260), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n289), .B1(new_n263), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n292), .B1(new_n287), .B2(new_n288), .ZN(new_n293));
  OAI21_X1  g107(.A(G472), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT68), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g110(.A(KEYINPUT68), .B(G472), .C1(new_n291), .C2(new_n293), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n284), .A2(new_n286), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  XOR2_X1   g112(.A(KEYINPUT69), .B(G217), .Z(new_n299));
  INV_X1    g113(.A(G234), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n299), .B1(new_n300), .B2(G902), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT77), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n292), .B1(new_n302), .B2(KEYINPUT25), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G140), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G125), .ZN(new_n306));
  INV_X1    g120(.A(G125), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G140), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT16), .ZN(new_n309));
  OR3_X1    g123(.A1(new_n307), .A2(KEYINPUT16), .A3(G140), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n216), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n310), .A3(G146), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n188), .A2(G128), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n232), .A2(G119), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT24), .B(G110), .ZN(new_n318));
  OR2_X1    g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G110), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT23), .B1(new_n232), .B2(G119), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT71), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI211_X1 g138(.A(KEYINPUT71), .B(KEYINPUT23), .C1(new_n232), .C2(G119), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n316), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(KEYINPUT23), .A2(G119), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT70), .B1(new_n327), .B2(G128), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT70), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n329), .A2(new_n232), .A3(KEYINPUT23), .A4(G119), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n321), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT72), .B1(new_n320), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n332), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT72), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n334), .A2(new_n335), .A3(new_n314), .A4(new_n319), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G953), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(G221), .A3(G234), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(KEYINPUT76), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT22), .B(G137), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n340), .B(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n325), .A2(new_n316), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT71), .B1(new_n315), .B2(KEYINPUT23), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n331), .B(new_n321), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT73), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT73), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n326), .A2(new_n347), .A3(new_n321), .A4(new_n331), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT74), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT74), .B1(new_n317), .B2(new_n318), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n349), .A2(KEYINPUT75), .A3(new_n353), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n306), .A2(new_n308), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n226), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n313), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n352), .B1(new_n346), .B2(new_n348), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(KEYINPUT75), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n337), .B(new_n342), .C1(new_n359), .C2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n349), .A2(new_n353), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT75), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n357), .B1(new_n360), .B2(KEYINPUT75), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n342), .B1(new_n368), .B2(new_n337), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n304), .B1(new_n363), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n302), .A2(KEYINPUT25), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n337), .B1(new_n359), .B2(new_n361), .ZN(new_n373));
  INV_X1    g187(.A(new_n342), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n362), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n376), .A2(new_n302), .A3(KEYINPUT25), .A4(new_n292), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n301), .B1(new_n372), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n301), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(G902), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT78), .B1(new_n378), .B2(new_n382), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n376), .A2(new_n304), .B1(new_n302), .B2(KEYINPUT25), .ZN(new_n384));
  AOI211_X1 g198(.A(new_n303), .B(new_n371), .C1(new_n375), .C2(new_n362), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n379), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT78), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(new_n381), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(G234), .A2(G237), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(G952), .A3(new_n338), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(KEYINPUT91), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n390), .A2(G902), .A3(G953), .ZN(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT21), .B(G898), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(G214), .B1(G237), .B2(G902), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(G210), .B1(G237), .B2(G902), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n230), .A2(new_n224), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G125), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT1), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(new_n226), .B2(G143), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n227), .B1(new_n404), .B2(new_n232), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(new_n307), .A3(new_n234), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n338), .A2(G224), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n407), .B(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G104), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT3), .B1(new_n410), .B2(G107), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT80), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT80), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n413), .B(KEYINPUT3), .C1(new_n410), .C2(G107), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT3), .ZN(new_n415));
  INV_X1    g229(.A(G107), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n416), .A3(G104), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n410), .A2(G107), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n412), .A2(new_n414), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G101), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n417), .A2(new_n418), .ZN(new_n421));
  INV_X1    g235(.A(G101), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n421), .A2(new_n422), .A3(new_n414), .A4(new_n412), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n420), .A2(KEYINPUT4), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n419), .A2(new_n425), .A3(G101), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n202), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n418), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n410), .A2(G107), .ZN(new_n429));
  OAI21_X1  g243(.A(G101), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n423), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n432));
  INV_X1    g246(.A(new_n189), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n194), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n197), .B2(new_n432), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n431), .A2(new_n196), .A3(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(G110), .B(G122), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n427), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  XOR2_X1   g252(.A(new_n437), .B(KEYINPUT84), .Z(new_n439));
  AOI21_X1  g253(.A(new_n439), .B1(new_n427), .B2(new_n436), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(KEYINPUT85), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n438), .A2(KEYINPUT6), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n427), .A2(new_n436), .ZN(new_n444));
  INV_X1    g258(.A(new_n439), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n442), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n409), .B1(new_n443), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(KEYINPUT86), .A2(KEYINPUT7), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n402), .A2(new_n406), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(KEYINPUT7), .A3(new_n408), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n408), .A2(KEYINPUT7), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n402), .A2(new_n406), .A3(new_n453), .A4(new_n450), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n427), .A2(new_n436), .A3(new_n437), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT5), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n434), .B1(new_n457), .B2(new_n197), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n196), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n431), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n437), .B(KEYINPUT8), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n435), .A2(new_n196), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n460), .B(new_n461), .C1(new_n431), .C2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n455), .A2(new_n456), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n292), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n400), .B1(new_n449), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n409), .ZN(new_n467));
  OAI22_X1  g281(.A1(new_n446), .A2(new_n447), .B1(new_n441), .B2(new_n456), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n440), .A2(new_n442), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n456), .A2(new_n463), .ZN(new_n471));
  AOI21_X1  g285(.A(G902), .B1(new_n471), .B2(new_n455), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(new_n399), .A3(new_n472), .ZN(new_n473));
  AOI211_X1 g287(.A(new_n396), .B(new_n398), .C1(new_n466), .C2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(G237), .ZN(new_n475));
  AND4_X1   g289(.A1(G143), .A2(new_n475), .A3(new_n338), .A4(G214), .ZN(new_n476));
  AOI21_X1  g290(.A(G143), .B1(new_n250), .B2(G214), .ZN(new_n477));
  OAI211_X1 g291(.A(KEYINPUT17), .B(G131), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n312), .A2(new_n313), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT88), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n312), .A2(new_n478), .A3(new_n481), .A4(new_n313), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n476), .A2(new_n477), .A3(G131), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n475), .A2(new_n338), .A3(G214), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n222), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n250), .A2(G143), .A3(G214), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n212), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT17), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n480), .A2(new_n482), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n356), .B1(new_n216), .B2(new_n355), .ZN(new_n492));
  NAND2_X1  g306(.A1(KEYINPUT18), .A2(G131), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n485), .A2(new_n486), .A3(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(KEYINPUT18), .B(G131), .C1(new_n476), .C2(new_n477), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  XOR2_X1   g310(.A(G113), .B(G122), .Z(new_n497));
  XOR2_X1   g311(.A(KEYINPUT87), .B(G104), .Z(new_n498));
  XOR2_X1   g312(.A(new_n497), .B(new_n498), .Z(new_n499));
  NAND3_X1  g313(.A1(new_n491), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT89), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT89), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n491), .A2(new_n502), .A3(new_n496), .A4(new_n499), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  XOR2_X1   g318(.A(new_n355), .B(KEYINPUT19), .Z(new_n505));
  OAI221_X1 g319(.A(new_n313), .B1(new_n487), .B2(new_n483), .C1(new_n505), .C2(new_n237), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n499), .B1(new_n506), .B2(new_n496), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT20), .ZN(new_n510));
  NOR2_X1   g324(.A1(G475), .A2(G902), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n507), .B1(new_n501), .B2(new_n503), .ZN(new_n513));
  INV_X1    g327(.A(new_n511), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT20), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n496), .ZN(new_n517));
  AOI22_X1  g331(.A1(KEYINPUT88), .A2(new_n479), .B1(new_n488), .B2(new_n489), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n517), .B1(new_n518), .B2(new_n482), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(new_n499), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n520), .B1(new_n503), .B2(new_n501), .ZN(new_n521));
  OAI21_X1  g335(.A(G475), .B1(new_n521), .B2(G902), .ZN(new_n522));
  INV_X1    g336(.A(G122), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G116), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n190), .A2(G122), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G107), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n524), .A2(new_n525), .A3(new_n416), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT13), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n232), .B2(G143), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n232), .A2(G143), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n222), .A2(G128), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(new_n530), .ZN(new_n535));
  OAI21_X1  g349(.A(G134), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n532), .A3(new_n204), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n529), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n534), .A2(new_n532), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G134), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n537), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n190), .A2(KEYINPUT14), .A3(G122), .ZN(new_n542));
  OAI211_X1 g356(.A(G107), .B(new_n542), .C1(new_n526), .C2(KEYINPUT14), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n528), .A3(new_n543), .ZN(new_n544));
  XOR2_X1   g358(.A(KEYINPUT9), .B(G234), .Z(new_n545));
  NAND3_X1  g359(.A1(new_n299), .A2(new_n545), .A3(new_n338), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n538), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT90), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n538), .A2(new_n544), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n546), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n538), .A2(new_n544), .A3(KEYINPUT90), .A4(new_n547), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n292), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT15), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n555), .B1(new_n556), .B2(G478), .ZN(new_n557));
  INV_X1    g371(.A(G478), .ZN(new_n558));
  AOI211_X1 g372(.A(KEYINPUT15), .B(new_n558), .C1(new_n554), .C2(new_n292), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n516), .A2(new_n522), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(G221), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(new_n545), .B2(new_n292), .ZN(new_n564));
  XOR2_X1   g378(.A(new_n564), .B(KEYINPUT79), .Z(new_n565));
  XNOR2_X1  g379(.A(G110), .B(G140), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n338), .A2(G227), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n234), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n220), .A2(new_n223), .B1(new_n571), .B2(G128), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n423), .B(new_n430), .C1(new_n570), .C2(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n573), .B1(new_n431), .B2(new_n239), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n214), .A2(new_n215), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT12), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n574), .A2(KEYINPUT12), .A3(new_n576), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT10), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n582), .B1(new_n405), .B2(new_n234), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n583), .A2(new_n431), .B1(new_n573), .B2(new_n582), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT81), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n214), .A2(new_n585), .A3(new_n215), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n585), .B1(new_n214), .B2(new_n215), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n230), .A2(new_n224), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n424), .A2(new_n589), .A3(new_n426), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n584), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n569), .B1(new_n581), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n431), .A2(KEYINPUT10), .A3(new_n239), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n573), .A2(new_n582), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n590), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n576), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(new_n591), .A3(new_n569), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT82), .B1(new_n592), .B2(new_n598), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n574), .A2(KEYINPUT12), .A3(new_n576), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT12), .B1(new_n574), .B2(new_n576), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OR2_X1    g416(.A1(new_n586), .A2(new_n587), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n595), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n568), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT82), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(new_n606), .A3(new_n597), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n599), .A2(new_n607), .A3(G469), .ZN(new_n608));
  INV_X1    g422(.A(G469), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(new_n292), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n575), .B1(new_n584), .B2(new_n590), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n568), .B1(new_n604), .B2(new_n611), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n591), .B(new_n569), .C1(new_n600), .C2(new_n601), .ZN(new_n613));
  AOI21_X1  g427(.A(G902), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n610), .B1(new_n614), .B2(new_n609), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n565), .B1(new_n608), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n474), .A2(new_n562), .A3(new_n616), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n298), .A2(new_n389), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(new_n422), .ZN(G3));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n554), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n620), .B1(new_n551), .B2(new_n546), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n548), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n621), .A2(G478), .A3(new_n292), .A4(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT92), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n555), .A2(new_n558), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n624), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT92), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n516), .A2(new_n522), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n474), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(G902), .B1(new_n281), .B2(new_n261), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n285), .B1(new_n633), .B2(G472), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n616), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n389), .A2(new_n631), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT34), .B(G104), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  AOI21_X1  g452(.A(new_n398), .B1(new_n466), .B2(new_n473), .ZN(new_n639));
  INV_X1    g453(.A(new_n396), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n389), .A2(new_n635), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n512), .A2(new_n515), .A3(KEYINPUT93), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT94), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n522), .A2(new_n644), .ZN(new_n645));
  OAI211_X1 g459(.A(KEYINPUT94), .B(G475), .C1(new_n521), .C2(G902), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n643), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(KEYINPUT93), .B1(new_n512), .B2(new_n515), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n647), .A2(new_n560), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT35), .B(G107), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  INV_X1    g466(.A(KEYINPUT95), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n342), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n373), .B(new_n654), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n655), .A2(new_n380), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n378), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(G472), .ZN(new_n658));
  OAI22_X1  g472(.A1(new_n632), .A2(new_n658), .B1(new_n273), .B2(new_n275), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n653), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n655), .A2(new_n380), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n386), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n634), .A2(new_n662), .A3(KEYINPUT95), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n617), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  NAND2_X1  g482(.A1(new_n662), .A2(new_n616), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n284), .A2(new_n286), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n296), .A2(new_n297), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT93), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n516), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n674), .A2(new_n643), .A3(new_n645), .A4(new_n646), .ZN(new_n675));
  INV_X1    g489(.A(G900), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n393), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n392), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n675), .A2(new_n560), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n672), .A2(new_n639), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G128), .ZN(G30));
  XOR2_X1   g495(.A(new_n678), .B(KEYINPUT39), .Z(new_n682));
  NAND2_X1  g496(.A1(new_n616), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT40), .Z(new_n684));
  NAND2_X1  g498(.A1(new_n290), .A2(new_n254), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n266), .A2(new_n263), .A3(new_n260), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n292), .ZN(new_n688));
  OAI21_X1  g502(.A(G472), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n670), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT38), .ZN(new_n691));
  INV_X1    g505(.A(new_n473), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n399), .B1(new_n470), .B2(new_n472), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n466), .A2(new_n473), .A3(KEYINPUT38), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n560), .B1(new_n516), .B2(new_n522), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n397), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n696), .A2(new_n698), .A3(new_n662), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n684), .A2(new_n690), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G143), .ZN(G45));
  AOI21_X1  g515(.A(new_n510), .B1(new_n509), .B2(new_n511), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n513), .A2(KEYINPUT20), .A3(new_n514), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n522), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n629), .A2(new_n627), .ZN(new_n705));
  INV_X1    g519(.A(new_n678), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n397), .B1(new_n692), .B2(new_n693), .ZN(new_n708));
  OAI21_X1  g522(.A(KEYINPUT96), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT96), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n630), .A2(new_n639), .A3(new_n710), .A4(new_n706), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n672), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT97), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT97), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n672), .A2(new_n715), .A3(new_n712), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  NAND2_X1  g532(.A1(new_n670), .A2(new_n671), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n383), .A2(new_n388), .ZN(new_n720));
  INV_X1    g534(.A(new_n631), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT99), .B1(new_n614), .B2(new_n609), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT98), .ZN(new_n723));
  OAI21_X1  g537(.A(G469), .B1(new_n614), .B2(new_n723), .ZN(new_n724));
  AOI211_X1 g538(.A(KEYINPUT98), .B(G902), .C1(new_n612), .C2(new_n613), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n722), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n569), .B1(new_n595), .B2(new_n603), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n602), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n569), .B1(new_n596), .B2(new_n591), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n292), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(KEYINPUT98), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n614), .A2(new_n723), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n731), .A2(KEYINPUT99), .A3(new_n732), .A4(G469), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n564), .B1(new_n726), .B2(new_n733), .ZN(new_n734));
  AND4_X1   g548(.A1(new_n719), .A2(new_n720), .A3(new_n721), .A4(new_n734), .ZN(new_n735));
  XOR2_X1   g549(.A(KEYINPUT41), .B(G113), .Z(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G15));
  INV_X1    g551(.A(KEYINPUT100), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n298), .A2(new_n389), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n649), .A2(new_n734), .A3(new_n474), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n649), .A2(new_n734), .A3(new_n474), .ZN(new_n742));
  NOR4_X1   g556(.A1(new_n742), .A2(new_n298), .A3(KEYINPUT100), .A4(new_n389), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G116), .ZN(G18));
  NOR2_X1   g559(.A1(new_n561), .A2(new_n396), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n734), .A2(new_n639), .A3(new_n662), .A4(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n298), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n188), .ZN(G21));
  AND3_X1   g563(.A1(new_n734), .A2(new_n474), .A3(new_n697), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n378), .A2(new_n382), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT101), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n634), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n386), .A2(new_n381), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT101), .B1(new_n754), .B2(new_n659), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n750), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G122), .ZN(G24));
  NAND2_X1  g572(.A1(new_n726), .A2(new_n733), .ZN(new_n759));
  INV_X1    g573(.A(new_n564), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n639), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n707), .A2(KEYINPUT102), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT102), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n630), .A2(new_n764), .A3(new_n706), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n657), .A2(new_n659), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n762), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G125), .ZN(G27));
  NAND2_X1  g583(.A1(new_n605), .A2(new_n597), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n609), .B1(new_n770), .B2(new_n292), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n730), .A2(G469), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n760), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n466), .A2(new_n473), .A3(new_n397), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n719), .A2(new_n720), .A3(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT42), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n763), .A2(new_n765), .A3(new_n777), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n276), .A2(new_n283), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n754), .B1(new_n671), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n766), .A2(new_n780), .A3(new_n775), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n776), .A2(new_n778), .B1(new_n781), .B2(KEYINPUT42), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G131), .ZN(G33));
  NAND3_X1  g597(.A1(new_n739), .A2(new_n679), .A3(new_n775), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G134), .ZN(G36));
  NAND3_X1  g599(.A1(new_n705), .A2(new_n516), .A3(new_n522), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT104), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n786), .A2(new_n787), .A3(KEYINPUT43), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT43), .B1(new_n786), .B2(new_n787), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(new_n659), .A3(new_n662), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT44), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n774), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n791), .A2(new_n792), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n610), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT45), .B1(new_n599), .B2(new_n607), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT45), .ZN(new_n799));
  OAI21_X1  g613(.A(G469), .B1(new_n770), .B2(new_n799), .ZN(new_n800));
  OAI211_X1 g614(.A(KEYINPUT46), .B(new_n797), .C1(new_n798), .C2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT103), .ZN(new_n802));
  INV_X1    g616(.A(new_n772), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n802), .B1(new_n801), .B2(new_n803), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n798), .A2(new_n800), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT46), .B1(new_n807), .B2(new_n797), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n805), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(new_n564), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n682), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n796), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(new_n206), .ZN(G39));
  INV_X1    g627(.A(KEYINPUT47), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n814), .B1(new_n809), .B2(new_n564), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n806), .A2(new_n808), .ZN(new_n816));
  OAI211_X1 g630(.A(KEYINPUT47), .B(new_n760), .C1(new_n816), .C2(new_n805), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n719), .A2(new_n720), .A3(new_n707), .A4(new_n774), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G140), .ZN(G42));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n822));
  NOR2_X1   g636(.A1(G952), .A2(G953), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n672), .A2(new_n715), .A3(new_n712), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n715), .B1(new_n672), .B2(new_n712), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n697), .A2(new_n639), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n662), .A2(new_n773), .A3(new_n678), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n690), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n680), .A2(new_n768), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n824), .B1(new_n827), .B2(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n680), .A2(new_n768), .A3(new_n831), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(new_n717), .A3(KEYINPUT52), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n739), .A2(new_n721), .A3(new_n734), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n746), .A2(new_n662), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n761), .A2(new_n838), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n719), .A2(new_n839), .B1(new_n750), .B2(new_n756), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n837), .B(new_n840), .C1(new_n741), .C2(new_n743), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n776), .A2(new_n778), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n781), .A2(KEYINPUT42), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT109), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n766), .A2(new_n767), .A3(new_n775), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT108), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n557), .A2(new_n559), .A3(new_n678), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n397), .A2(new_n466), .A3(new_n473), .A4(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n645), .A2(new_n646), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n849), .A2(new_n674), .A3(new_n643), .A4(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n847), .B1(new_n672), .B2(new_n852), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n298), .A2(new_n851), .A3(KEYINPUT108), .A4(new_n669), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n784), .B(new_n846), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n839), .A2(new_n719), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n837), .A2(new_n858), .A3(new_n757), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT109), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n744), .A2(new_n859), .A3(new_n782), .A4(new_n860), .ZN(new_n861));
  AND4_X1   g675(.A1(new_n836), .A2(new_n845), .A3(new_n857), .A4(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT106), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n863), .B1(new_n618), .B2(new_n636), .ZN(new_n864));
  INV_X1    g678(.A(new_n635), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n720), .A2(new_n721), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n719), .A2(new_n720), .ZN(new_n867));
  OAI211_X1 g681(.A(KEYINPUT106), .B(new_n866), .C1(new_n867), .C2(new_n617), .ZN(new_n868));
  INV_X1    g682(.A(new_n560), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n516), .A2(new_n522), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n642), .A2(new_n871), .B1(new_n664), .B2(new_n665), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n864), .A2(new_n868), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT107), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT107), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n864), .A2(new_n868), .A3(new_n872), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n841), .A2(new_n844), .A3(new_n855), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n836), .A3(new_n878), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n862), .A2(new_n877), .B1(new_n856), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g694(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n856), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n877), .A2(new_n836), .A3(new_n878), .A4(KEYINPUT53), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n880), .A2(new_n881), .B1(new_n884), .B2(KEYINPUT54), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n788), .A2(new_n789), .A3(new_n392), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n734), .A2(new_n398), .A3(new_n696), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n887), .A3(new_n756), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT111), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT50), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT111), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n886), .A2(new_n887), .A3(new_n891), .A4(new_n756), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT112), .B1(new_n888), .B2(new_n890), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n889), .A2(KEYINPUT112), .A3(new_n890), .A4(new_n892), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n734), .A2(new_n794), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n886), .A2(new_n898), .A3(new_n767), .ZN(new_n899));
  INV_X1    g713(.A(new_n690), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n389), .A2(new_n392), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n901), .A3(new_n898), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n704), .A2(new_n705), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n759), .A2(new_n565), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n815), .A2(new_n817), .A3(new_n905), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n886), .A2(new_n756), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n907), .A2(new_n794), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n904), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n897), .A2(new_n909), .A3(KEYINPUT51), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT113), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT113), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n897), .A2(new_n909), .A3(new_n912), .A4(KEYINPUT51), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT51), .B1(new_n897), .B2(new_n909), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n886), .A2(new_n898), .A3(new_n780), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT48), .Z(new_n917));
  NAND2_X1  g731(.A1(new_n338), .A2(G952), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n918), .B1(new_n907), .B2(new_n762), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n704), .A2(new_n705), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n919), .B1(new_n920), .B2(new_n902), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n915), .A2(new_n917), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n914), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n823), .B1(new_n885), .B2(new_n924), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n754), .A2(new_n398), .A3(new_n565), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT105), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT49), .B1(new_n726), .B2(new_n733), .ZN(new_n928));
  AOI211_X1 g742(.A(new_n786), .B(new_n928), .C1(new_n695), .C2(new_n694), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n726), .A2(new_n733), .A3(KEYINPUT49), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n927), .A2(new_n929), .A3(new_n900), .A4(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n822), .B1(new_n925), .B2(new_n932), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n845), .A2(new_n861), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n934), .A2(new_n877), .A3(new_n836), .A4(new_n857), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n935), .A2(new_n882), .A3(new_n881), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT54), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n882), .B2(new_n883), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n936), .A2(new_n923), .A3(new_n938), .ZN(new_n939));
  OAI211_X1 g753(.A(KEYINPUT114), .B(new_n931), .C1(new_n939), .C2(new_n823), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n933), .A2(new_n940), .ZN(G75));
  INV_X1    g755(.A(KEYINPUT116), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n338), .A2(G952), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(G210), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n880), .A2(new_n945), .A3(new_n292), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n468), .A2(new_n469), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(new_n467), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT55), .Z(new_n949));
  XNOR2_X1  g763(.A(KEYINPUT115), .B(KEYINPUT56), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n944), .B1(new_n946), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n949), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n935), .A2(new_n882), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n955), .A2(G210), .A3(G902), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT56), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n942), .B1(new_n953), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n949), .B1(new_n946), .B2(KEYINPUT56), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n943), .B1(new_n956), .B2(new_n951), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n960), .A2(KEYINPUT116), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n959), .A2(new_n962), .ZN(G51));
  NOR2_X1   g777(.A1(new_n880), .A2(new_n881), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n964), .A2(new_n936), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n610), .B(KEYINPUT57), .Z(new_n966));
  OAI22_X1  g780(.A1(new_n965), .A2(new_n966), .B1(new_n729), .B2(new_n728), .ZN(new_n967));
  OR3_X1    g781(.A1(new_n880), .A2(new_n292), .A3(new_n807), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n943), .B1(new_n967), .B2(new_n968), .ZN(G54));
  NOR2_X1   g783(.A1(new_n880), .A2(new_n292), .ZN(new_n970));
  NAND2_X1  g784(.A1(KEYINPUT58), .A2(G475), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT117), .Z(new_n972));
  AND3_X1   g786(.A1(new_n970), .A2(new_n509), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n509), .B1(new_n970), .B2(new_n972), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n973), .A2(new_n974), .A3(new_n943), .ZN(G60));
  AND2_X1   g789(.A1(new_n621), .A2(new_n623), .ZN(new_n976));
  INV_X1    g790(.A(new_n885), .ZN(new_n977));
  XNOR2_X1  g791(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n978));
  NAND2_X1  g792(.A1(G478), .A2(G902), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n976), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n976), .A2(new_n980), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n944), .B1(new_n965), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n981), .A2(new_n983), .ZN(G63));
  NAND2_X1  g798(.A1(G217), .A2(G902), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT60), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n986), .B1(new_n935), .B2(new_n882), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n655), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(KEYINPUT119), .A2(KEYINPUT61), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n943), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n991), .B1(new_n987), .B2(new_n376), .ZN(new_n992));
  OAI211_X1 g806(.A(KEYINPUT119), .B(KEYINPUT61), .C1(new_n989), .C2(new_n992), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n987), .A2(new_n376), .ZN(new_n994));
  NAND2_X1  g808(.A1(KEYINPUT119), .A2(KEYINPUT61), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n994), .A2(new_n995), .A3(new_n988), .A4(new_n991), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n993), .A2(new_n996), .ZN(G66));
  INV_X1    g811(.A(G224), .ZN(new_n998));
  OAI21_X1  g812(.A(G953), .B1(new_n394), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n841), .B1(new_n874), .B2(new_n876), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n999), .B1(new_n1000), .B2(G953), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n947), .B1(G898), .B2(new_n338), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT120), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1001), .B(new_n1003), .ZN(G69));
  NOR2_X1   g818(.A1(new_n246), .A2(new_n247), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n505), .B(KEYINPUT121), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1005), .B(new_n1006), .Z(new_n1007));
  AOI21_X1  g821(.A(new_n1007), .B1(G900), .B2(G953), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n782), .A2(new_n784), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT123), .Z(new_n1010));
  INV_X1    g824(.A(new_n811), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n780), .A2(new_n829), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n812), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n680), .A2(new_n768), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n827), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1010), .A2(new_n820), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1008), .B1(new_n1016), .B2(G953), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n338), .B1(G227), .B2(G900), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT124), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AND2_X1   g834(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  AOI211_X1 g835(.A(new_n774), .B(new_n683), .C1(new_n920), .C2(new_n870), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(new_n739), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  AOI211_X1 g838(.A(new_n1024), .B(new_n812), .C1(new_n818), .C2(new_n819), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1015), .A2(new_n700), .ZN(new_n1026));
  OR2_X1    g840(.A1(new_n1026), .A2(KEYINPUT62), .ZN(new_n1027));
  AND3_X1   g841(.A1(new_n1026), .A2(KEYINPUT122), .A3(KEYINPUT62), .ZN(new_n1028));
  AOI21_X1  g842(.A(KEYINPUT122), .B1(new_n1026), .B2(KEYINPUT62), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n1025), .B(new_n1027), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1030), .A2(new_n338), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1031), .A2(new_n1007), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1033), .ZN(new_n1034));
  AND3_X1   g848(.A1(new_n1021), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1034), .B1(new_n1021), .B2(new_n1032), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n1035), .A2(new_n1036), .ZN(G72));
  NAND2_X1  g851(.A1(G472), .A2(G902), .ZN(new_n1038));
  XOR2_X1   g852(.A(new_n1038), .B(KEYINPUT63), .Z(new_n1039));
  INV_X1    g853(.A(new_n1000), .ZN(new_n1040));
  OAI211_X1 g854(.A(KEYINPUT125), .B(new_n1039), .C1(new_n1030), .C2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1041), .A2(new_n686), .ZN(new_n1042));
  OR2_X1    g856(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1043));
  NAND4_X1  g857(.A1(new_n1043), .A2(new_n1000), .A3(new_n1027), .A4(new_n1025), .ZN(new_n1044));
  AOI21_X1  g858(.A(KEYINPUT125), .B1(new_n1044), .B2(new_n1039), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n1039), .B1(new_n1016), .B2(new_n1040), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n248), .A2(new_n263), .A3(new_n260), .ZN(new_n1048));
  XNOR2_X1  g862(.A(new_n1048), .B(KEYINPUT126), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n943), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g864(.A(KEYINPUT127), .ZN(new_n1051));
  AND3_X1   g865(.A1(new_n685), .A2(new_n1039), .A3(new_n1048), .ZN(new_n1052));
  AND3_X1   g866(.A1(new_n884), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1051), .B1(new_n884), .B2(new_n1052), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n1050), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g869(.A1(new_n1046), .A2(new_n1055), .ZN(G57));
endmodule


