//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011;
  INV_X1    g000(.A(KEYINPUT100), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(KEYINPUT16), .A3(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G8gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT97), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n205), .B(new_n207), .C1(new_n204), .C2(new_n203), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n206), .A2(KEYINPUT97), .ZN(new_n209));
  XOR2_X1   g008(.A(new_n208), .B(new_n209), .Z(new_n210));
  INV_X1    g009(.A(KEYINPUT98), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(G43gat), .B(G50gat), .Z(new_n213));
  OR2_X1    g012(.A1(new_n213), .A2(KEYINPUT94), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(KEYINPUT94), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(KEYINPUT15), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G29gat), .ZN(new_n217));
  INV_X1    g016(.A(G36gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n219), .B(KEYINPUT14), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT15), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT95), .ZN(new_n222));
  INV_X1    g021(.A(G50gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(G43gat), .ZN(new_n224));
  INV_X1    g023(.A(G43gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(G50gat), .ZN(new_n226));
  NOR3_X1   g025(.A1(new_n222), .A2(new_n223), .A3(G43gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n221), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G29gat), .A2(G36gat), .ZN(new_n229));
  XOR2_X1   g028(.A(new_n229), .B(KEYINPUT96), .Z(new_n230));
  NAND4_X1  g029(.A1(new_n216), .A2(new_n220), .A3(new_n228), .A4(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n220), .A2(new_n229), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n232), .A2(KEYINPUT15), .A3(new_n215), .A4(new_n214), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n208), .B(new_n209), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT98), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n212), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT99), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n237), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n236), .A2(KEYINPUT98), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n234), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n212), .A2(KEYINPUT99), .A3(new_n235), .A4(new_n237), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G229gat), .A2(G233gat), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n246), .B(KEYINPUT13), .Z(new_n247));
  NAND2_X1  g046(.A1(new_n235), .A2(KEYINPUT17), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT17), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n210), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(new_n243), .A3(new_n246), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT18), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n245), .A2(new_n247), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G113gat), .B(G141gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(G197gat), .ZN(new_n256));
  XOR2_X1   g055(.A(KEYINPUT11), .B(G169gat), .Z(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n258), .B(KEYINPUT12), .Z(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n251), .A2(new_n243), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n261), .A2(KEYINPUT18), .A3(new_n246), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n254), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n260), .B1(new_n254), .B2(new_n262), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n202), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n254), .A2(new_n262), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n259), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(KEYINPUT100), .A3(new_n263), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G57gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n272), .A2(G64gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT101), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT101), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n275), .B1(new_n272), .B2(G64gat), .ZN(new_n276));
  INV_X1    g075(.A(G64gat), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n274), .B(new_n276), .C1(G57gat), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G71gat), .A2(G78gat), .ZN(new_n279));
  OR2_X1    g078(.A1(G71gat), .A2(G78gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT9), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n277), .A2(G57gat), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT9), .B1(new_n273), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(new_n279), .A3(new_n280), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT21), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G231gat), .A2(G233gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G127gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n212), .B(new_n237), .C1(new_n288), .C2(new_n287), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(G155gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G183gat), .B(G211gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n295), .A2(new_n299), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G85gat), .A2(G92gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n304), .B(KEYINPUT7), .ZN(new_n305));
  NAND2_X1  g104(.A1(G99gat), .A2(G106gat), .ZN(new_n306));
  INV_X1    g105(.A(G85gat), .ZN(new_n307));
  INV_X1    g106(.A(G92gat), .ZN(new_n308));
  AOI22_X1  g107(.A1(KEYINPUT8), .A2(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G99gat), .B(G106gat), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n310), .B(new_n311), .Z(new_n312));
  NAND3_X1  g111(.A1(new_n248), .A2(new_n250), .A3(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n310), .B(new_n311), .ZN(new_n314));
  AND2_X1   g113(.A1(G232gat), .A2(G233gat), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n234), .A2(new_n314), .B1(KEYINPUT41), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G190gat), .B(G218gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n315), .A2(KEYINPUT41), .ZN(new_n320));
  XNOR2_X1  g119(.A(G134gat), .B(G162gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  OR2_X1    g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n319), .A2(new_n322), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G120gat), .B(G148gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(G176gat), .B(G204gat), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n327), .B(new_n328), .Z(new_n329));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n287), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n314), .A2(new_n283), .A3(new_n286), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT104), .ZN(new_n333));
  NAND2_X1  g132(.A1(G230gat), .A2(G233gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n332), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n333), .B1(new_n332), .B2(new_n335), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT10), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n330), .A2(new_n340), .A3(new_n331), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n314), .A2(KEYINPUT10), .A3(new_n283), .A4(new_n286), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(new_n334), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n329), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT106), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n329), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n337), .A2(new_n348), .A3(new_n338), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT102), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n335), .B1(new_n343), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n341), .A2(KEYINPUT102), .A3(new_n342), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(KEYINPUT103), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT103), .B1(new_n351), .B2(new_n352), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n349), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n356), .A2(KEYINPUT105), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT105), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n351), .A2(new_n352), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT103), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n353), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n358), .B1(new_n362), .B2(new_n349), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n347), .B1(new_n357), .B2(new_n363), .ZN(new_n364));
  NOR3_X1   g163(.A1(new_n303), .A2(new_n326), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT2), .ZN(new_n366));
  INV_X1    g165(.A(G141gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(G148gat), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n367), .A2(G148gat), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n366), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G162gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G155gat), .ZN(new_n373));
  INV_X1    g172(.A(G155gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G162gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n373), .A2(new_n375), .ZN(new_n378));
  AND2_X1   g177(.A1(KEYINPUT82), .A2(G148gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(KEYINPUT82), .A2(G148gat), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n379), .A2(new_n380), .A3(new_n367), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n378), .B1(new_n381), .B2(new_n369), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT83), .B(G162gat), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n366), .B1(new_n383), .B2(G155gat), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n377), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G211gat), .B(G218gat), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G211gat), .A2(G218gat), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT77), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT22), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(G197gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(G204gat), .ZN(new_n393));
  INV_X1    g192(.A(G204gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(G197gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n391), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n389), .B1(new_n388), .B2(new_n390), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n387), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n397), .ZN(new_n399));
  XNOR2_X1  g198(.A(G197gat), .B(G204gat), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n399), .A2(new_n386), .A3(new_n400), .A4(new_n391), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT29), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n385), .B1(new_n402), .B2(KEYINPUT3), .ZN(new_n403));
  OR2_X1    g202(.A1(KEYINPUT82), .A2(G148gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(KEYINPUT82), .A2(G148gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(G141gat), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n376), .B1(new_n406), .B2(new_n368), .ZN(new_n407));
  AND2_X1   g206(.A1(KEYINPUT83), .A2(G162gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(KEYINPUT83), .A2(G162gat), .ZN(new_n409));
  OAI21_X1  g208(.A(G155gat), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT2), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n407), .A2(new_n411), .B1(new_n376), .B2(new_n371), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT3), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT29), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n401), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n403), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT87), .B1(new_n414), .B2(new_n415), .ZN(new_n417));
  NAND2_X1  g216(.A1(G228gat), .A2(G233gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n418), .ZN(new_n420));
  OAI221_X1 g219(.A(new_n403), .B1(KEYINPUT87), .B2(new_n420), .C1(new_n414), .C2(new_n415), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(G22gat), .ZN(new_n423));
  INV_X1    g222(.A(G22gat), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n419), .A2(new_n424), .A3(new_n421), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G78gat), .B(G106gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT31), .B(G50gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  AOI21_X1  g228(.A(new_n424), .B1(new_n419), .B2(new_n421), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT88), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n426), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n423), .A2(new_n431), .A3(new_n425), .A4(new_n429), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437));
  INV_X1    g236(.A(G134gat), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n438), .A2(KEYINPUT71), .A3(G127gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(G127gat), .B(G134gat), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n439), .B1(new_n440), .B2(KEYINPUT71), .ZN(new_n441));
  INV_X1    g240(.A(G120gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(G113gat), .ZN(new_n443));
  INV_X1    g242(.A(G113gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(G120gat), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT1), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT72), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n443), .A2(new_n445), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT1), .ZN(new_n451));
  AND4_X1   g250(.A1(new_n449), .A2(new_n450), .A3(new_n440), .A4(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n449), .B1(new_n446), .B2(new_n440), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n448), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n437), .B1(new_n454), .B2(new_n385), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n450), .A2(new_n440), .A3(new_n451), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT72), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n446), .A2(new_n449), .A3(new_n440), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n412), .A2(new_n459), .A3(KEYINPUT4), .A4(new_n448), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n455), .A2(KEYINPUT85), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT85), .B1(new_n455), .B2(new_n460), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT5), .ZN(new_n464));
  NAND2_X1  g263(.A1(G225gat), .A2(G233gat), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n454), .B1(new_n412), .B2(new_n413), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n385), .A2(KEYINPUT3), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n464), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT86), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n465), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n385), .A2(KEYINPUT3), .B1(new_n459), .B2(new_n448), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n412), .A2(new_n413), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT84), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n473), .A2(new_n474), .A3(new_n455), .A4(new_n460), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n455), .A2(new_n460), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT84), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n454), .B(new_n385), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n464), .B1(new_n479), .B2(new_n470), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n475), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n468), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT86), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n482), .B(new_n483), .C1(new_n462), .C2(new_n461), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n469), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G1gat), .B(G29gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT0), .ZN(new_n487));
  XNOR2_X1  g286(.A(G57gat), .B(G85gat), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n487), .B(new_n488), .Z(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n469), .A2(new_n481), .A3(new_n489), .A4(new_n484), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n485), .A2(KEYINPUT6), .A3(new_n490), .ZN(new_n495));
  XNOR2_X1  g294(.A(G8gat), .B(G36gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(KEYINPUT79), .ZN(new_n497));
  XNOR2_X1  g296(.A(G64gat), .B(G92gat), .ZN(new_n498));
  XOR2_X1   g297(.A(new_n497), .B(new_n498), .Z(new_n499));
  INV_X1    g298(.A(G169gat), .ZN(new_n500));
  INV_X1    g299(.A(G176gat), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT23), .ZN(new_n502));
  AND3_X1   g301(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT66), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G183gat), .A2(G190gat), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT67), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT24), .ZN(new_n511));
  NAND3_X1  g310(.A1(KEYINPUT67), .A2(G183gat), .A3(G190gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(G183gat), .A2(G190gat), .ZN(new_n514));
  AND2_X1   g313(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n514), .B1(new_n515), .B2(G190gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT25), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n500), .A2(new_n501), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT23), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n502), .B(KEYINPUT66), .C1(new_n503), .C2(new_n504), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n507), .A2(new_n517), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n511), .ZN(new_n524));
  OR2_X1    g323(.A1(G183gat), .A2(G190gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n520), .A2(G169gat), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT64), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n501), .ZN(new_n530));
  NAND2_X1  g329(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G169gat), .A2(G176gat), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT65), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n519), .A2(new_n520), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n527), .A2(new_n532), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n518), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n508), .ZN(new_n542));
  NAND2_X1  g341(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT27), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT27), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n545), .A2(KEYINPUT68), .A3(G183gat), .ZN(new_n546));
  INV_X1    g345(.A(G190gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT28), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT27), .B(G183gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(KEYINPUT28), .A3(new_n547), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n542), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT69), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n519), .A2(new_n554), .A3(KEYINPUT26), .ZN(new_n555));
  NOR2_X1   g354(.A1(G169gat), .A2(G176gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT26), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT69), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT70), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n556), .A2(new_n560), .A3(new_n557), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT70), .B1(new_n519), .B2(KEYINPUT26), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n559), .A2(new_n537), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n553), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n541), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT29), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n565), .A2(new_n566), .B1(G226gat), .B2(G233gat), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n540), .A2(new_n523), .B1(new_n553), .B2(new_n563), .ZN(new_n568));
  NAND2_X1  g367(.A1(G226gat), .A2(G233gat), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT78), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n569), .B1(new_n568), .B2(KEYINPUT29), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT78), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n415), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n565), .A2(G226gat), .A3(G233gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n572), .A2(new_n576), .A3(new_n415), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n499), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n415), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n573), .B1(new_n572), .B2(new_n576), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT78), .B1(new_n582), .B2(new_n569), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n580), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n499), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n584), .A2(KEYINPUT30), .A3(new_n577), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n579), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g386(.A1(new_n494), .A2(new_n495), .B1(KEYINPUT80), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT80), .ZN(new_n589));
  INV_X1    g388(.A(new_n587), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n584), .A2(new_n577), .A3(new_n585), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT30), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT81), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n591), .A2(KEYINPUT81), .A3(new_n592), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n589), .A2(new_n590), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n436), .B1(new_n588), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n454), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n565), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n541), .A2(new_n564), .A3(new_n454), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT34), .ZN(new_n603));
  INV_X1    g402(.A(G227gat), .ZN(new_n604));
  INV_X1    g403(.A(G233gat), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n602), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n603), .B1(new_n602), .B2(new_n607), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G15gat), .B(G43gat), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT73), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(KEYINPUT74), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n612), .B(KEYINPUT73), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT74), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G71gat), .B(G99gat), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n615), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n619), .B1(new_n615), .B2(new_n618), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n600), .A2(new_n606), .A3(new_n601), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT75), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n623), .A2(KEYINPUT32), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n626), .B1(new_n625), .B2(new_n627), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(KEYINPUT33), .B1(new_n620), .B2(new_n621), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n623), .A2(new_n631), .A3(KEYINPUT32), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT76), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n623), .A2(new_n631), .A3(KEYINPUT76), .A4(KEYINPUT32), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n611), .B1(new_n630), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n623), .A2(new_n624), .ZN(new_n638));
  INV_X1    g437(.A(new_n622), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n627), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT75), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n642));
  AND4_X1   g441(.A1(new_n611), .A2(new_n641), .A3(new_n636), .A4(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT36), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n637), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n641), .A2(new_n636), .A3(new_n642), .ZN(new_n646));
  INV_X1    g445(.A(new_n611), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n641), .A2(new_n636), .A3(new_n611), .A4(new_n642), .ZN(new_n649));
  AOI21_X1  g448(.A(KEYINPUT36), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT89), .B1(new_n598), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n494), .A2(new_n495), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n587), .A2(KEYINPUT80), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n590), .A2(new_n589), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n595), .A2(new_n596), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n653), .A2(new_n654), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n435), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n648), .A2(new_n649), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(new_n644), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT89), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n479), .A2(new_n470), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT39), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n466), .A2(new_n467), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT85), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n477), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n455), .A2(KEYINPUT85), .A3(new_n460), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n666), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n665), .B1(new_n670), .B2(new_n465), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n470), .B1(new_n463), .B2(new_n666), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n671), .B(new_n489), .C1(KEYINPUT39), .C2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT40), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n673), .A2(KEYINPUT90), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n674), .B1(new_n673), .B2(KEYINPUT90), .ZN(new_n676));
  INV_X1    g475(.A(new_n491), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n656), .A2(new_n590), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n435), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT91), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n495), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n653), .B2(KEYINPUT91), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT37), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n584), .A2(new_n684), .A3(new_n577), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n415), .B1(new_n581), .B2(new_n583), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n572), .A2(new_n576), .A3(new_n580), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(KEYINPUT37), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT38), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n685), .A2(new_n688), .A3(new_n689), .A4(new_n499), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n690), .A2(new_n591), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n685), .A2(new_n499), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n684), .B1(new_n584), .B2(new_n577), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT38), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n683), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n696), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n652), .A2(new_n662), .A3(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n637), .A2(new_n643), .A3(new_n435), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT92), .B(KEYINPUT35), .Z(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n701), .A2(new_n683), .A3(new_n679), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n436), .A2(new_n648), .A3(new_n649), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT35), .B1(new_n657), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT93), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n699), .A2(new_n588), .A3(new_n597), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n707), .A2(KEYINPUT93), .A3(KEYINPUT35), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n702), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n271), .B(new_n365), .C1(new_n698), .C2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT107), .ZN(new_n711));
  OR3_X1    g510(.A1(new_n701), .A2(new_n683), .A3(new_n679), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n707), .A2(KEYINPUT93), .A3(KEYINPUT35), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT93), .B1(new_n707), .B2(KEYINPUT35), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n652), .A2(new_n662), .A3(new_n697), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n270), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n717), .A2(new_n718), .A3(new_n365), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n711), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n653), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G1gat), .ZN(G1324gat));
  INV_X1    g522(.A(KEYINPUT42), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n715), .A2(new_n716), .ZN(new_n725));
  AND4_X1   g524(.A1(new_n718), .A2(new_n725), .A3(new_n271), .A4(new_n365), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n718), .B1(new_n717), .B2(new_n365), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n679), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G8gat), .ZN(new_n729));
  XNOR2_X1  g528(.A(KEYINPUT16), .B(G8gat), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n720), .A2(new_n679), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n724), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n679), .ZN(new_n734));
  AOI211_X1 g533(.A(new_n734), .B(new_n730), .C1(new_n711), .C2(new_n719), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(KEYINPUT42), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n733), .A2(KEYINPUT108), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n206), .B1(new_n720), .B2(new_n679), .ZN(new_n739));
  OAI21_X1  g538(.A(KEYINPUT42), .B1(new_n739), .B2(new_n735), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n732), .A2(new_n724), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n737), .A2(new_n742), .ZN(G1325gat));
  INV_X1    g542(.A(new_n720), .ZN(new_n744));
  OR3_X1    g543(.A1(new_n744), .A2(G15gat), .A3(new_n659), .ZN(new_n745));
  OAI21_X1  g544(.A(G15gat), .B1(new_n744), .B2(new_n660), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(G1326gat));
  NAND2_X1  g546(.A1(new_n720), .A2(new_n435), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT43), .B(G22gat), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1327gat));
  INV_X1    g549(.A(new_n364), .ZN(new_n751));
  AND4_X1   g550(.A1(new_n717), .A2(new_n303), .A3(new_n326), .A4(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n752), .A2(new_n217), .A3(new_n721), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT45), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n598), .A2(new_n651), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n697), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT110), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n697), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n709), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n755), .B1(new_n761), .B2(new_n325), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n725), .A2(KEYINPUT44), .A3(new_n326), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n302), .B(KEYINPUT109), .Z(new_n764));
  NAND2_X1  g563(.A1(new_n268), .A2(new_n263), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n764), .A2(new_n765), .A3(new_n751), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n762), .A2(new_n763), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(G29gat), .B1(new_n768), .B2(new_n653), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n769), .ZN(G1328gat));
  NAND3_X1  g569(.A1(new_n752), .A2(new_n218), .A3(new_n679), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT46), .Z(new_n772));
  OAI21_X1  g571(.A(KEYINPUT111), .B1(new_n768), .B2(new_n734), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G36gat), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n768), .A2(KEYINPUT111), .A3(new_n734), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n772), .B1(new_n774), .B2(new_n775), .ZN(G1329gat));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n768), .A2(new_n660), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n225), .ZN(new_n779));
  INV_X1    g578(.A(new_n659), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n752), .A2(new_n225), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(new_n778), .B2(new_n225), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n779), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  OAI221_X1 g583(.A(new_n781), .B1(new_n777), .B2(KEYINPUT47), .C1(new_n778), .C2(new_n225), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(G1330gat));
  NAND4_X1  g585(.A1(new_n762), .A2(new_n435), .A3(new_n763), .A4(new_n767), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G50gat), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n752), .A2(new_n223), .A3(new_n435), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT113), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT48), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n790), .B(new_n791), .ZN(G1331gat));
  NAND2_X1  g591(.A1(new_n758), .A2(new_n760), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n715), .ZN(new_n794));
  NOR4_X1   g593(.A1(new_n751), .A2(new_n765), .A3(new_n303), .A4(new_n326), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(new_n653), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(new_n272), .ZN(G1332gat));
  NOR2_X1   g597(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT116), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n796), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n794), .A2(KEYINPUT114), .A3(new_n795), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n734), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT115), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n806), .A2(KEYINPUT115), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n801), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n809), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n811), .A2(new_n807), .A3(new_n800), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(G1333gat));
  AND2_X1   g612(.A1(new_n803), .A2(new_n804), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n814), .A2(G71gat), .A3(new_n651), .ZN(new_n815));
  INV_X1    g614(.A(G71gat), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n816), .B1(new_n796), .B2(new_n659), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n815), .A2(KEYINPUT50), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT50), .B1(new_n815), .B2(new_n817), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n818), .A2(new_n819), .ZN(G1334gat));
  NAND2_X1  g619(.A1(new_n814), .A2(new_n435), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g621(.A1(new_n302), .A2(new_n765), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n794), .A2(new_n326), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n751), .B1(new_n824), .B2(KEYINPUT51), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n794), .A2(new_n826), .A3(new_n326), .A4(new_n823), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n828), .A2(new_n307), .A3(new_n721), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n823), .A2(new_n364), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n762), .A2(new_n763), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(G85gat), .B1(new_n831), .B2(new_n653), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n829), .A2(new_n832), .ZN(G1336gat));
  OAI211_X1 g632(.A(KEYINPUT52), .B(G92gat), .C1(new_n831), .C2(new_n734), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n734), .A2(G92gat), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n825), .A2(new_n827), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n834), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n825), .A2(new_n837), .A3(new_n827), .A4(new_n835), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT118), .B1(new_n831), .B2(new_n734), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(G92gat), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n831), .A2(KEYINPUT118), .A3(new_n734), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n841), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n840), .B1(new_n845), .B2(new_n838), .ZN(G1337gat));
  INV_X1    g645(.A(G99gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n828), .A2(new_n847), .A3(new_n780), .ZN(new_n848));
  OAI21_X1  g647(.A(G99gat), .B1(new_n831), .B2(new_n660), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(G1338gat));
  NOR2_X1   g649(.A1(new_n436), .A2(G106gat), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n825), .A2(new_n827), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(G106gat), .B1(new_n831), .B2(new_n436), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g653(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n854), .B(new_n855), .ZN(G1339gat));
  OAI22_X1  g655(.A1(new_n245), .A2(new_n247), .B1(new_n261), .B2(new_n246), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n258), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n263), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n364), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n356), .A2(KEYINPUT105), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n362), .A2(new_n358), .A3(new_n349), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT55), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT54), .B1(new_n343), .B2(new_n334), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n866), .B1(new_n361), .B2(new_n353), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n348), .B1(new_n344), .B2(KEYINPUT54), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n865), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n868), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n354), .A2(new_n355), .ZN(new_n871));
  OAI211_X1 g670(.A(KEYINPUT55), .B(new_n870), .C1(new_n871), .C2(new_n866), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n864), .A2(new_n765), .A3(new_n869), .A4(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n326), .B1(new_n861), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n864), .A2(new_n872), .A3(new_n869), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(new_n325), .A3(new_n859), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n764), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n765), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n365), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n703), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n721), .A3(new_n734), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n881), .A2(new_n444), .A3(new_n270), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n721), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n883), .B(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n734), .A3(new_n765), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n882), .B1(new_n886), .B2(new_n444), .ZN(G1340gat));
  NOR2_X1   g686(.A1(new_n751), .A2(G120gat), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n885), .A2(new_n734), .A3(new_n888), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n881), .A2(new_n751), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n890), .A2(KEYINPUT121), .A3(G120gat), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT121), .B1(new_n890), .B2(G120gat), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n889), .B(KEYINPUT122), .C1(new_n891), .C2(new_n892), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1341gat));
  OAI21_X1  g696(.A(G127gat), .B1(new_n881), .B2(new_n764), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n885), .A2(new_n734), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n302), .A2(new_n292), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(G1342gat));
  NOR2_X1   g700(.A1(new_n325), .A2(new_n679), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n438), .A3(new_n902), .ZN(new_n903));
  OR2_X1    g702(.A1(new_n903), .A2(KEYINPUT56), .ZN(new_n904));
  INV_X1    g703(.A(new_n902), .ZN(new_n905));
  OAI21_X1  g704(.A(G134gat), .B1(new_n883), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n903), .A2(KEYINPUT56), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(G1343gat));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n861), .B1(new_n270), .B2(new_n875), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n876), .B1(new_n910), .B2(new_n325), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n879), .B1(new_n911), .B2(new_n302), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n435), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT57), .ZN(new_n914));
  AOI211_X1 g713(.A(KEYINPUT57), .B(new_n436), .C1(new_n877), .C2(new_n879), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n660), .A2(new_n721), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(new_n679), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n914), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n909), .B1(new_n919), .B2(new_n270), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT57), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n921), .B1(new_n912), .B2(new_n435), .ZN(new_n922));
  INV_X1    g721(.A(new_n918), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n922), .A2(new_n915), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(KEYINPUT124), .A3(new_n271), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n920), .A2(G141gat), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n436), .B1(new_n877), .B2(new_n879), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n270), .A2(G141gat), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n927), .A2(new_n918), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(KEYINPUT58), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n914), .A2(new_n916), .A3(new_n765), .A4(new_n918), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n929), .B1(new_n932), .B2(G141gat), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT58), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n929), .ZN(new_n937));
  NOR4_X1   g736(.A1(new_n922), .A2(new_n915), .A3(new_n878), .A4(new_n923), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(new_n367), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT123), .B1(new_n939), .B2(KEYINPUT58), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n931), .B1(new_n936), .B2(new_n940), .ZN(G1344gat));
  INV_X1    g740(.A(new_n927), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n942), .A2(new_n923), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n379), .A2(new_n380), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n943), .A2(new_n944), .A3(new_n364), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT59), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n365), .A2(new_n270), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT125), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n911), .A2(new_n302), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n921), .B(new_n435), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n942), .A2(KEYINPUT57), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n952), .A2(new_n364), .A3(new_n918), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n946), .B1(new_n953), .B2(G148gat), .ZN(new_n954));
  AOI211_X1 g753(.A(KEYINPUT59), .B(new_n944), .C1(new_n924), .C2(new_n364), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n945), .B1(new_n954), .B2(new_n955), .ZN(G1345gat));
  OAI21_X1  g755(.A(G155gat), .B1(new_n919), .B2(new_n764), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n943), .A2(new_n374), .A3(new_n302), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1346gat));
  OAI21_X1  g758(.A(new_n383), .B1(new_n919), .B2(new_n325), .ZN(new_n960));
  OR3_X1    g759(.A1(new_n917), .A2(new_n383), .A3(new_n905), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n960), .B1(new_n942), .B2(new_n961), .ZN(G1347gat));
  NOR2_X1   g761(.A1(new_n734), .A2(new_n721), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n880), .A2(new_n963), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n964), .A2(new_n500), .A3(new_n270), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n877), .A2(new_n879), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(new_n653), .ZN(new_n967));
  OR2_X1    g766(.A1(new_n967), .A2(KEYINPUT126), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n734), .B1(new_n967), .B2(KEYINPUT126), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n968), .A2(new_n699), .A3(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(new_n765), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n965), .B1(new_n972), .B2(new_n500), .ZN(G1348gat));
  AOI21_X1  g772(.A(G176gat), .B1(new_n971), .B2(new_n364), .ZN(new_n974));
  INV_X1    g773(.A(new_n964), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n751), .B1(new_n530), .B2(new_n531), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(G1349gat));
  OAI21_X1  g776(.A(G183gat), .B1(new_n964), .B2(new_n764), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n302), .A2(new_n551), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n978), .B1(new_n970), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g780(.A(G190gat), .B1(new_n964), .B2(new_n325), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n982), .A2(KEYINPUT61), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n982), .A2(KEYINPUT61), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n326), .A2(new_n547), .ZN(new_n985));
  OAI22_X1  g784(.A1(new_n983), .A2(new_n984), .B1(new_n970), .B2(new_n985), .ZN(G1351gat));
  NOR3_X1   g785(.A1(new_n651), .A2(new_n721), .A3(new_n734), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n952), .A2(new_n987), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n988), .A2(new_n392), .A3(new_n270), .ZN(new_n989));
  AND2_X1   g788(.A1(new_n968), .A2(new_n969), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n651), .A2(new_n436), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n990), .A2(KEYINPUT127), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n968), .A2(new_n969), .A3(new_n991), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT127), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n992), .A2(new_n765), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n989), .B1(new_n996), .B2(new_n392), .ZN(G1352gat));
  NAND4_X1  g796(.A1(new_n990), .A2(new_n394), .A3(new_n364), .A4(new_n991), .ZN(new_n998));
  OR2_X1    g797(.A1(new_n998), .A2(KEYINPUT62), .ZN(new_n999));
  OAI21_X1  g798(.A(G204gat), .B1(new_n988), .B2(new_n751), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n998), .A2(KEYINPUT62), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(G1353gat));
  NOR2_X1   g801(.A1(new_n303), .A2(G211gat), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n992), .A2(new_n995), .A3(new_n1003), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n952), .A2(new_n302), .A3(new_n987), .ZN(new_n1005));
  AND3_X1   g804(.A1(new_n1005), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1006));
  AOI21_X1  g805(.A(KEYINPUT63), .B1(new_n1005), .B2(G211gat), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(G1354gat));
  NOR2_X1   g807(.A1(new_n325), .A2(G218gat), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n992), .A2(new_n995), .A3(new_n1009), .ZN(new_n1010));
  OAI21_X1  g809(.A(G218gat), .B1(new_n988), .B2(new_n325), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1010), .A2(new_n1011), .ZN(G1355gat));
endmodule


