//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n829, new_n830, new_n831, new_n832, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G57gat), .ZN(new_n204));
  INV_X1    g003(.A(G85gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT77), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT67), .B(G120gat), .ZN(new_n209));
  INV_X1    g008(.A(G113gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212));
  XNOR2_X1  g011(.A(G127gat), .B(G134gat), .ZN(new_n213));
  OR2_X1    g012(.A1(KEYINPUT67), .A2(G120gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(KEYINPUT67), .A2(G120gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(G113gat), .A3(new_n215), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n211), .A2(new_n212), .A3(new_n213), .A4(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n213), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT1), .B1(G113gat), .B2(G120gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(G113gat), .B2(G120gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT2), .ZN(new_n223));
  INV_X1    g022(.A(G155gat), .ZN(new_n224));
  INV_X1    g023(.A(G162gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT74), .ZN(new_n229));
  INV_X1    g028(.A(G148gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(KEYINPUT74), .A2(G148gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(G141gat), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G141gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(new_n230), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n228), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n223), .B1(G141gat), .B2(G148gat), .ZN(new_n237));
  AND2_X1   g036(.A1(G141gat), .A2(G148gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n227), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT73), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(new_n224), .A3(new_n225), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT73), .B1(G155gat), .B2(G162gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT76), .B1(new_n236), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G141gat), .A2(G148gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n235), .A2(new_n223), .A3(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n247), .A2(new_n227), .A3(new_n242), .A4(new_n241), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n228), .A2(new_n233), .A3(new_n235), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT76), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n222), .B1(new_n245), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT4), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n208), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n248), .A2(new_n249), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n216), .A2(new_n213), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT1), .B1(new_n209), .B2(new_n210), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n257), .A2(new_n258), .B1(new_n218), .B2(new_n220), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n256), .A2(new_n259), .A3(new_n253), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n250), .B1(new_n248), .B2(new_n249), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n263), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n254), .A2(new_n260), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT78), .ZN(new_n266));
  NAND2_X1  g065(.A1(G225gat), .A2(G233gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT3), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n248), .A2(new_n249), .A3(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n222), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT75), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n269), .A2(KEYINPUT75), .A3(new_n222), .A4(new_n271), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n268), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n265), .A2(new_n266), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n266), .B1(new_n265), .B2(new_n276), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n222), .B(new_n255), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(new_n268), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n277), .A2(new_n278), .A3(new_n282), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n222), .A2(new_n253), .A3(new_n255), .ZN(new_n284));
  AOI221_X4 g083(.A(new_n284), .B1(new_n263), .B2(new_n253), .C1(new_n274), .C2(new_n275), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT79), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n285), .A2(new_n286), .A3(new_n279), .A4(new_n267), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n274), .A2(new_n275), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n263), .A2(new_n253), .ZN(new_n289));
  INV_X1    g088(.A(new_n284), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n288), .A2(new_n279), .A3(new_n289), .A4(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT79), .B1(new_n291), .B2(new_n268), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n207), .B1(new_n283), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(KEYINPUT80), .A2(KEYINPUT6), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n265), .A2(new_n276), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT78), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n265), .A2(new_n266), .A3(new_n276), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(new_n281), .A3(new_n298), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n299), .A2(new_n206), .A3(new_n292), .A4(new_n287), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n294), .A2(new_n295), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n292), .A3(new_n287), .ZN(new_n302));
  INV_X1    g101(.A(new_n295), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n207), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G211gat), .B(G218gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n309));
  INV_X1    g108(.A(G197gat), .ZN(new_n310));
  INV_X1    g109(.A(G204gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G197gat), .A2(G204gat), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n309), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(new_n308), .B(new_n314), .Z(new_n315));
  INV_X1    g114(.A(KEYINPUT72), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT64), .ZN(new_n317));
  NOR2_X1   g116(.A1(G169gat), .A2(G176gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n317), .B1(new_n318), .B2(KEYINPUT23), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT23), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n320), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(KEYINPUT23), .ZN(new_n323));
  INV_X1    g122(.A(G183gat), .ZN(new_n324));
  INV_X1    g123(.A(G190gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(KEYINPUT24), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n329), .B1(new_n327), .B2(KEYINPUT24), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n322), .A2(new_n323), .A3(new_n328), .A4(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT25), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n327), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT24), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n330), .B1(new_n337), .B2(new_n326), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n338), .A2(KEYINPUT25), .A3(new_n323), .A4(new_n322), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  OR2_X1    g139(.A1(new_n324), .A2(KEYINPUT27), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT28), .B1(new_n341), .B2(KEYINPUT65), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT27), .B(G183gat), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n342), .B(new_n325), .C1(KEYINPUT65), .C2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n343), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT28), .B1(new_n345), .B2(G190gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT26), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n318), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT66), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n350), .A2(new_n335), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n348), .A2(new_n349), .A3(new_n329), .A4(new_n352), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n344), .A2(new_n346), .A3(new_n351), .A4(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n340), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n355), .A2(new_n356), .B1(G226gat), .B2(G233gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n358), .B1(new_n340), .B2(new_n354), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n316), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n355), .A2(new_n356), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n358), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT72), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n315), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n308), .B(new_n314), .ZN(new_n365));
  NOR3_X1   g164(.A1(new_n357), .A2(new_n365), .A3(new_n359), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G8gat), .B(G36gat), .ZN(new_n368));
  INV_X1    g167(.A(G64gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(G92gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n372), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n374), .B1(new_n364), .B2(new_n366), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(KEYINPUT30), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT30), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n377), .B(new_n374), .C1(new_n364), .C2(new_n366), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n305), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT81), .ZN(new_n381));
  XOR2_X1   g180(.A(G78gat), .B(G106gat), .Z(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT31), .B(G50gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n271), .A2(new_n356), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n315), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT3), .B1(new_n365), .B2(new_n356), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n245), .A2(new_n251), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G228gat), .A2(G233gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(KEYINPUT82), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  OR2_X1    g191(.A1(new_n387), .A2(new_n256), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n390), .B1(new_n315), .B2(new_n385), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n389), .A2(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT83), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n384), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G22gat), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n399), .B1(new_n395), .B2(new_n396), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n395), .A2(new_n396), .A3(new_n399), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n398), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n402), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n397), .B1(new_n404), .B2(new_n400), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT81), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n305), .A2(new_n407), .A3(new_n379), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n381), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT39), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n280), .A2(new_n268), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n412));
  AOI211_X1 g211(.A(new_n410), .B(new_n411), .C1(new_n412), .C2(new_n268), .ZN(new_n413));
  NOR3_X1   g212(.A1(new_n285), .A2(KEYINPUT39), .A3(new_n267), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n413), .A2(new_n414), .A3(new_n207), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n302), .A2(new_n207), .B1(new_n415), .B2(KEYINPUT40), .ZN(new_n416));
  OR2_X1    g215(.A1(new_n415), .A2(KEYINPUT40), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n416), .A2(new_n417), .A3(new_n378), .A4(new_n376), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT6), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n294), .A2(new_n419), .A3(new_n300), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n302), .A2(KEYINPUT6), .A3(new_n207), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT37), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n422), .B1(new_n364), .B2(new_n366), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n360), .A2(new_n363), .A3(new_n315), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n365), .B1(new_n357), .B2(new_n359), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(KEYINPUT37), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT38), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n423), .A2(new_n426), .A3(new_n427), .A4(new_n372), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n420), .A2(new_n421), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n423), .A2(new_n372), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n364), .A2(new_n422), .A3(new_n366), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT38), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n375), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n418), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n406), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n409), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n340), .A2(new_n259), .A3(new_n354), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT68), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n355), .A2(new_n222), .ZN(new_n441));
  NAND2_X1  g240(.A1(G227gat), .A2(G233gat), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n340), .A2(new_n354), .A3(KEYINPUT68), .A4(new_n259), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  XOR2_X1   g243(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT32), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n448));
  INV_X1    g247(.A(new_n442), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT33), .B1(new_n448), .B2(new_n449), .ZN(new_n451));
  XNOR2_X1  g250(.A(G15gat), .B(G43gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n452), .B(G71gat), .ZN(new_n453));
  INV_X1    g252(.A(G99gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n450), .A2(new_n451), .A3(new_n456), .ZN(new_n457));
  AOI221_X4 g256(.A(new_n447), .B1(KEYINPUT33), .B2(new_n455), .C1(new_n448), .C2(new_n449), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n446), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n451), .A2(new_n456), .ZN(new_n460));
  INV_X1    g259(.A(new_n450), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n446), .ZN(new_n463));
  INV_X1    g262(.A(new_n458), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT70), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n459), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT36), .ZN(new_n468));
  OAI211_X1 g267(.A(KEYINPUT70), .B(new_n446), .C1(new_n457), .C2(new_n458), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n459), .A2(new_n465), .A3(KEYINPUT36), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n437), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n406), .B1(new_n469), .B2(new_n467), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n379), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(KEYINPUT84), .B(KEYINPUT35), .Z(new_n478));
  AOI21_X1  g277(.A(new_n478), .B1(new_n420), .B2(new_n421), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n459), .A2(new_n465), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n406), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n381), .A2(new_n481), .A3(new_n408), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n477), .A2(new_n479), .B1(new_n482), .B2(KEYINPUT35), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n473), .A2(new_n483), .ZN(new_n484));
  XOR2_X1   g283(.A(G15gat), .B(G22gat), .Z(new_n485));
  INV_X1    g284(.A(G1gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G15gat), .B(G22gat), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT16), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n488), .B1(new_n489), .B2(G1gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT89), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(G8gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n487), .B(new_n490), .C1(new_n492), .C2(G8gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(KEYINPUT90), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT90), .B1(new_n495), .B2(new_n496), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(G71gat), .B(G78gat), .Z(new_n501));
  INV_X1    g300(.A(KEYINPUT92), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n502), .A2(new_n369), .A3(G57gat), .ZN(new_n503));
  INV_X1    g302(.A(G57gat), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT92), .B1(new_n504), .B2(G64gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(G64gat), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT93), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n501), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT9), .ZN(new_n510));
  INV_X1    g309(.A(G71gat), .ZN(new_n511));
  INV_X1    g310(.A(G78gat), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n509), .B(new_n513), .C1(new_n508), .C2(new_n507), .ZN(new_n514));
  XNOR2_X1  g313(.A(G57gat), .B(G64gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n501), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(KEYINPUT21), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n514), .A2(new_n516), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT21), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n500), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n499), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n497), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(new_n519), .A3(new_n518), .ZN(new_n524));
  XOR2_X1   g323(.A(G127gat), .B(G155gat), .Z(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n521), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n526), .B1(new_n521), .B2(new_n524), .ZN(new_n528));
  INV_X1    g327(.A(G231gat), .ZN(new_n529));
  INV_X1    g328(.A(G233gat), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OR3_X1    g330(.A1(new_n527), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n531), .B1(new_n527), .B2(new_n528), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G183gat), .B(G211gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT20), .ZN(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n532), .A2(new_n533), .A3(new_n538), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G85gat), .A2(G92gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  NAND2_X1  g343(.A1(G99gat), .A2(G106gat), .ZN(new_n545));
  AOI22_X1  g344(.A1(KEYINPUT8), .A2(new_n545), .B1(new_n205), .B2(new_n371), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n546), .A2(KEYINPUT96), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(KEYINPUT96), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G99gat), .B(G106gat), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n550), .B(new_n544), .C1(new_n547), .C2(new_n548), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G43gat), .B(G50gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT87), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT15), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(G50gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n558), .A2(KEYINPUT87), .A3(G43gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n555), .A2(KEYINPUT15), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT14), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n562), .B1(G29gat), .B2(G36gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(G29gat), .A2(G36gat), .ZN(new_n564));
  MUX2_X1   g363(.A(new_n563), .B(new_n562), .S(new_n564), .Z(new_n565));
  NAND3_X1  g364(.A1(new_n560), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT88), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n565), .A2(new_n561), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n567), .B1(new_n570), .B2(new_n566), .ZN(new_n571));
  NOR3_X1   g370(.A1(new_n569), .A2(new_n571), .A3(KEYINPUT17), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n566), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT88), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n573), .B1(new_n575), .B2(new_n568), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n554), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n577), .A2(KEYINPUT97), .B1(KEYINPUT41), .B2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G190gat), .B(G218gat), .Z(new_n580));
  NAND2_X1  g379(.A1(new_n575), .A2(new_n568), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n581), .A2(new_n553), .A3(new_n552), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT97), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n583), .B(new_n554), .C1(new_n572), .C2(new_n576), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n579), .A2(new_n580), .A3(new_n582), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT98), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n579), .A2(new_n582), .A3(new_n584), .ZN(new_n587));
  INV_X1    g386(.A(new_n580), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n578), .A2(KEYINPUT41), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT95), .ZN(new_n591));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n586), .A2(new_n589), .A3(new_n585), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n586), .A2(new_n593), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n589), .A2(new_n585), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n554), .A2(new_n518), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n552), .A2(new_n514), .A3(new_n553), .A4(new_n516), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G230gat), .A2(G233gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT99), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n600), .A2(KEYINPUT99), .A3(new_n602), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT100), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT10), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n599), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n598), .A2(new_n609), .A3(new_n599), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n602), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G120gat), .B(G148gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT101), .ZN(new_n614));
  INV_X1    g413(.A(G176gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(new_n311), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT100), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n605), .A2(new_n619), .A3(new_n606), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n608), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n617), .B1(new_n607), .B2(new_n612), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n542), .A2(new_n594), .A3(new_n597), .A4(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(KEYINPUT102), .Z(new_n626));
  INV_X1    g425(.A(KEYINPUT91), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n569), .A2(new_n571), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n627), .B1(new_n500), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n523), .A2(new_n581), .A3(KEYINPUT91), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G229gat), .A2(G233gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n495), .A2(new_n496), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n572), .B2(new_n576), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT18), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n500), .A2(new_n628), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n631), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n632), .B(KEYINPUT13), .Z(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n631), .A2(KEYINPUT18), .A3(new_n632), .A4(new_n634), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n637), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G113gat), .B(G141gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(G197gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT11), .ZN(new_n646));
  INV_X1    g445(.A(G169gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT85), .B(KEYINPUT12), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n648), .B(new_n649), .Z(new_n650));
  AND3_X1   g449(.A1(new_n643), .A2(KEYINPUT86), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n650), .B1(new_n643), .B2(KEYINPUT86), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n484), .A2(new_n626), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT103), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT103), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n484), .A2(new_n656), .A3(new_n626), .A4(new_n653), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n305), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g460(.A1(new_n489), .A2(new_n494), .ZN(new_n662));
  AOI211_X1 g461(.A(new_n379), .B(new_n662), .C1(new_n655), .C2(new_n657), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n489), .A2(new_n494), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT42), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n658), .A2(new_n476), .ZN(new_n668));
  AOI22_X1  g467(.A1(new_n663), .A2(new_n664), .B1(new_n668), .B2(G8gat), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n667), .B1(new_n669), .B2(new_n666), .ZN(G1325gat));
  INV_X1    g469(.A(G15gat), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n472), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n470), .A2(KEYINPUT104), .A3(new_n471), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n671), .B1(new_n658), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n467), .A2(new_n469), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  AOI211_X1 g479(.A(G15gat), .B(new_n680), .C1(new_n655), .C2(new_n657), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n678), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT105), .B1(new_n677), .B2(new_n681), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(G1326gat));
  NAND2_X1  g485(.A1(new_n658), .A2(new_n406), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT43), .B(G22gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  NAND2_X1  g488(.A1(new_n597), .A2(new_n594), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n484), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n653), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(new_n542), .A3(new_n623), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n694), .A2(G29gat), .A3(new_n305), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n483), .ZN(new_n698));
  AOI221_X4 g497(.A(KEYINPUT106), .B1(new_n673), .B2(new_n674), .C1(new_n409), .C2(new_n436), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n437), .B2(new_n675), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n698), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT44), .B1(new_n702), .B2(new_n690), .ZN(new_n703));
  OAI211_X1 g502(.A(KEYINPUT44), .B(new_n690), .C1(new_n473), .C2(new_n483), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n693), .ZN(new_n707));
  OAI21_X1  g506(.A(G29gat), .B1(new_n707), .B2(new_n305), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n697), .A2(new_n708), .ZN(G1328gat));
  OR3_X1    g508(.A1(new_n694), .A2(G36gat), .A3(new_n379), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n710), .A2(KEYINPUT46), .ZN(new_n711));
  OAI21_X1  g510(.A(G36gat), .B1(new_n707), .B2(new_n379), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(KEYINPUT46), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(G1329gat));
  NAND4_X1  g513(.A1(new_n706), .A2(G43gat), .A3(new_n676), .A4(new_n693), .ZN(new_n715));
  INV_X1    g514(.A(G43gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(new_n694), .B2(new_n680), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n690), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n722), .A2(new_n406), .A3(new_n704), .A4(new_n693), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G50gat), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT48), .B1(new_n724), .B2(KEYINPUT107), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n691), .A2(new_n558), .A3(new_n406), .A4(new_n693), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n724), .B(new_n726), .C1(KEYINPUT107), .C2(KEYINPUT48), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(G1331gat));
  INV_X1    g529(.A(new_n542), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(new_n690), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n702), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n653), .A2(new_n624), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n305), .B(KEYINPUT108), .Z(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(new_n504), .ZN(G1332gat));
  NOR2_X1   g537(.A1(new_n735), .A2(new_n379), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  AND2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n739), .B2(new_n740), .ZN(G1333gat));
  OAI21_X1  g542(.A(new_n511), .B1(new_n735), .B2(new_n680), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n676), .A2(G71gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n735), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g546(.A1(new_n735), .A2(new_n435), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(new_n512), .ZN(G1335gat));
  NOR2_X1   g548(.A1(new_n653), .A2(new_n542), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n706), .A2(new_n623), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G85gat), .B1(new_n751), .B2(new_n305), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n702), .A2(new_n690), .A3(new_n750), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT51), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n702), .A2(new_n755), .A3(new_n690), .A4(new_n750), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n623), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n659), .A2(new_n205), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n752), .B1(new_n759), .B2(new_n760), .ZN(G1336gat));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n762));
  AOI22_X1  g561(.A1(new_n754), .A2(new_n756), .B1(new_n762), .B2(new_n753), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n379), .A2(G92gat), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n623), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n753), .A2(new_n762), .A3(new_n755), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n763), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n750), .ZN(new_n768));
  NOR4_X1   g567(.A1(new_n703), .A2(new_n705), .A3(new_n624), .A4(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n371), .B1(new_n769), .B2(new_n476), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT52), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(G92gat), .B1(new_n751), .B2(new_n379), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n758), .A2(new_n623), .A3(new_n764), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n771), .A2(new_n775), .ZN(G1337gat));
  NOR3_X1   g575(.A1(new_n751), .A2(new_n454), .A3(new_n675), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n758), .A2(new_n623), .A3(new_n679), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n454), .ZN(G1338gat));
  INV_X1    g578(.A(G106gat), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n406), .A2(new_n780), .A3(new_n623), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n763), .A2(new_n766), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n780), .B1(new_n769), .B2(new_n406), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT53), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n757), .B2(new_n781), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(new_n787), .ZN(G1339gat));
  NOR2_X1   g587(.A1(new_n625), .A2(new_n653), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n610), .A2(new_n611), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n601), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n610), .A2(new_n611), .A3(new_n602), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(KEYINPUT54), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  INV_X1    g593(.A(new_n617), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n612), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n793), .A2(new_n794), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n794), .B1(new_n793), .B2(new_n797), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n621), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT110), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT110), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n803), .B(new_n621), .C1(new_n799), .C2(new_n800), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n637), .A2(new_n641), .A3(new_n642), .A4(new_n650), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n639), .A2(new_n640), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n632), .B1(new_n631), .B2(new_n634), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n648), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n805), .A2(new_n690), .A3(new_n810), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n623), .A2(new_n806), .A3(new_n809), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n805), .B2(new_n653), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n813), .B2(new_n690), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n789), .B1(new_n814), .B2(new_n731), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n815), .A2(new_n476), .A3(new_n736), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n816), .A2(new_n481), .ZN(new_n817));
  XOR2_X1   g616(.A(new_n817), .B(KEYINPUT111), .Z(new_n818));
  NAND3_X1  g617(.A1(new_n818), .A2(new_n210), .A3(new_n653), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n815), .A2(new_n475), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n476), .A2(new_n305), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(G113gat), .B1(new_n822), .B2(new_n692), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n823), .ZN(G1340gat));
  INV_X1    g623(.A(G120gat), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n818), .A2(new_n825), .A3(new_n623), .ZN(new_n826));
  OAI21_X1  g625(.A(G120gat), .B1(new_n822), .B2(new_n624), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(G1341gat));
  INV_X1    g627(.A(G127gat), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n822), .A2(new_n829), .A3(new_n731), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n817), .A2(new_n542), .ZN(new_n831));
  XOR2_X1   g630(.A(new_n831), .B(KEYINPUT112), .Z(new_n832));
  AOI21_X1  g631(.A(new_n830), .B1(new_n832), .B2(new_n829), .ZN(G1342gat));
  INV_X1    g632(.A(G134gat), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n817), .A2(new_n834), .A3(new_n690), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT56), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(KEYINPUT114), .Z(new_n837));
  NOR2_X1   g636(.A1(new_n835), .A2(KEYINPUT56), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n838), .B(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n690), .ZN(new_n841));
  OAI21_X1  g640(.A(G134gat), .B1(new_n822), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n837), .A2(new_n840), .A3(new_n842), .ZN(G1343gat));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n675), .A2(new_n821), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n805), .A2(new_n690), .A3(new_n810), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n643), .A2(KEYINPUT86), .ZN(new_n848));
  INV_X1    g647(.A(new_n650), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n621), .ZN(new_n851));
  INV_X1    g650(.A(new_n800), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(new_n798), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n643), .A2(KEYINPUT86), .A3(new_n650), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n850), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n812), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n690), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n731), .B1(new_n847), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n789), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n435), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n846), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n815), .A2(KEYINPUT57), .A3(new_n435), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n862), .A2(new_n863), .A3(KEYINPUT115), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT115), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n855), .A2(new_n856), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n841), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n542), .B1(new_n867), .B2(new_n811), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n406), .B1(new_n868), .B2(new_n789), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n845), .B1(new_n869), .B2(KEYINPUT57), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n814), .A2(new_n731), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n861), .B(new_n406), .C1(new_n871), .C2(new_n789), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n865), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n864), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n844), .B(G141gat), .C1(new_n874), .C2(new_n692), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT115), .B1(new_n862), .B2(new_n863), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n870), .A2(new_n872), .A3(new_n865), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n692), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT116), .B1(new_n878), .B2(new_n234), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n675), .A2(new_n406), .ZN(new_n880));
  NOR4_X1   g679(.A1(new_n815), .A2(new_n476), .A3(new_n880), .A4(new_n736), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n234), .A3(new_n653), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n875), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT58), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n882), .B(KEYINPUT117), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n870), .A2(new_n872), .A3(new_n653), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT58), .B1(new_n886), .B2(G141gat), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n884), .A2(new_n888), .ZN(G1344gat));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n626), .A2(new_n692), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n893), .B1(new_n841), .B2(new_n801), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n690), .A2(KEYINPUT119), .A3(new_n853), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n810), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n542), .B1(new_n896), .B2(new_n867), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n861), .B(new_n406), .C1(new_n892), .C2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT57), .B1(new_n815), .B2(new_n435), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n898), .A2(new_n623), .A3(new_n846), .A4(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n891), .B1(new_n900), .B2(G148gat), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n876), .A2(new_n877), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT59), .B1(new_n902), .B2(new_n623), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n231), .A2(new_n232), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n901), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n881), .A2(new_n904), .A3(new_n623), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT118), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n908), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n890), .B1(new_n906), .B2(new_n912), .ZN(new_n913));
  AOI211_X1 g712(.A(KEYINPUT59), .B(new_n904), .C1(new_n902), .C2(new_n623), .ZN(new_n914));
  OAI211_X1 g713(.A(KEYINPUT120), .B(new_n911), .C1(new_n914), .C2(new_n901), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1345gat));
  AOI21_X1  g715(.A(G155gat), .B1(new_n881), .B2(new_n542), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n874), .A2(new_n731), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g718(.A(G162gat), .B1(new_n881), .B2(new_n690), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n874), .A2(new_n841), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(G162gat), .ZN(G1347gat));
  OAI211_X1 g721(.A(new_n305), .B(new_n476), .C1(new_n871), .C2(new_n789), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n923), .A2(new_n406), .A3(new_n480), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(new_n647), .A3(new_n653), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n736), .A2(new_n476), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT121), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n820), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G169gat), .B1(new_n928), .B2(new_n692), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n925), .A2(new_n929), .ZN(G1348gat));
  NOR3_X1   g729(.A1(new_n928), .A2(new_n615), .A3(new_n624), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n924), .A2(new_n623), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n932), .B2(new_n615), .ZN(G1349gat));
  INV_X1    g732(.A(new_n928), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n324), .B1(new_n934), .B2(new_n542), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n731), .A2(new_n345), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n924), .B2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n938), .A2(KEYINPUT60), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(KEYINPUT60), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT123), .Z(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  OR3_X1    g741(.A1(new_n937), .A2(new_n939), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n937), .B2(new_n939), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1350gat));
  NAND3_X1  g744(.A1(new_n924), .A2(new_n325), .A3(new_n690), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n325), .B1(new_n934), .B2(new_n690), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n948));
  OR2_X1    g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n947), .A2(new_n948), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n950), .B1(new_n949), .B2(new_n951), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n946), .B1(new_n952), .B2(new_n953), .ZN(G1351gat));
  NAND2_X1  g753(.A1(new_n927), .A2(new_n675), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT125), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n898), .A2(new_n899), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(G197gat), .B1(new_n958), .B2(new_n692), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n923), .A2(new_n880), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n960), .A2(new_n310), .A3(new_n653), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(G1352gat));
  OAI21_X1  g761(.A(G204gat), .B1(new_n958), .B2(new_n624), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n960), .A2(new_n311), .A3(new_n623), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(KEYINPUT62), .ZN(new_n965));
  OR2_X1    g764(.A1(new_n964), .A2(KEYINPUT62), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(G1353gat));
  NAND2_X1  g766(.A1(new_n957), .A2(new_n542), .ZN(new_n968));
  OAI21_X1  g767(.A(G211gat), .B1(new_n968), .B2(new_n955), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n969), .A2(KEYINPUT63), .ZN(new_n970));
  INV_X1    g769(.A(G211gat), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n960), .A2(new_n971), .A3(new_n542), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT126), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n969), .A2(KEYINPUT63), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n970), .A2(new_n973), .A3(new_n974), .ZN(G1354gat));
  INV_X1    g774(.A(G218gat), .ZN(new_n976));
  NOR3_X1   g775(.A1(new_n958), .A2(new_n976), .A3(new_n841), .ZN(new_n977));
  INV_X1    g776(.A(new_n960), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n976), .B1(new_n978), .B2(new_n841), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n979), .A2(KEYINPUT127), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n979), .A2(KEYINPUT127), .ZN(new_n981));
  NOR3_X1   g780(.A1(new_n977), .A2(new_n980), .A3(new_n981), .ZN(G1355gat));
endmodule


