//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT72), .ZN(new_n188));
  NOR2_X1   g002(.A1(G472), .A2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G134), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(G134), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT64), .A3(G137), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G131), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT11), .B1(new_n195), .B2(G137), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT11), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(new_n192), .A3(G134), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G131), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n192), .A2(G134), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n210), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n209), .A2(new_n211), .A3(G143), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n213), .B(G146), .C1(new_n209), .C2(KEYINPUT1), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n197), .A2(KEYINPUT65), .A3(G131), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n200), .A2(new_n208), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n212), .A2(new_n214), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT0), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(new_n209), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n221), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n212), .B(new_n214), .C1(new_n222), .C2(new_n209), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI211_X1 g041(.A(G131), .B(new_n206), .C1(new_n201), .C2(new_n203), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n205), .B1(new_n204), .B2(new_n207), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n220), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(G116), .B(G119), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  OR2_X1    g047(.A1(KEYINPUT2), .A2(G113), .ZN(new_n234));
  AND3_X1   g048(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n232), .B(new_n234), .C1(new_n236), .C2(new_n235), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT67), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(new_n239), .A3(KEYINPUT67), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n231), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n208), .A2(new_n218), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n197), .A2(KEYINPUT65), .A3(G131), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT65), .B1(new_n197), .B2(G131), .ZN(new_n247));
  NOR3_X1   g061(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n229), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n249), .A2(new_n208), .B1(new_n225), .B2(new_n226), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT30), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT30), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n220), .A2(new_n230), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n244), .B1(new_n254), .B2(new_n243), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n256), .B(G101), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT68), .B(G953), .ZN(new_n258));
  INV_X1    g072(.A(G237), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(G210), .A3(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n257), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT70), .B(KEYINPUT31), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n255), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n220), .A2(new_n252), .A3(new_n230), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n252), .B1(new_n220), .B2(new_n230), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n243), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OR2_X1    g080(.A1(new_n231), .A2(new_n243), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n261), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n266), .A2(KEYINPUT69), .A3(new_n261), .A4(new_n267), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n263), .B1(new_n272), .B2(KEYINPUT31), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n244), .A2(KEYINPUT28), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n231), .A2(new_n243), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n267), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT71), .B(KEYINPUT28), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n274), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OR2_X1    g092(.A1(new_n278), .A2(new_n261), .ZN(new_n279));
  AOI211_X1 g093(.A(new_n188), .B(new_n190), .C1(new_n273), .C2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT69), .B1(new_n255), .B2(new_n261), .ZN(new_n281));
  INV_X1    g095(.A(new_n271), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT31), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n263), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(new_n279), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT72), .B1(new_n285), .B2(new_n189), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n187), .B1(new_n280), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT29), .B1(new_n278), .B2(new_n261), .ZN(new_n288));
  INV_X1    g102(.A(new_n255), .ZN(new_n289));
  INV_X1    g103(.A(new_n261), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n276), .A2(KEYINPUT28), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(new_n274), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n276), .A2(KEYINPUT73), .A3(KEYINPUT28), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n295), .A2(KEYINPUT29), .A3(new_n261), .A4(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n292), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G472), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n285), .A2(KEYINPUT32), .A3(new_n189), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n287), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G214), .B1(G237), .B2(G902), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G107), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(KEYINPUT83), .A3(G104), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT3), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n307), .A2(G104), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n312), .A2(new_n307), .A3(KEYINPUT83), .A4(G104), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n309), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(new_n315), .A3(G101), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(G101), .ZN(new_n317));
  INV_X1    g131(.A(G101), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n309), .A2(new_n311), .A3(new_n318), .A4(new_n313), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(KEYINPUT4), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n242), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n316), .B(new_n320), .C1(new_n321), .C2(new_n240), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT5), .ZN(new_n323));
  INV_X1    g137(.A(G119), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n324), .A3(G116), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n233), .B2(new_n323), .ZN(new_n326));
  INV_X1    g140(.A(G113), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n239), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G104), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(G107), .ZN(new_n330));
  OAI21_X1  g144(.A(G101), .B1(new_n310), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n319), .A2(new_n331), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G110), .B(G122), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n322), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT85), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT85), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n322), .A2(new_n333), .A3(new_n337), .A4(new_n334), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n322), .A2(new_n333), .ZN(new_n339));
  INV_X1    g153(.A(new_n334), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n336), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT86), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n339), .A2(new_n343), .A3(new_n340), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT6), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n339), .A2(new_n343), .A3(KEYINPUT6), .A4(new_n340), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n342), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n227), .A2(G125), .ZN(new_n349));
  INV_X1    g163(.A(new_n218), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n349), .B1(G125), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G953), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G224), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n351), .B(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n336), .A2(new_n338), .ZN(new_n356));
  XOR2_X1   g170(.A(new_n334), .B(KEYINPUT8), .Z(new_n357));
  NAND2_X1  g171(.A1(new_n328), .A2(new_n332), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n357), .B1(new_n333), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n351), .B(KEYINPUT87), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n353), .A2(KEYINPUT7), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n351), .A2(KEYINPUT87), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n356), .B(new_n362), .C1(new_n361), .C2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n355), .A2(new_n298), .A3(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G210), .B1(G237), .B2(G902), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(G902), .B1(new_n348), .B2(new_n354), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(new_n366), .A3(new_n364), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n306), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G475), .ZN(new_n372));
  AND2_X1   g186(.A1(KEYINPUT68), .A2(G953), .ZN(new_n373));
  NOR2_X1   g187(.A1(KEYINPUT68), .A2(G953), .ZN(new_n374));
  OAI211_X1 g188(.A(G214), .B(new_n259), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n213), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n258), .A2(G143), .A3(G214), .A4(new_n259), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(new_n377), .A3(new_n205), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT88), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(new_n377), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G131), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT17), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT88), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n376), .A2(new_n377), .A3(new_n383), .A4(new_n205), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n379), .A2(new_n381), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G140), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G125), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(KEYINPUT16), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G125), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(KEYINPUT75), .A3(G140), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT75), .ZN(new_n393));
  XNOR2_X1  g207(.A(G125), .B(G140), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT16), .ZN(new_n396));
  OAI211_X1 g210(.A(G146), .B(new_n389), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n390), .A2(G140), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(new_n387), .A3(new_n393), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n396), .B1(new_n399), .B2(new_n391), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n211), .B1(new_n400), .B2(new_n388), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n380), .A2(KEYINPUT17), .A3(G131), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n385), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT76), .B1(new_n394), .B2(new_n211), .ZN(new_n405));
  AND4_X1   g219(.A1(KEYINPUT76), .A2(new_n398), .A3(new_n387), .A4(new_n211), .ZN(new_n406));
  OR2_X1    g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n399), .A2(new_n391), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n407), .B1(new_n211), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT18), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n376), .B(new_n377), .C1(new_n410), .C2(new_n205), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n409), .B(new_n411), .C1(new_n410), .C2(new_n381), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n404), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(G113), .B(G122), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(new_n329), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(KEYINPUT91), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(G902), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n404), .A2(new_n412), .A3(new_n416), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n372), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n413), .A2(new_n415), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n399), .A2(KEYINPUT19), .A3(new_n391), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT19), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT89), .B1(new_n394), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n399), .A2(KEYINPUT89), .A3(KEYINPUT19), .A4(new_n391), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n211), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT90), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n379), .A2(new_n381), .A3(new_n384), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT90), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n427), .A2(new_n431), .A3(new_n211), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n429), .A2(new_n397), .A3(new_n430), .A4(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n415), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n434), .A3(new_n412), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n421), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT20), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n436), .A2(new_n437), .A3(new_n372), .A4(new_n298), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n421), .A2(new_n435), .A3(new_n372), .A4(new_n298), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT20), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n420), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT97), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n213), .A2(G128), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n213), .A2(KEYINPUT93), .A3(G128), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT93), .B1(new_n213), .B2(G128), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n444), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n448), .A2(G134), .ZN(new_n449));
  INV_X1    g263(.A(G122), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G116), .ZN(new_n451));
  INV_X1    g265(.A(G116), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G122), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT92), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT92), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n451), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G107), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n455), .A2(new_n307), .A3(new_n457), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT13), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT94), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT94), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT13), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n446), .B2(new_n447), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT95), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n468), .A3(new_n444), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT93), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n470), .B1(new_n209), .B2(G143), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n471), .A2(new_n445), .B1(new_n463), .B2(new_n465), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT95), .B1(new_n472), .B2(new_n443), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n471), .A2(new_n445), .A3(new_n463), .A4(new_n465), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n469), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n449), .B(new_n461), .C1(new_n475), .C2(new_n195), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n452), .A2(KEYINPUT14), .A3(G122), .ZN(new_n477));
  OAI211_X1 g291(.A(G107), .B(new_n477), .C1(new_n454), .C2(KEYINPUT14), .ZN(new_n478));
  XOR2_X1   g292(.A(new_n478), .B(KEYINPUT96), .Z(new_n479));
  XNOR2_X1  g293(.A(new_n448), .B(G134), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(new_n480), .A3(new_n460), .ZN(new_n481));
  XOR2_X1   g295(.A(KEYINPUT9), .B(G234), .Z(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(G217), .A3(new_n352), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n476), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n484), .B1(new_n476), .B2(new_n481), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n442), .B(new_n298), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G478), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n489), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n476), .A2(new_n481), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n483), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n476), .A2(new_n481), .A3(new_n484), .ZN(new_n494));
  AOI21_X1  g308(.A(G902), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n491), .B1(new_n495), .B2(new_n442), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n490), .B1(new_n496), .B2(new_n487), .ZN(new_n497));
  INV_X1    g311(.A(G952), .ZN(new_n498));
  AOI211_X1 g312(.A(G953), .B(new_n498), .C1(G234), .C2(G237), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI211_X1 g314(.A(new_n298), .B(new_n258), .C1(G234), .C2(G237), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT21), .B(G898), .Z(new_n503));
  OAI21_X1  g317(.A(new_n500), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n441), .A2(new_n497), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(G469), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n228), .A2(new_n229), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n218), .A2(new_n319), .A3(new_n331), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n218), .B1(new_n319), .B2(new_n331), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT12), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n320), .A2(new_n227), .A3(new_n316), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT84), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT10), .ZN(new_n516));
  OR2_X1    g330(.A1(new_n509), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n515), .A2(KEYINPUT10), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n516), .B1(new_n509), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n514), .A2(new_n517), .A3(new_n507), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n258), .A2(G227), .ZN(new_n521));
  XNOR2_X1  g335(.A(G110), .B(G140), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n513), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n514), .A2(new_n517), .A3(new_n519), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n508), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n523), .B1(new_n527), .B2(new_n520), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n506), .B(new_n298), .C1(new_n525), .C2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(G469), .A2(G902), .ZN(new_n530));
  INV_X1    g344(.A(new_n523), .ZN(new_n531));
  INV_X1    g345(.A(new_n520), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n531), .B1(new_n513), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n527), .A2(new_n520), .A3(new_n523), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(G469), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n529), .A2(new_n530), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G221), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n537), .B1(new_n482), .B2(new_n298), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n371), .A2(new_n505), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT79), .ZN(new_n543));
  OAI211_X1 g357(.A(G221), .B(G234), .C1(new_n373), .C2(new_n374), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT78), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT78), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n258), .A2(new_n546), .A3(G221), .A4(G234), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT22), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n548), .B1(new_n545), .B2(new_n547), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n550), .A2(new_n551), .A3(new_n192), .ZN(new_n552));
  OR2_X1    g366(.A1(KEYINPUT68), .A2(G953), .ZN(new_n553));
  NAND2_X1  g367(.A1(KEYINPUT68), .A2(G953), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n537), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n546), .B1(new_n555), .B2(G234), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n544), .A2(KEYINPUT78), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT22), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(G137), .B1(new_n558), .B2(new_n549), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n543), .B1(new_n552), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n192), .B1(new_n550), .B2(new_n551), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n558), .A2(G137), .A3(new_n549), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n562), .A3(KEYINPUT79), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT23), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n565), .B1(new_n324), .B2(G128), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n566), .B(new_n567), .C1(G119), .C2(new_n209), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT74), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n209), .B2(G119), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n324), .A2(KEYINPUT74), .A3(G128), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n570), .A2(new_n571), .B1(G119), .B2(new_n209), .ZN(new_n572));
  XOR2_X1   g386(.A(KEYINPUT24), .B(G110), .Z(new_n573));
  OAI22_X1  g387(.A1(G110), .A2(new_n568), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n397), .A2(new_n574), .A3(new_n407), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT77), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n405), .A2(new_n406), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n388), .B1(new_n408), .B2(KEYINPUT16), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n578), .B1(new_n579), .B2(G146), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(KEYINPUT77), .A3(new_n574), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n397), .A2(new_n401), .ZN(new_n582));
  AOI22_X1  g396(.A1(G110), .A2(new_n568), .B1(new_n572), .B2(new_n573), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n577), .A2(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT80), .B1(new_n564), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(new_n583), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT77), .B1(new_n580), .B2(new_n574), .ZN(new_n587));
  AND4_X1   g401(.A1(KEYINPUT77), .A2(new_n397), .A3(new_n574), .A4(new_n407), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT80), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n589), .A2(new_n590), .A3(new_n563), .A4(new_n560), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n585), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n584), .B1(new_n552), .B2(new_n559), .ZN(new_n593));
  AND2_X1   g407(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n594));
  NOR2_X1   g408(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n592), .A2(new_n298), .A3(new_n593), .A4(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(G217), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(G234), .B2(new_n298), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n585), .A2(new_n298), .A3(new_n593), .A4(new_n591), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n600), .B1(new_n601), .B2(new_n594), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT82), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n597), .A2(new_n602), .A3(KEYINPUT82), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n592), .A2(new_n593), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n599), .A2(G902), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n605), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n304), .A2(new_n542), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G101), .ZN(G3));
  INV_X1    g428(.A(KEYINPUT31), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n270), .B2(new_n271), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n278), .A2(new_n261), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n616), .A2(new_n617), .A3(new_n263), .ZN(new_n618));
  OAI21_X1  g432(.A(G472), .B1(new_n618), .B2(G902), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n619), .B1(new_n280), .B2(new_n286), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n611), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n541), .ZN(new_n622));
  XOR2_X1   g436(.A(new_n622), .B(KEYINPUT98), .Z(new_n623));
  INV_X1    g437(.A(new_n420), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n439), .A2(KEYINPUT20), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n439), .A2(KEYINPUT20), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(KEYINPUT33), .B1(new_n485), .B2(new_n486), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n493), .A2(new_n629), .A3(new_n494), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n628), .A2(new_n630), .A3(G478), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n495), .A2(new_n488), .ZN(new_n632));
  NAND2_X1  g446(.A1(G478), .A2(G902), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n627), .A2(new_n635), .ZN(new_n636));
  AND4_X1   g450(.A1(new_n298), .A2(new_n355), .A3(new_n366), .A4(new_n364), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n366), .B1(new_n369), .B2(new_n364), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n305), .B(new_n504), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n623), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT34), .B(G104), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  INV_X1    g456(.A(new_n497), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n420), .B(KEYINPUT99), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n438), .A2(new_n440), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n623), .A2(new_n639), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT35), .B(G107), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  INV_X1    g463(.A(new_n620), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n597), .A2(new_n602), .A3(KEYINPUT82), .ZN(new_n651));
  AOI21_X1  g465(.A(KEYINPUT82), .B1(new_n597), .B2(new_n602), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n564), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(KEYINPUT36), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(new_n589), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n609), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n542), .A2(new_n650), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT100), .B(KEYINPUT37), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G110), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n659), .B(new_n661), .ZN(G12));
  XNOR2_X1  g476(.A(KEYINPUT101), .B(G900), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n499), .B1(new_n501), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n643), .A2(new_n644), .A3(new_n645), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT102), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n371), .A2(new_n541), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n667), .A2(new_n304), .A3(new_n668), .A4(new_n658), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n671));
  INV_X1    g485(.A(G472), .ZN(new_n672));
  INV_X1    g486(.A(new_n276), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n272), .B1(new_n261), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n672), .B1(new_n674), .B2(new_n298), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n188), .B1(new_n618), .B2(new_n190), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n285), .A2(KEYINPUT72), .A3(new_n189), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n675), .B1(new_n678), .B2(new_n187), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n671), .B1(new_n679), .B2(new_n301), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT32), .B1(new_n676), .B2(new_n677), .ZN(new_n681));
  INV_X1    g495(.A(new_n301), .ZN(new_n682));
  NOR4_X1   g496(.A1(new_n681), .A2(KEYINPUT104), .A3(new_n682), .A4(new_n675), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n684), .A2(new_n306), .A3(new_n658), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n368), .A2(new_n370), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT103), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT38), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n441), .A2(new_n497), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n664), .B(KEYINPUT39), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n540), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT40), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n685), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G143), .ZN(G45));
  NOR2_X1   g510(.A1(new_n636), .A2(new_n664), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n304), .A2(new_n668), .A3(new_n658), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  NOR2_X1   g513(.A1(new_n639), .A2(new_n636), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n525), .A2(new_n528), .ZN(new_n701));
  OAI21_X1  g515(.A(G469), .B1(new_n701), .B2(G902), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n529), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n538), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n304), .A2(new_n700), .A3(new_n612), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT41), .B(G113), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G15));
  NOR2_X1   g521(.A1(new_n639), .A2(new_n646), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n304), .A2(new_n612), .A3(new_n708), .A4(new_n704), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G116), .ZN(G18));
  AND2_X1   g524(.A1(new_n371), .A2(new_n704), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n304), .A2(new_n505), .A3(new_n658), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  NAND2_X1  g527(.A1(new_n295), .A2(new_n296), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n290), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n190), .B1(new_n715), .B2(new_n273), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n619), .A2(new_n717), .ZN(new_n718));
  OAI211_X1 g532(.A(KEYINPUT105), .B(G472), .C1(new_n618), .C2(G902), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n716), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n639), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n689), .A2(new_n704), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n720), .A2(new_n721), .A3(new_n612), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G122), .ZN(G24));
  NAND4_X1  g538(.A1(new_n720), .A2(new_n711), .A3(new_n658), .A4(new_n697), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G125), .ZN(G27));
  NOR2_X1   g540(.A1(new_n686), .A2(new_n306), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n612), .B(new_n727), .C1(new_n681), .C2(new_n302), .ZN(new_n728));
  INV_X1    g542(.A(new_n697), .ZN(new_n729));
  NOR4_X1   g543(.A1(new_n728), .A2(KEYINPUT42), .A3(new_n540), .A4(new_n729), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n636), .A2(new_n540), .A3(new_n664), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n187), .B1(new_n618), .B2(new_n190), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n300), .A3(new_n301), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n612), .A2(new_n727), .A3(new_n731), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT42), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n730), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G131), .ZN(G33));
  AOI21_X1  g552(.A(new_n611), .B1(new_n287), .B2(new_n303), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n667), .A2(new_n739), .A3(new_n541), .A4(new_n727), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G134), .ZN(G36));
  NAND2_X1  g555(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n627), .A2(new_n634), .ZN(new_n744));
  MUX2_X1   g558(.A(new_n742), .B(new_n743), .S(new_n744), .Z(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n620), .A3(new_n658), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n747), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n727), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT109), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n533), .A2(new_n534), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(G469), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT106), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n753), .A2(KEYINPUT106), .A3(G469), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(KEYINPUT46), .A3(new_n530), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT107), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n530), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT46), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT107), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n758), .A2(new_n764), .A3(KEYINPUT46), .A4(new_n530), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n760), .A2(new_n763), .A3(new_n529), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n539), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n692), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n748), .A2(new_n769), .A3(new_n727), .A4(new_n749), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n751), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n767), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n766), .A2(KEYINPUT47), .A3(new_n539), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n304), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n727), .A2(new_n611), .A3(new_n697), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G140), .ZN(G42));
  OAI21_X1  g593(.A(new_n688), .B1(KEYINPUT49), .B2(new_n703), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n780), .A2(new_n306), .A3(new_n538), .ZN(new_n781));
  AOI211_X1 g595(.A(new_n683), .B(new_n680), .C1(KEYINPUT49), .C2(new_n703), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n781), .A2(new_n612), .A3(new_n744), .A4(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n745), .A2(new_n499), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n784), .A2(new_n612), .A3(new_n720), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n704), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n688), .A2(new_n306), .ZN(new_n787));
  OAI21_X1  g601(.A(KEYINPUT115), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT50), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n790));
  OAI211_X1 g604(.A(KEYINPUT115), .B(new_n790), .C1(new_n786), .C2(new_n787), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n727), .A2(new_n704), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n784), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n658), .A3(new_n720), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT116), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n774), .B(new_n775), .C1(new_n539), .C2(new_n703), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n727), .A3(new_n785), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n792), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n611), .A2(new_n500), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n684), .A2(new_n793), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n627), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n634), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT117), .ZN(new_n805));
  OR3_X1    g619(.A1(new_n799), .A2(new_n800), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n800), .B1(new_n799), .B2(new_n805), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n653), .A2(new_n657), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n665), .A2(KEYINPUT111), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n540), .B1(new_n813), .B2(new_n664), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n811), .A2(KEYINPUT112), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n371), .A2(new_n689), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n653), .A2(new_n657), .A3(new_n812), .A4(new_n814), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT112), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n815), .B(new_n819), .C1(new_n680), .C2(new_n683), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n669), .A2(new_n698), .A3(new_n725), .ZN(new_n822));
  OAI21_X1  g636(.A(KEYINPUT52), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n669), .A2(new_n698), .A3(new_n725), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT52), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(new_n825), .A3(new_n820), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT42), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n739), .A2(new_n828), .A3(new_n541), .A4(new_n727), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n740), .B(new_n735), .C1(new_n829), .C2(new_n729), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n705), .A2(new_n709), .A3(new_n712), .A4(new_n723), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT110), .B1(new_n627), .B2(new_n497), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n636), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n441), .A2(new_n634), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT110), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n639), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n621), .A2(new_n837), .A3(new_n541), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n613), .A3(new_n659), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n832), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n720), .A2(new_n731), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n541), .B(new_n665), .C1(new_n681), .C2(new_n302), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n644), .A2(new_n497), .A3(new_n645), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(new_n658), .A3(new_n727), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n831), .A2(new_n840), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n810), .B1(new_n827), .B2(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n838), .A2(new_n613), .A3(new_n659), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n709), .A2(new_n723), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n705), .A2(new_n712), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n845), .A2(new_n848), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(new_n830), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(KEYINPUT53), .A3(new_n823), .A4(new_n826), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n847), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n827), .A2(new_n846), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(KEYINPUT114), .A3(KEYINPUT53), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n856), .A2(new_n810), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT53), .B1(new_n827), .B2(new_n846), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n862), .A3(KEYINPUT54), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n785), .A2(new_n711), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n498), .A2(G953), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n865), .B(new_n866), .C1(new_n636), .C2(new_n802), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n611), .B1(new_n303), .B2(new_n732), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n794), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n794), .A2(KEYINPUT118), .A3(new_n869), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(KEYINPUT48), .A3(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n868), .B(new_n874), .C1(KEYINPUT48), .C2(new_n872), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT119), .Z(new_n876));
  NOR3_X1   g690(.A1(new_n808), .A2(new_n864), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(G952), .A2(G953), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n783), .B1(new_n877), .B2(new_n878), .ZN(G75));
  INV_X1    g693(.A(new_n858), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(G210), .A3(G902), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT121), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n348), .B(new_n354), .ZN(new_n883));
  XOR2_X1   g697(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n884));
  XNOR2_X1  g698(.A(new_n883), .B(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n882), .A2(new_n885), .B1(new_n886), .B2(new_n881), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n888));
  AND4_X1   g702(.A1(new_n888), .A2(new_n881), .A3(new_n886), .A4(new_n885), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n258), .A2(G952), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(G51));
  NOR3_X1   g705(.A1(new_n858), .A2(new_n298), .A3(new_n758), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n530), .B(KEYINPUT57), .Z(new_n893));
  AND3_X1   g707(.A1(new_n855), .A2(KEYINPUT54), .A3(new_n857), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT54), .B1(new_n855), .B2(new_n857), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n701), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n892), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT122), .B1(new_n898), .B2(new_n890), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n900));
  INV_X1    g714(.A(new_n890), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n855), .A2(KEYINPUT54), .A3(new_n857), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n860), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n701), .B1(new_n903), .B2(new_n893), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n900), .B(new_n901), .C1(new_n904), .C2(new_n892), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n899), .A2(new_n905), .ZN(G54));
  NAND4_X1  g720(.A1(new_n880), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n907));
  INV_X1    g721(.A(new_n436), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n907), .A2(new_n908), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n909), .A2(new_n910), .A3(new_n890), .ZN(G60));
  NAND2_X1  g725(.A1(new_n628), .A2(new_n630), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n633), .B(KEYINPUT59), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n903), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n912), .B1(new_n864), .B2(new_n913), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n914), .A2(new_n915), .A3(new_n890), .ZN(G63));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT60), .Z(new_n918));
  AOI21_X1  g732(.A(new_n608), .B1(new_n880), .B2(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n855), .A2(new_n857), .A3(new_n656), .A4(new_n918), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n901), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT61), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n923), .A2(KEYINPUT61), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n922), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n923), .B(KEYINPUT61), .C1(new_n919), .C2(new_n921), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(G66));
  AOI21_X1  g742(.A(new_n352), .B1(new_n503), .B2(G224), .ZN(new_n929));
  INV_X1    g743(.A(new_n840), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n929), .B1(new_n930), .B2(new_n258), .ZN(new_n931));
  INV_X1    g745(.A(G898), .ZN(new_n932));
  INV_X1    g746(.A(new_n258), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n348), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT124), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n931), .B(new_n935), .ZN(G69));
  XNOR2_X1  g750(.A(new_n254), .B(new_n427), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n933), .A2(G900), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n822), .B1(new_n776), .B2(new_n777), .ZN(new_n939));
  INV_X1    g753(.A(new_n816), .ZN(new_n940));
  AOI22_X1  g754(.A1(new_n751), .A2(new_n770), .B1(new_n869), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n768), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n939), .B(new_n831), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n937), .B(new_n938), .C1(new_n943), .C2(new_n933), .ZN(new_n944));
  NAND2_X1  g758(.A1(G227), .A2(G900), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n933), .A2(new_n945), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT126), .Z(new_n947));
  NAND2_X1  g761(.A1(new_n834), .A2(new_n836), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n739), .A2(new_n693), .A3(new_n727), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n771), .A2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n771), .A2(KEYINPUT125), .A3(new_n949), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n695), .A2(new_n824), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT62), .Z(new_n956));
  NAND3_X1  g770(.A1(new_n954), .A2(new_n778), .A3(new_n956), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n957), .A2(new_n258), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n944), .B(new_n947), .C1(new_n958), .C2(new_n937), .ZN(new_n959));
  INV_X1    g773(.A(new_n947), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n937), .B1(new_n957), .B2(new_n258), .ZN(new_n961));
  INV_X1    g775(.A(new_n944), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n959), .A2(new_n963), .ZN(G72));
  NAND4_X1  g778(.A1(new_n954), .A2(new_n778), .A3(new_n840), .A4(new_n956), .ZN(new_n965));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  AOI211_X1 g781(.A(new_n290), .B(new_n255), .C1(new_n965), .C2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n943), .B2(new_n930), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n969), .A2(new_n290), .A3(new_n255), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n272), .A2(new_n291), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n861), .A2(new_n862), .A3(new_n967), .A4(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n970), .A2(new_n901), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(KEYINPUT127), .B1(new_n968), .B2(new_n973), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n970), .A2(new_n901), .A3(new_n972), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n965), .A2(new_n967), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n976), .A2(new_n261), .A3(new_n289), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n975), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n974), .A2(new_n979), .ZN(G57));
endmodule


