//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n801, new_n803, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1027, new_n1028, new_n1029;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT11), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G197gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209));
  INV_X1    g008(.A(G43gat), .ZN(new_n210));
  INV_X1    g009(.A(G50gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G43gat), .A2(G50gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT14), .ZN(new_n215));
  INV_X1    g014(.A(G29gat), .ZN(new_n216));
  INV_X1    g015(.A(G36gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n218), .A2(new_n219), .B1(G29gat), .B2(G36gat), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n214), .B1(new_n220), .B2(KEYINPUT88), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n212), .A2(new_n209), .A3(new_n213), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n220), .B(new_n222), .C1(new_n214), .C2(KEYINPUT88), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G15gat), .B(G22gat), .ZN(new_n227));
  INV_X1    g026(.A(G1gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(KEYINPUT16), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(new_n228), .B2(new_n227), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G8gat), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n230), .A2(G8gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n226), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n231), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n224), .A2(new_n225), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238));
  XOR2_X1   g037(.A(new_n238), .B(KEYINPUT13), .Z(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT91), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n237), .A2(KEYINPUT91), .A3(new_n239), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT17), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n235), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT17), .B1(new_n224), .B2(new_n225), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n234), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n248), .A2(KEYINPUT18), .A3(new_n238), .A4(new_n233), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT90), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n249), .A2(new_n250), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n244), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n248), .A2(new_n233), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT89), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n254), .A2(new_n255), .A3(new_n238), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n248), .A2(new_n238), .A3(new_n233), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT89), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT18), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n208), .B1(new_n253), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT18), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n257), .A2(KEYINPUT89), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n257), .A2(KEYINPUT89), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n249), .B(new_n250), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n264), .A2(new_n265), .A3(new_n244), .A4(new_n207), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G183gat), .B(G211gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT94), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G127gat), .B(G155gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n271), .B(KEYINPUT93), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(G57gat), .B(G64gat), .Z(new_n274));
  INV_X1    g073(.A(KEYINPUT9), .ZN(new_n275));
  INV_X1    g074(.A(G71gat), .ZN(new_n276));
  INV_X1    g075(.A(G78gat), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G71gat), .B(G78gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n274), .A2(new_n280), .A3(new_n278), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT92), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT21), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n285), .B1(new_n284), .B2(new_n286), .ZN(new_n289));
  INV_X1    g088(.A(G231gat), .ZN(new_n290));
  INV_X1    g089(.A(G233gat), .ZN(new_n291));
  OAI22_X1  g090(.A1(new_n288), .A2(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n284), .A2(new_n286), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT92), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n290), .A2(new_n291), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(new_n295), .A3(new_n287), .ZN(new_n296));
  XOR2_X1   g095(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n297));
  NAND3_X1  g096(.A1(new_n292), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n297), .B1(new_n292), .B2(new_n296), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n273), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n300), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n302), .A2(new_n272), .A3(new_n298), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n234), .B1(new_n286), .B2(new_n284), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n304), .B1(new_n301), .B2(new_n303), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n270), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n304), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n272), .B1(new_n302), .B2(new_n298), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n299), .A2(new_n300), .A3(new_n273), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(new_n312), .A3(new_n269), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  AND2_X1   g114(.A1(G232gat), .A2(G233gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n316), .A2(KEYINPUT41), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT95), .ZN(new_n318));
  XNOR2_X1  g117(.A(G134gat), .B(G162gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT96), .B(G92gat), .ZN(new_n321));
  INV_X1    g120(.A(G85gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(G99gat), .A2(G106gat), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n325), .B1(KEYINPUT8), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n323), .A2(new_n324), .A3(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(G99gat), .B(G106gat), .Z(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n329), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n331), .A2(new_n323), .A3(new_n324), .A4(new_n327), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n333), .B1(new_n246), .B2(new_n247), .ZN(new_n334));
  INV_X1    g133(.A(new_n333), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n226), .A2(new_n335), .B1(KEYINPUT41), .B2(new_n316), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G190gat), .B(G218gat), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n338), .B(KEYINPUT97), .Z(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n334), .A2(new_n339), .A3(new_n336), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n320), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT98), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n343), .A2(new_n344), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n341), .A2(new_n342), .A3(new_n320), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT99), .ZN(new_n349));
  OR2_X1    g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n349), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT10), .ZN(new_n355));
  OR3_X1    g154(.A1(new_n333), .A2(new_n355), .A3(new_n284), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT101), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT100), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n282), .A2(new_n358), .A3(new_n283), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n333), .ZN(new_n361));
  INV_X1    g160(.A(new_n283), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n280), .B1(new_n274), .B2(new_n278), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT100), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n364), .A2(new_n359), .A3(new_n332), .A4(new_n330), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n357), .B1(new_n366), .B2(new_n355), .ZN(new_n367));
  AOI211_X1 g166(.A(KEYINPUT101), .B(KEYINPUT10), .C1(new_n361), .C2(new_n365), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n356), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G230gat), .A2(G233gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n370), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n361), .A2(new_n365), .A3(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G120gat), .B(G148gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(G176gat), .B(G204gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n371), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n377), .B1(new_n371), .B2(new_n373), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NOR3_X1   g181(.A1(new_n315), .A2(new_n354), .A3(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G78gat), .B(G106gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT29), .ZN(new_n386));
  OR3_X1    g185(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(G155gat), .A2(G162gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G141gat), .A2(G148gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(G141gat), .A2(G148gat), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT76), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(G141gat), .ZN(new_n395));
  INV_X1    g194(.A(G148gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT76), .B1(new_n397), .B2(new_n390), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n389), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n388), .ZN(new_n401));
  NOR3_X1   g200(.A1(KEYINPUT75), .A2(G155gat), .A3(G162gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT2), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n397), .A2(new_n404), .A3(new_n390), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n399), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n386), .B1(new_n407), .B2(KEYINPUT3), .ZN(new_n408));
  NAND2_X1  g207(.A1(G211gat), .A2(G218gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(G211gat), .A2(G218gat), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(G204gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(G197gat), .ZN(new_n415));
  INV_X1    g214(.A(G197gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(G204gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n418), .A2(KEYINPUT70), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT70), .ZN(new_n421));
  XNOR2_X1  g220(.A(G197gat), .B(G204gat), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT22), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n409), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n421), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n413), .B1(new_n420), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT70), .B1(new_n418), .B2(new_n419), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n422), .A2(new_n421), .A3(new_n424), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n412), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n408), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n426), .A2(new_n386), .A3(new_n429), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT82), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n426), .A2(KEYINPUT82), .A3(new_n386), .A4(new_n429), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT3), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n393), .B1(new_n391), .B2(new_n392), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n397), .A2(KEYINPUT76), .A3(new_n390), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n439), .A2(new_n389), .B1(new_n403), .B2(new_n405), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n431), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G228gat), .A2(G233gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(G22gat), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT3), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n432), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n442), .B1(new_n446), .B2(new_n407), .ZN(new_n447));
  XOR2_X1   g246(.A(new_n430), .B(KEYINPUT71), .Z(new_n448));
  INV_X1    g247(.A(KEYINPUT83), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n408), .B(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n447), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n443), .A2(new_n444), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n444), .B1(new_n443), .B2(new_n451), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n385), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n443), .A2(new_n451), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(G22gat), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n443), .A2(new_n444), .A3(new_n451), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(new_n384), .ZN(new_n458));
  XOR2_X1   g257(.A(KEYINPUT31), .B(G50gat), .Z(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n454), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n460), .B1(new_n454), .B2(new_n458), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(G183gat), .ZN(new_n464));
  INV_X1    g263(.A(G190gat), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT24), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT24), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n467), .A2(G183gat), .A3(G190gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n469), .B1(G183gat), .B2(G190gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(G169gat), .A2(G176gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT23), .ZN(new_n472));
  INV_X1    g271(.A(G176gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n204), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(G169gat), .A2(G176gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT23), .ZN(new_n477));
  NOR2_X1   g276(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n475), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT64), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n480), .B1(new_n475), .B2(new_n477), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n470), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT26), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n471), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n474), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n476), .A2(new_n483), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n485), .A2(new_n486), .B1(G183gat), .B2(G190gat), .ZN(new_n487));
  AND2_X1   g286(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n488));
  NOR2_X1   g287(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(KEYINPUT27), .B(G183gat), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT28), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT28), .B1(new_n490), .B2(new_n491), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n487), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n490), .A2(new_n464), .B1(new_n466), .B2(new_n468), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n475), .A2(new_n477), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT25), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n482), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(G134gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT66), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT66), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(G134gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(new_n502), .A3(G127gat), .ZN(new_n503));
  INV_X1    g302(.A(G127gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT67), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT67), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(G127gat), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n507), .A3(G134gat), .ZN(new_n508));
  INV_X1    g307(.A(G120gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(G113gat), .ZN(new_n510));
  INV_X1    g309(.A(G113gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(G120gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT1), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n503), .A2(new_n508), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G127gat), .B(G134gat), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n513), .A2(new_n516), .A3(new_n514), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n498), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G227gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n520), .A2(new_n291), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n508), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n513), .A2(new_n514), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n513), .A2(new_n516), .A3(new_n514), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n482), .A2(new_n526), .A3(new_n494), .A4(new_n497), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n519), .A2(new_n521), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT33), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT68), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT68), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n528), .A2(new_n532), .A3(new_n529), .ZN(new_n533));
  XOR2_X1   g332(.A(G15gat), .B(G43gat), .Z(new_n534));
  XNOR2_X1  g333(.A(G71gat), .B(G99gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n537), .B1(new_n528), .B2(KEYINPUT32), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n531), .A2(new_n533), .A3(new_n538), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n528), .B(KEYINPUT32), .C1(new_n529), .C2(new_n537), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n519), .A2(new_n527), .ZN(new_n543));
  INV_X1    g342(.A(new_n521), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n545), .A2(KEYINPUT34), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(KEYINPUT34), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT69), .B1(new_n542), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n548), .B1(new_n539), .B2(new_n540), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT69), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n542), .A2(new_n548), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n549), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n463), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT5), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n524), .A2(new_n399), .A3(new_n406), .A4(new_n525), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT78), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n518), .A2(new_n440), .A3(KEYINPUT78), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n526), .A2(new_n407), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G225gat), .A2(G233gat), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n556), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT4), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n559), .A2(new_n566), .A3(new_n560), .ZN(new_n567));
  AND4_X1   g366(.A1(new_n406), .A2(new_n524), .A3(new_n399), .A4(new_n525), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n564), .B1(new_n568), .B2(KEYINPUT4), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n440), .A2(new_n445), .B1(new_n524), .B2(new_n525), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT77), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n571), .B1(new_n440), .B2(new_n445), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n407), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n567), .A2(new_n569), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n565), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n560), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT4), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n557), .A2(new_n566), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n564), .A2(KEYINPUT5), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n578), .A2(new_n574), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G1gat), .B(G29gat), .Z(new_n583));
  XNOR2_X1  g382(.A(G57gat), .B(G85gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n585), .B(new_n586), .Z(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT85), .ZN(new_n590));
  XOR2_X1   g389(.A(KEYINPUT80), .B(KEYINPUT6), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n579), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n566), .B1(new_n559), .B2(new_n560), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n595), .A2(new_n580), .B1(new_n575), .B2(new_n565), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n592), .B1(new_n596), .B2(new_n587), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT85), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n598), .A3(new_n588), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n590), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n582), .A2(new_n588), .A3(new_n592), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT35), .ZN(new_n603));
  INV_X1    g402(.A(G226gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n604), .A2(new_n291), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n498), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n605), .B1(new_n498), .B2(new_n386), .ZN(new_n608));
  NOR3_X1   g407(.A1(new_n607), .A2(new_n608), .A3(new_n430), .ZN(new_n609));
  INV_X1    g408(.A(new_n608), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT72), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n611), .B1(new_n498), .B2(new_n605), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n498), .A2(new_n611), .A3(new_n605), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n610), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n448), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n609), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT30), .ZN(new_n618));
  XNOR2_X1  g417(.A(G8gat), .B(G36gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT73), .ZN(new_n620));
  XNOR2_X1  g419(.A(G64gat), .B(G92gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n617), .A2(new_n618), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n622), .B(KEYINPUT74), .Z(new_n625));
  OAI21_X1  g424(.A(KEYINPUT30), .B1(new_n617), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n610), .A2(new_n429), .A3(new_n426), .A4(new_n606), .ZN(new_n627));
  INV_X1    g426(.A(new_n614), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n628), .A2(new_n608), .A3(new_n612), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n627), .B1(new_n629), .B2(new_n448), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n630), .A2(new_n622), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n624), .B1(new_n626), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n602), .A2(new_n603), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n555), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT87), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n452), .A2(new_n453), .A3(new_n385), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n384), .B1(new_n456), .B2(new_n457), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n459), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n454), .A2(new_n458), .A3(new_n460), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n541), .A2(new_n546), .A3(new_n547), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(new_n550), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n635), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n463), .A2(KEYINPUT87), .A3(new_n642), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n576), .A2(new_n587), .A3(new_n581), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n589), .A2(KEYINPUT81), .A3(new_n646), .A4(new_n591), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n601), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT81), .B1(new_n597), .B2(new_n589), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n632), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n644), .A2(new_n645), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n634), .B1(new_n652), .B2(KEYINPUT35), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n650), .B1(new_n639), .B2(new_n638), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n608), .A2(new_n612), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n448), .B1(new_n655), .B2(new_n614), .ZN(new_n656));
  OAI21_X1  g455(.A(KEYINPUT37), .B1(new_n656), .B2(new_n609), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT37), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n627), .B(new_n658), .C1(new_n629), .C2(new_n448), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n657), .A2(new_n622), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n631), .B1(new_n660), .B2(KEYINPUT38), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n430), .B1(new_n607), .B2(new_n608), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n615), .B2(new_n616), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(KEYINPUT37), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT86), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n625), .A2(KEYINPUT38), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n659), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n663), .A2(KEYINPUT86), .A3(KEYINPUT37), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n666), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n661), .A2(new_n670), .A3(new_n601), .A4(new_n600), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n630), .A2(KEYINPUT30), .A3(new_n622), .ZN(new_n672));
  INV_X1    g471(.A(new_n625), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n618), .B1(new_n630), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n617), .A2(new_n623), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n590), .A2(new_n599), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n562), .A2(new_n564), .ZN(new_n678));
  OAI211_X1 g477(.A(KEYINPUT39), .B(new_n678), .C1(new_n595), .C2(new_n563), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT39), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n680), .B(new_n564), .C1(new_n593), .C2(new_n594), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT84), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n681), .A2(new_n682), .A3(new_n587), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n682), .B1(new_n681), .B2(new_n587), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n679), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n679), .B(KEYINPUT40), .C1(new_n683), .C2(new_n684), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n676), .A2(new_n677), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n671), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n654), .B1(new_n463), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT36), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n641), .A2(new_n550), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n549), .A2(new_n552), .A3(new_n553), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n694), .B2(new_n692), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n267), .B(new_n383), .C1(new_n653), .C2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n648), .A2(new_n649), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(new_n228), .ZN(G1324gat));
  NOR2_X1   g500(.A1(new_n697), .A2(new_n632), .ZN(new_n702));
  XOR2_X1   g501(.A(KEYINPUT16), .B(G8gat), .Z(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n702), .A2(KEYINPUT42), .A3(new_n703), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n702), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT102), .B1(new_n709), .B2(G8gat), .ZN(new_n710));
  OAI211_X1 g509(.A(KEYINPUT102), .B(G8gat), .C1(new_n697), .C2(new_n632), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n708), .B(KEYINPUT103), .C1(new_n710), .C2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n710), .A2(new_n712), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n706), .A2(new_n707), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n713), .A2(new_n717), .ZN(G1325gat));
  INV_X1    g517(.A(new_n693), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n554), .B2(KEYINPUT36), .ZN(new_n720));
  OAI21_X1  g519(.A(G15gat), .B1(new_n697), .B2(new_n720), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n694), .A2(G15gat), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n697), .B2(new_n722), .ZN(G1326gat));
  NOR2_X1   g522(.A1(new_n697), .A2(new_n463), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT104), .ZN(new_n725));
  XNOR2_X1  g524(.A(KEYINPUT43), .B(G22gat), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1327gat));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n691), .B2(new_n695), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n690), .A2(new_n463), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n640), .A2(new_n651), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n732), .A2(KEYINPUT106), .A3(new_n720), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(KEYINPUT107), .B1(new_n734), .B2(new_n653), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n652), .A2(KEYINPUT35), .ZN(new_n736));
  INV_X1    g535(.A(new_n634), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n738), .A2(new_n739), .A3(new_n733), .A4(new_n729), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n353), .A2(KEYINPUT44), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n735), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n653), .A2(new_n696), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT44), .B1(new_n743), .B2(new_n353), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n314), .A2(KEYINPUT105), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT105), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n307), .B2(new_n313), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n267), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n749), .A2(new_n750), .A3(new_n382), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n745), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G29gat), .B1(new_n752), .B2(new_n699), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n743), .A2(new_n750), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n314), .A2(new_n382), .A3(new_n353), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n756), .A2(G29gat), .A3(new_n699), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n757), .A2(KEYINPUT45), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(KEYINPUT45), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n753), .A2(new_n758), .A3(new_n759), .ZN(G1328gat));
  OAI21_X1  g559(.A(G36gat), .B1(new_n752), .B2(new_n632), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n632), .A2(G36gat), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n756), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n754), .A2(KEYINPUT108), .A3(new_n755), .A4(new_n763), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n765), .A2(KEYINPUT46), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT46), .B1(new_n765), .B2(new_n766), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n761), .B1(new_n767), .B2(new_n768), .ZN(G1329gat));
  OAI21_X1  g568(.A(new_n210), .B1(new_n756), .B2(new_n694), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n720), .A2(new_n210), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n770), .B1(new_n752), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT47), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT47), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n775), .B(new_n770), .C1(new_n752), .C2(new_n772), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(G1330gat));
  OAI21_X1  g576(.A(G50gat), .B1(new_n752), .B2(new_n463), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n463), .A2(G50gat), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT109), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n756), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n778), .A2(KEYINPUT48), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT48), .ZN(new_n784));
  INV_X1    g583(.A(new_n751), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n742), .B2(new_n744), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n211), .B1(new_n786), .B2(new_n640), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n784), .B1(new_n787), .B2(new_n781), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n783), .A2(new_n788), .ZN(G1331gat));
  NOR4_X1   g588(.A1(new_n315), .A2(new_n354), .A3(new_n267), .A4(new_n381), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n735), .A2(new_n740), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(new_n699), .ZN(new_n792));
  XOR2_X1   g591(.A(new_n792), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g592(.A1(new_n791), .A2(new_n632), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n794), .A2(KEYINPUT49), .A3(G64gat), .ZN(new_n795));
  XOR2_X1   g594(.A(KEYINPUT49), .B(G64gat), .Z(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n794), .B2(new_n796), .ZN(G1333gat));
  OAI21_X1  g596(.A(G71gat), .B1(new_n791), .B2(new_n720), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n554), .A2(new_n276), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n791), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n800), .B(new_n801), .ZN(G1334gat));
  NOR2_X1   g601(.A1(new_n791), .A2(new_n463), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(new_n277), .ZN(G1335gat));
  NOR2_X1   g603(.A1(new_n314), .A2(new_n267), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n382), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n742), .B2(new_n744), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(G85gat), .B1(new_n808), .B2(new_n699), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n805), .A2(new_n354), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  OAI211_X1 g610(.A(KEYINPUT51), .B(new_n811), .C1(new_n734), .C2(new_n653), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT110), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n738), .A2(new_n733), .A3(new_n729), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT110), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n814), .A2(new_n815), .A3(KEYINPUT51), .A4(new_n811), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT106), .B1(new_n732), .B2(new_n720), .ZN(new_n818));
  AOI211_X1 g617(.A(new_n728), .B(new_n695), .C1(new_n730), .C2(new_n731), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n653), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n817), .B1(new_n820), .B2(new_n810), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n813), .A2(new_n816), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n382), .A2(new_n322), .A3(new_n698), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n809), .B1(new_n823), .B2(new_n824), .ZN(G1336gat));
  AOI21_X1  g624(.A(new_n321), .B1(new_n807), .B2(new_n676), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n381), .A2(G92gat), .A3(new_n632), .ZN(new_n827));
  XOR2_X1   g626(.A(new_n827), .B(KEYINPUT111), .Z(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n821), .B2(new_n812), .ZN(new_n829));
  OAI21_X1  g628(.A(KEYINPUT52), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT112), .ZN(new_n831));
  INV_X1    g630(.A(new_n828), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n822), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n831), .B1(new_n822), .B2(new_n832), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n836));
  AOI211_X1 g635(.A(new_n632), .B(new_n806), .C1(new_n742), .C2(new_n744), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(new_n321), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n830), .B1(new_n835), .B2(new_n838), .ZN(G1337gat));
  OAI21_X1  g638(.A(G99gat), .B1(new_n808), .B2(new_n720), .ZN(new_n840));
  OR3_X1    g639(.A1(new_n694), .A2(G99gat), .A3(new_n381), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n840), .B1(new_n823), .B2(new_n841), .ZN(G1338gat));
  INV_X1    g641(.A(G106gat), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n843), .B1(new_n807), .B2(new_n640), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n821), .A2(new_n812), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n463), .A2(G106gat), .A3(new_n381), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT53), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n822), .A2(new_n846), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n848), .B1(new_n844), .B2(new_n851), .ZN(G1339gat));
  OR2_X1    g651(.A1(new_n746), .A2(new_n748), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n356), .B(new_n372), .C1(new_n367), .C2(new_n368), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n371), .A2(KEYINPUT54), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n369), .A2(new_n856), .A3(new_n370), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n855), .A2(KEYINPUT55), .A3(new_n376), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n378), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n376), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT55), .B1(new_n861), .B2(new_n855), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n237), .A2(new_n239), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT113), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n254), .A2(new_n238), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n206), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n266), .A2(new_n866), .ZN(new_n867));
  NOR4_X1   g666(.A1(new_n353), .A2(new_n859), .A3(new_n862), .A4(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT55), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n371), .A2(KEYINPUT54), .A3(new_n854), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(new_n860), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n267), .A2(new_n871), .A3(new_n378), .A4(new_n858), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n266), .B(new_n866), .C1(new_n379), .C2(new_n380), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n354), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n853), .B1(new_n868), .B2(new_n874), .ZN(new_n875));
  NOR4_X1   g674(.A1(new_n315), .A2(new_n354), .A3(new_n267), .A4(new_n382), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n699), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n878), .A2(new_n632), .ZN(new_n879));
  INV_X1    g678(.A(new_n555), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n881), .A2(new_n511), .A3(new_n750), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n644), .A2(new_n645), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  XOR2_X1   g683(.A(new_n884), .B(KEYINPUT114), .Z(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(new_n632), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n267), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n882), .B1(new_n887), .B2(new_n511), .ZN(G1340gat));
  NOR2_X1   g687(.A1(new_n381), .A2(G120gat), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT115), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(G120gat), .B1(new_n881), .B2(new_n381), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(G1341gat));
  NAND2_X1  g692(.A1(new_n886), .A2(new_n314), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n505), .A2(new_n507), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n853), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n880), .A3(new_n896), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n897), .A2(KEYINPUT116), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(KEYINPUT116), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n894), .A2(new_n895), .B1(new_n898), .B2(new_n899), .ZN(G1342gat));
  OAI21_X1  g699(.A(G134gat), .B1(new_n881), .B2(new_n353), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n353), .A2(new_n676), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n902), .A2(new_n500), .A3(new_n502), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n885), .A2(KEYINPUT56), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT56), .B1(new_n885), .B2(new_n903), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n901), .B1(new_n904), .B2(new_n905), .ZN(G1343gat));
  NOR2_X1   g705(.A1(new_n750), .A2(G141gat), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n720), .A2(new_n640), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n908), .B(KEYINPUT119), .Z(new_n909));
  NAND3_X1  g708(.A1(new_n879), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT57), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n872), .A2(new_n873), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n353), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n859), .A2(new_n862), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n914), .A2(new_n354), .A3(new_n266), .A4(new_n866), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n749), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n911), .B(new_n640), .C1(new_n916), .C2(new_n876), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n695), .A2(new_n699), .A3(new_n676), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT117), .B1(new_n859), .B2(new_n862), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT117), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n871), .A2(new_n921), .A3(new_n378), .A4(new_n858), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n750), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(new_n873), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n353), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n314), .B1(new_n925), .B2(new_n915), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n640), .B1(new_n926), .B2(new_n876), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n919), .B1(new_n927), .B2(KEYINPUT57), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n395), .B1(new_n928), .B2(new_n267), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT118), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n910), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI211_X1 g730(.A(KEYINPUT118), .B(new_n395), .C1(new_n928), .C2(new_n267), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT58), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n909), .A2(new_n878), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(KEYINPUT120), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT120), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n909), .A2(new_n936), .A3(new_n878), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n676), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(KEYINPUT58), .B1(new_n938), .B2(new_n907), .ZN(new_n939));
  INV_X1    g738(.A(new_n929), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n933), .A2(new_n941), .ZN(G1344gat));
  NAND3_X1  g741(.A1(new_n938), .A2(new_n396), .A3(new_n382), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT59), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT121), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n925), .A2(new_n915), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n945), .B(new_n877), .C1(new_n946), .C2(new_n314), .ZN(new_n947));
  OAI21_X1  g746(.A(KEYINPUT121), .B1(new_n926), .B2(new_n876), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n463), .A2(KEYINPUT57), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n875), .A2(new_n877), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(new_n640), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(KEYINPUT57), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n950), .A2(new_n382), .A3(new_n918), .A4(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n944), .B1(new_n954), .B2(G148gat), .ZN(new_n955));
  AOI211_X1 g754(.A(KEYINPUT59), .B(new_n396), .C1(new_n928), .C2(new_n382), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n943), .B1(new_n955), .B2(new_n956), .ZN(G1345gat));
  INV_X1    g756(.A(new_n928), .ZN(new_n958));
  OAI21_X1  g757(.A(G155gat), .B1(new_n958), .B2(new_n853), .ZN(new_n959));
  INV_X1    g758(.A(G155gat), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n938), .A2(new_n960), .A3(new_n314), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT122), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT122), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n959), .A2(new_n961), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(G1346gat));
  OAI21_X1  g765(.A(G162gat), .B1(new_n958), .B2(new_n353), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n935), .A2(new_n937), .ZN(new_n968));
  INV_X1    g767(.A(G162gat), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n968), .A2(new_n969), .A3(new_n902), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n967), .A2(new_n970), .ZN(G1347gat));
  NAND2_X1  g770(.A1(new_n699), .A2(new_n676), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n972), .A2(KEYINPUT123), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n972), .A2(KEYINPUT123), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n973), .A2(new_n974), .A3(new_n555), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n951), .A2(new_n975), .ZN(new_n976));
  NOR3_X1   g775(.A1(new_n976), .A2(new_n204), .A3(new_n750), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n698), .B1(new_n875), .B2(new_n877), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n978), .A2(new_n883), .A3(new_n676), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(new_n267), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n977), .B1(new_n980), .B2(new_n204), .ZN(G1348gat));
  NAND3_X1  g780(.A1(new_n979), .A2(new_n473), .A3(new_n382), .ZN(new_n982));
  OAI21_X1  g781(.A(G176gat), .B1(new_n976), .B2(new_n381), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(G1349gat));
  INV_X1    g783(.A(new_n976), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n464), .B1(new_n985), .B2(new_n749), .ZN(new_n986));
  AND2_X1   g785(.A1(new_n314), .A2(new_n491), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n986), .B1(new_n979), .B2(new_n987), .ZN(new_n988));
  XOR2_X1   g787(.A(new_n988), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g788(.A1(new_n951), .A2(new_n354), .A3(new_n975), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(G190gat), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n991), .A2(KEYINPUT124), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT124), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n990), .A2(new_n993), .A3(G190gat), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT61), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n992), .A2(KEYINPUT61), .A3(new_n994), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n979), .A2(new_n490), .A3(new_n354), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT125), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g801(.A1(new_n997), .A2(KEYINPUT125), .A3(new_n998), .A4(new_n999), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(G1351gat));
  NOR2_X1   g803(.A1(new_n908), .A2(new_n632), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n978), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g805(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g806(.A(G197gat), .B1(new_n1007), .B2(new_n267), .ZN(new_n1008));
  NOR3_X1   g807(.A1(new_n973), .A2(new_n974), .A3(new_n695), .ZN(new_n1009));
  AND3_X1   g808(.A1(new_n950), .A2(new_n953), .A3(new_n1009), .ZN(new_n1010));
  NOR2_X1   g809(.A1(new_n750), .A2(new_n416), .ZN(new_n1011));
  AOI21_X1  g810(.A(new_n1008), .B1(new_n1010), .B2(new_n1011), .ZN(G1352gat));
  NOR3_X1   g811(.A1(new_n1006), .A2(G204gat), .A3(new_n381), .ZN(new_n1013));
  XNOR2_X1  g812(.A(new_n1013), .B(KEYINPUT62), .ZN(new_n1014));
  NAND4_X1  g813(.A1(new_n950), .A2(new_n382), .A3(new_n953), .A4(new_n1009), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1015), .A2(G204gat), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1017), .A2(KEYINPUT126), .ZN(new_n1018));
  INV_X1    g817(.A(KEYINPUT126), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n1014), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1018), .A2(new_n1020), .ZN(G1353gat));
  OR3_X1    g820(.A1(new_n1006), .A2(G211gat), .A3(new_n315), .ZN(new_n1022));
  NAND4_X1  g821(.A1(new_n950), .A2(new_n314), .A3(new_n953), .A4(new_n1009), .ZN(new_n1023));
  AND3_X1   g822(.A1(new_n1023), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1024));
  AOI21_X1  g823(.A(KEYINPUT63), .B1(new_n1023), .B2(G211gat), .ZN(new_n1025));
  OAI21_X1  g824(.A(new_n1022), .B1(new_n1024), .B2(new_n1025), .ZN(G1354gat));
  AOI21_X1  g825(.A(G218gat), .B1(new_n1007), .B2(new_n354), .ZN(new_n1027));
  NAND2_X1  g826(.A1(new_n354), .A2(G218gat), .ZN(new_n1028));
  XNOR2_X1  g827(.A(new_n1028), .B(KEYINPUT127), .ZN(new_n1029));
  AOI21_X1  g828(.A(new_n1027), .B1(new_n1010), .B2(new_n1029), .ZN(G1355gat));
endmodule


