

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754;

  XNOR2_X1 U379 ( .A(n380), .B(n437), .ZN(n374) );
  NOR2_X1 U380 ( .A1(n751), .A2(n753), .ZN(n560) );
  XNOR2_X1 U381 ( .A(G104), .B(G122), .ZN(n381) );
  XNOR2_X1 U382 ( .A(n381), .B(G113), .ZN(n470) );
  INV_X2 U383 ( .A(G953), .ZN(n743) );
  XNOR2_X2 U384 ( .A(n586), .B(n585), .ZN(n594) );
  NOR2_X2 U385 ( .A1(n541), .A2(n550), .ZN(n364) );
  NAND2_X1 U386 ( .A1(n515), .A2(n514), .ZN(n660) );
  NOR2_X2 U387 ( .A1(G953), .A2(G237), .ZN(n424) );
  BUF_X1 U388 ( .A(G128), .Z(n357) );
  AND2_X1 U389 ( .A1(n497), .A2(n496), .ZN(n498) );
  NOR2_X2 U390 ( .A1(n577), .A2(n576), .ZN(n642) );
  XNOR2_X1 U391 ( .A(n478), .B(n477), .ZN(n515) );
  XOR2_X1 U392 ( .A(n634), .B(KEYINPUT122), .Z(n635) );
  XNOR2_X1 U393 ( .A(n376), .B(n375), .ZN(n634) );
  XNOR2_X1 U394 ( .A(n377), .B(n416), .ZN(n376) );
  XNOR2_X1 U395 ( .A(n413), .B(n473), .ZN(n375) );
  XNOR2_X1 U396 ( .A(n383), .B(G119), .ZN(n382) );
  XNOR2_X1 U397 ( .A(KEYINPUT3), .B(KEYINPUT73), .ZN(n428) );
  XNOR2_X1 U398 ( .A(G119), .B(G110), .ZN(n411) );
  BUF_X1 U399 ( .A(n739), .Z(n355) );
  BUF_X1 U400 ( .A(n562), .Z(n356) );
  XNOR2_X1 U401 ( .A(n372), .B(n371), .ZN(n562) );
  BUF_X1 U402 ( .A(n373), .Z(n358) );
  XNOR2_X1 U403 ( .A(n382), .B(n428), .ZN(n373) );
  XNOR2_X2 U404 ( .A(KEYINPUT66), .B(G101), .ZN(n429) );
  XNOR2_X1 U405 ( .A(n642), .B(n366), .ZN(n365) );
  INV_X1 U406 ( .A(KEYINPUT84), .ZN(n366) );
  XNOR2_X1 U407 ( .A(n384), .B(KEYINPUT75), .ZN(n565) );
  XNOR2_X1 U408 ( .A(n364), .B(KEYINPUT78), .ZN(n545) );
  XNOR2_X1 U409 ( .A(n390), .B(n389), .ZN(n514) );
  INV_X1 U410 ( .A(G478), .ZN(n389) );
  OR2_X1 U411 ( .A1(n724), .A2(G902), .ZN(n390) );
  NAND2_X1 U412 ( .A1(n521), .A2(n645), .ZN(n530) );
  AND2_X1 U413 ( .A1(n660), .A2(n663), .ZN(n679) );
  XNOR2_X1 U414 ( .A(G116), .B(G113), .ZN(n422) );
  XNOR2_X1 U415 ( .A(n429), .B(n430), .ZN(n362) );
  NOR2_X1 U416 ( .A1(n581), .A2(n580), .ZN(n582) );
  INV_X1 U417 ( .A(KEYINPUT19), .ZN(n371) );
  XNOR2_X1 U418 ( .A(n429), .B(n397), .ZN(n439) );
  XNOR2_X1 U419 ( .A(KEYINPUT74), .B(G110), .ZN(n397) );
  XNOR2_X1 U420 ( .A(n435), .B(n434), .ZN(n709) );
  NOR2_X1 U421 ( .A1(n660), .A2(n452), .ZN(n379) );
  INV_X1 U422 ( .A(KEYINPUT94), .ZN(n460) );
  NAND2_X1 U423 ( .A1(n612), .A2(n476), .ZN(n432) );
  XNOR2_X1 U424 ( .A(n485), .B(n486), .ZN(n724) );
  NAND2_X1 U425 ( .A1(n561), .A2(n385), .ZN(n384) );
  INV_X1 U426 ( .A(KEYINPUT47), .ZN(n385) );
  XNOR2_X1 U427 ( .A(n679), .B(KEYINPUT83), .ZN(n561) );
  NOR2_X1 U428 ( .A1(n643), .A2(n530), .ZN(n531) );
  XNOR2_X1 U429 ( .A(n406), .B(G146), .ZN(n443) );
  INV_X1 U430 ( .A(G125), .ZN(n406) );
  NOR2_X1 U431 ( .A1(n391), .A2(G953), .ZN(n440) );
  INV_X1 U432 ( .A(G224), .ZN(n391) );
  NAND2_X1 U433 ( .A1(n675), .A2(n674), .ZN(n678) );
  INV_X1 U434 ( .A(KEYINPUT38), .ZN(n361) );
  XNOR2_X1 U435 ( .A(n363), .B(n427), .ZN(n612) );
  XNOR2_X1 U436 ( .A(n431), .B(n426), .ZN(n363) );
  XNOR2_X1 U437 ( .A(n393), .B(n425), .ZN(n426) );
  XNOR2_X1 U438 ( .A(n373), .B(n470), .ZN(n380) );
  XNOR2_X1 U439 ( .A(n412), .B(n407), .ZN(n377) );
  XNOR2_X1 U440 ( .A(n411), .B(n410), .ZN(n412) );
  INV_X1 U441 ( .A(KEYINPUT23), .ZN(n410) );
  XNOR2_X1 U442 ( .A(n443), .B(KEYINPUT10), .ZN(n473) );
  XNOR2_X1 U443 ( .A(G122), .B(KEYINPUT102), .ZN(n388) );
  NOR2_X1 U444 ( .A1(n564), .A2(n563), .ZN(n578) );
  NOR2_X1 U445 ( .A1(n634), .A2(G902), .ZN(n419) );
  XNOR2_X1 U446 ( .A(n542), .B(n433), .ZN(n567) );
  XNOR2_X1 U447 ( .A(n612), .B(KEYINPUT62), .ZN(n613) );
  XNOR2_X1 U448 ( .A(n427), .B(n401), .ZN(n718) );
  XNOR2_X1 U449 ( .A(G107), .B(G104), .ZN(n400) );
  XNOR2_X1 U450 ( .A(n615), .B(KEYINPUT91), .ZN(n721) );
  OR2_X1 U451 ( .A1(n564), .A2(n710), .ZN(n559) );
  BUF_X1 U452 ( .A(n574), .Z(n577) );
  NOR2_X1 U453 ( .A1(n515), .A2(n514), .ZN(n516) );
  OR2_X1 U454 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X1 U455 ( .A(n725), .B(n724), .ZN(n368) );
  AND2_X1 U456 ( .A1(n420), .A2(G217), .ZN(n359) );
  XOR2_X1 U457 ( .A(n534), .B(KEYINPUT45), .Z(n360) );
  XNOR2_X1 U458 ( .A(n591), .B(n361), .ZN(n555) );
  XNOR2_X2 U459 ( .A(n450), .B(n449), .ZN(n591) );
  INV_X1 U460 ( .A(n530), .ZN(n529) );
  XNOR2_X1 U461 ( .A(n358), .B(n362), .ZN(n431) );
  INV_X2 U462 ( .A(KEYINPUT72), .ZN(n383) );
  NOR2_X1 U463 ( .A1(n508), .A2(n709), .ZN(n463) );
  NAND2_X1 U464 ( .A1(n579), .A2(n365), .ZN(n580) );
  NAND2_X1 U465 ( .A1(n533), .A2(n367), .ZN(n535) );
  NAND2_X1 U466 ( .A1(n531), .A2(n532), .ZN(n367) );
  NOR2_X1 U467 ( .A1(n368), .A2(n726), .ZN(G63) );
  NAND2_X1 U468 ( .A1(n369), .A2(n494), .ZN(n495) );
  NAND2_X1 U469 ( .A1(n511), .A2(n369), .ZN(n513) );
  XNOR2_X1 U470 ( .A(n369), .B(n460), .ZN(n508) );
  XNOR2_X2 U471 ( .A(n370), .B(n459), .ZN(n369) );
  NOR2_X2 U472 ( .A1(G902), .A2(n718), .ZN(n403) );
  NOR2_X2 U473 ( .A1(n688), .A2(n687), .ZN(n510) );
  NAND2_X1 U474 ( .A1(n562), .A2(n458), .ZN(n370) );
  NOR2_X2 U475 ( .A1(n591), .A2(n452), .ZN(n372) );
  XNOR2_X1 U476 ( .A(n374), .B(n446), .ZN(n621) );
  XNOR2_X1 U477 ( .A(n374), .B(G101), .ZN(n727) );
  NOR2_X1 U478 ( .A1(n588), .A2(n591), .ZN(n568) );
  NAND2_X1 U479 ( .A1(n567), .A2(n378), .ZN(n588) );
  AND2_X1 U480 ( .A1(n566), .A2(n379), .ZN(n378) );
  XNOR2_X1 U481 ( .A(n387), .B(n386), .ZN(n483) );
  INV_X1 U482 ( .A(n481), .ZN(n386) );
  XNOR2_X2 U483 ( .A(G143), .B(G128), .ZN(n481) );
  XNOR2_X1 U484 ( .A(n482), .B(n388), .ZN(n387) );
  BUF_X1 U485 ( .A(n716), .Z(n723) );
  AND2_X2 U486 ( .A1(n504), .A2(n684), .ZN(n639) );
  BUF_X1 U487 ( .A(n528), .Z(n643) );
  XOR2_X2 U488 ( .A(n403), .B(n402), .Z(n554) );
  NAND2_X1 U489 ( .A1(n503), .A2(n549), .ZN(n687) );
  XNOR2_X2 U490 ( .A(n432), .B(G472), .ZN(n542) );
  XOR2_X1 U491 ( .A(KEYINPUT25), .B(n359), .Z(n392) );
  XOR2_X1 U492 ( .A(n423), .B(n422), .Z(n393) );
  INV_X1 U493 ( .A(KEYINPUT76), .ZN(n430) );
  INV_X1 U494 ( .A(KEYINPUT48), .ZN(n585) );
  XNOR2_X1 U495 ( .A(n466), .B(n465), .ZN(n472) );
  BUF_X1 U496 ( .A(n603), .Z(n669) );
  XNOR2_X1 U497 ( .A(n472), .B(n471), .ZN(n475) );
  NOR2_X1 U498 ( .A1(n574), .A2(n555), .ZN(n546) );
  XNOR2_X1 U499 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n547) );
  XNOR2_X1 U500 ( .A(n718), .B(n717), .ZN(n719) );
  XNOR2_X1 U501 ( .A(n548), .B(n547), .ZN(n751) );
  XNOR2_X1 U502 ( .A(n720), .B(n719), .ZN(n722) );
  XNOR2_X1 U503 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n394) );
  XNOR2_X2 U504 ( .A(n394), .B(n481), .ZN(n438) );
  XNOR2_X1 U505 ( .A(G134), .B(G137), .ZN(n395) );
  XNOR2_X2 U506 ( .A(n438), .B(n395), .ZN(n742) );
  XNOR2_X2 U507 ( .A(n742), .B(G146), .ZN(n427) );
  XOR2_X2 U508 ( .A(G131), .B(G140), .Z(n474) );
  NAND2_X1 U509 ( .A1(G227), .A2(n743), .ZN(n396) );
  XNOR2_X1 U510 ( .A(n474), .B(n396), .ZN(n398) );
  XNOR2_X1 U511 ( .A(n398), .B(n439), .ZN(n399) );
  XNOR2_X1 U512 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U513 ( .A(KEYINPUT71), .B(G469), .ZN(n402) );
  INV_X1 U514 ( .A(KEYINPUT65), .ZN(n404) );
  XNOR2_X1 U515 ( .A(n404), .B(KEYINPUT1), .ZN(n405) );
  XNOR2_X2 U516 ( .A(n554), .B(n405), .ZN(n688) );
  XNOR2_X1 U517 ( .A(KEYINPUT24), .B(KEYINPUT95), .ZN(n407) );
  XOR2_X1 U518 ( .A(KEYINPUT96), .B(G140), .Z(n409) );
  XNOR2_X1 U519 ( .A(n357), .B(G137), .ZN(n408) );
  XNOR2_X1 U520 ( .A(n409), .B(n408), .ZN(n413) );
  NAND2_X1 U521 ( .A1(n743), .A2(G234), .ZN(n415) );
  XNOR2_X1 U522 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n414) );
  XNOR2_X1 U523 ( .A(n415), .B(n414), .ZN(n480) );
  NAND2_X1 U524 ( .A1(n480), .A2(G221), .ZN(n416) );
  XOR2_X1 U525 ( .A(KEYINPUT20), .B(KEYINPUT97), .Z(n418) );
  XNOR2_X1 U526 ( .A(KEYINPUT15), .B(G902), .ZN(n606) );
  NAND2_X1 U527 ( .A1(G234), .A2(n606), .ZN(n417) );
  XNOR2_X1 U528 ( .A(n418), .B(n417), .ZN(n420) );
  XNOR2_X2 U529 ( .A(n419), .B(n392), .ZN(n503) );
  AND2_X1 U530 ( .A1(n420), .A2(G221), .ZN(n421) );
  XNOR2_X1 U531 ( .A(n421), .B(KEYINPUT21), .ZN(n549) );
  XOR2_X1 U532 ( .A(KEYINPUT5), .B(G131), .Z(n423) );
  XOR2_X1 U533 ( .A(KEYINPUT77), .B(n424), .Z(n464) );
  NAND2_X1 U534 ( .A1(n464), .A2(G210), .ZN(n425) );
  INV_X1 U535 ( .A(G902), .ZN(n476) );
  XOR2_X1 U536 ( .A(KEYINPUT6), .B(KEYINPUT104), .Z(n433) );
  NAND2_X1 U537 ( .A1(n510), .A2(n567), .ZN(n435) );
  INV_X1 U538 ( .A(KEYINPUT33), .ZN(n434) );
  XOR2_X1 U539 ( .A(G116), .B(G107), .Z(n479) );
  INV_X1 U540 ( .A(KEYINPUT16), .ZN(n436) );
  XNOR2_X1 U541 ( .A(n479), .B(n436), .ZN(n437) );
  XNOR2_X1 U542 ( .A(n439), .B(n438), .ZN(n445) );
  XNOR2_X1 U543 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n441) );
  XNOR2_X1 U544 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U545 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U546 ( .A(n445), .B(n444), .ZN(n446) );
  INV_X1 U547 ( .A(n606), .ZN(n596) );
  OR2_X2 U548 ( .A1(n621), .A2(n596), .ZN(n450) );
  INV_X1 U549 ( .A(G237), .ZN(n447) );
  NAND2_X1 U550 ( .A1(n476), .A2(n447), .ZN(n451) );
  NAND2_X1 U551 ( .A1(n451), .A2(G210), .ZN(n448) );
  XNOR2_X1 U552 ( .A(n448), .B(KEYINPUT92), .ZN(n449) );
  NAND2_X1 U553 ( .A1(n451), .A2(G214), .ZN(n674) );
  INV_X1 U554 ( .A(n674), .ZN(n452) );
  NOR2_X1 U555 ( .A1(G898), .A2(n743), .ZN(n453) );
  XOR2_X1 U556 ( .A(KEYINPUT93), .B(n453), .Z(n728) );
  NAND2_X1 U557 ( .A1(n728), .A2(G902), .ZN(n454) );
  NAND2_X1 U558 ( .A1(n743), .A2(G952), .ZN(n538) );
  NAND2_X1 U559 ( .A1(n454), .A2(n538), .ZN(n457) );
  NAND2_X1 U560 ( .A1(G237), .A2(G234), .ZN(n456) );
  INV_X1 U561 ( .A(KEYINPUT14), .ZN(n455) );
  XNOR2_X1 U562 ( .A(n456), .B(n455), .ZN(n703) );
  INV_X1 U563 ( .A(n703), .ZN(n540) );
  AND2_X1 U564 ( .A1(n457), .A2(n540), .ZN(n458) );
  INV_X1 U565 ( .A(KEYINPUT0), .ZN(n459) );
  INV_X1 U566 ( .A(KEYINPUT79), .ZN(n461) );
  XNOR2_X1 U567 ( .A(n461), .B(KEYINPUT34), .ZN(n462) );
  XNOR2_X1 U568 ( .A(n463), .B(n462), .ZN(n488) );
  NAND2_X1 U569 ( .A1(n464), .A2(G214), .ZN(n466) );
  XOR2_X1 U570 ( .A(KEYINPUT101), .B(KEYINPUT100), .Z(n465) );
  XOR2_X1 U571 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n468) );
  XNOR2_X1 U572 ( .A(G143), .B(KEYINPUT11), .ZN(n467) );
  XNOR2_X1 U573 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U574 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U575 ( .A(n474), .B(n473), .ZN(n740) );
  XNOR2_X1 U576 ( .A(n475), .B(n740), .ZN(n628) );
  NAND2_X1 U577 ( .A1(n628), .A2(n476), .ZN(n478) );
  XOR2_X1 U578 ( .A(KEYINPUT13), .B(G475), .Z(n477) );
  XNOR2_X1 U579 ( .A(G134), .B(n479), .ZN(n486) );
  NAND2_X1 U580 ( .A1(n480), .A2(G217), .ZN(n484) );
  XNOR2_X1 U581 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n482) );
  XNOR2_X1 U582 ( .A(n484), .B(n483), .ZN(n485) );
  INV_X1 U583 ( .A(n514), .ZN(n493) );
  NAND2_X1 U584 ( .A1(n515), .A2(n493), .ZN(n575) );
  INV_X1 U585 ( .A(n575), .ZN(n487) );
  NAND2_X1 U586 ( .A1(n488), .A2(n487), .ZN(n489) );
  XNOR2_X2 U587 ( .A(n489), .B(KEYINPUT35), .ZN(n528) );
  XNOR2_X1 U588 ( .A(n528), .B(KEYINPUT67), .ZN(n506) );
  NOR2_X1 U589 ( .A1(n688), .A2(n503), .ZN(n490) );
  XNOR2_X1 U590 ( .A(n490), .B(KEYINPUT105), .ZN(n491) );
  NOR2_X1 U591 ( .A1(n567), .A2(n491), .ZN(n492) );
  XNOR2_X1 U592 ( .A(n492), .B(KEYINPUT80), .ZN(n497) );
  OR2_X1 U593 ( .A1(n515), .A2(n493), .ZN(n677) );
  INV_X1 U594 ( .A(n549), .ZN(n683) );
  NOR2_X1 U595 ( .A1(n677), .A2(n683), .ZN(n494) );
  XNOR2_X1 U596 ( .A(n495), .B(KEYINPUT22), .ZN(n520) );
  INV_X1 U597 ( .A(n520), .ZN(n496) );
  XNOR2_X1 U598 ( .A(n498), .B(KEYINPUT32), .ZN(n754) );
  INV_X1 U599 ( .A(n688), .ZN(n499) );
  OR2_X1 U600 ( .A1(n542), .A2(n499), .ZN(n500) );
  OR2_X1 U601 ( .A1(n520), .A2(n500), .ZN(n502) );
  INV_X1 U602 ( .A(KEYINPUT64), .ZN(n501) );
  XNOR2_X1 U603 ( .A(n502), .B(n501), .ZN(n504) );
  INV_X1 U604 ( .A(n503), .ZN(n684) );
  NOR2_X1 U605 ( .A1(n754), .A2(n639), .ZN(n505) );
  NAND2_X1 U606 ( .A1(n505), .A2(n506), .ZN(n524) );
  INV_X1 U607 ( .A(KEYINPUT44), .ZN(n522) );
  OR2_X2 U608 ( .A1(n554), .A2(n687), .ZN(n541) );
  OR2_X1 U609 ( .A1(n542), .A2(n541), .ZN(n507) );
  XNOR2_X2 U610 ( .A(n509), .B(KEYINPUT98), .ZN(n648) );
  NAND2_X1 U611 ( .A1(n542), .A2(n510), .ZN(n695) );
  INV_X1 U612 ( .A(n695), .ZN(n511) );
  INV_X1 U613 ( .A(KEYINPUT31), .ZN(n512) );
  XNOR2_X1 U614 ( .A(n513), .B(n512), .ZN(n662) );
  NAND2_X1 U615 ( .A1(n648), .A2(n662), .ZN(n517) );
  XNOR2_X2 U616 ( .A(KEYINPUT103), .B(n516), .ZN(n663) );
  NAND2_X1 U617 ( .A1(n517), .A2(n561), .ZN(n521) );
  NAND2_X1 U618 ( .A1(n688), .A2(n503), .ZN(n518) );
  OR2_X1 U619 ( .A1(n567), .A2(n518), .ZN(n519) );
  OR2_X1 U620 ( .A1(n520), .A2(n519), .ZN(n645) );
  AND2_X1 U621 ( .A1(n522), .A2(n529), .ZN(n523) );
  NAND2_X1 U622 ( .A1(n524), .A2(n523), .ZN(n533) );
  INV_X1 U623 ( .A(KEYINPUT67), .ZN(n525) );
  NAND2_X1 U624 ( .A1(n525), .A2(KEYINPUT44), .ZN(n526) );
  OR2_X2 U625 ( .A1(n754), .A2(n526), .ZN(n527) );
  NOR2_X2 U626 ( .A1(n527), .A2(n639), .ZN(n532) );
  INV_X1 U627 ( .A(KEYINPUT88), .ZN(n534) );
  XNOR2_X2 U628 ( .A(n535), .B(n360), .ZN(n730) );
  NOR2_X1 U629 ( .A1(G900), .A2(n743), .ZN(n536) );
  NAND2_X1 U630 ( .A1(G902), .A2(n536), .ZN(n537) );
  NAND2_X1 U631 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U632 ( .A1(n540), .A2(n539), .ZN(n550) );
  NAND2_X1 U633 ( .A1(n542), .A2(n674), .ZN(n543) );
  XOR2_X1 U634 ( .A(n543), .B(KEYINPUT30), .Z(n544) );
  NAND2_X1 U635 ( .A1(n545), .A2(n544), .ZN(n574) );
  XNOR2_X1 U636 ( .A(n546), .B(KEYINPUT39), .ZN(n587) );
  NOR2_X1 U637 ( .A1(n587), .A2(n660), .ZN(n548) );
  NAND2_X1 U638 ( .A1(n684), .A2(n549), .ZN(n551) );
  NOR2_X1 U639 ( .A1(n551), .A2(n550), .ZN(n566) );
  NAND2_X1 U640 ( .A1(n542), .A2(n566), .ZN(n552) );
  XNOR2_X1 U641 ( .A(KEYINPUT28), .B(n552), .ZN(n553) );
  OR2_X1 U642 ( .A1(n554), .A2(n553), .ZN(n564) );
  INV_X1 U643 ( .A(n555), .ZN(n675) );
  NOR2_X1 U644 ( .A1(n677), .A2(n678), .ZN(n557) );
  XNOR2_X1 U645 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n556) );
  XOR2_X1 U646 ( .A(n557), .B(n556), .Z(n710) );
  XOR2_X1 U647 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n558) );
  XNOR2_X1 U648 ( .A(n559), .B(n558), .ZN(n753) );
  XNOR2_X1 U649 ( .A(n560), .B(KEYINPUT46), .ZN(n584) );
  INV_X1 U650 ( .A(n356), .ZN(n563) );
  NAND2_X1 U651 ( .A1(n565), .A2(n578), .ZN(n573) );
  XOR2_X1 U652 ( .A(KEYINPUT36), .B(n568), .Z(n569) );
  NOR2_X1 U653 ( .A1(n688), .A2(n569), .ZN(n665) );
  NAND2_X1 U654 ( .A1(KEYINPUT47), .A2(n679), .ZN(n570) );
  XOR2_X1 U655 ( .A(KEYINPUT82), .B(n570), .Z(n571) );
  NOR2_X1 U656 ( .A1(n665), .A2(n571), .ZN(n572) );
  NAND2_X1 U657 ( .A1(n573), .A2(n572), .ZN(n581) );
  OR2_X1 U658 ( .A1(n591), .A2(n575), .ZN(n576) );
  INV_X1 U659 ( .A(n578), .ZN(n657) );
  NAND2_X1 U660 ( .A1(n657), .A2(KEYINPUT47), .ZN(n579) );
  XNOR2_X1 U661 ( .A(n582), .B(KEYINPUT70), .ZN(n583) );
  NAND2_X1 U662 ( .A1(n584), .A2(n583), .ZN(n586) );
  NOR2_X1 U663 ( .A1(n587), .A2(n663), .ZN(n668) );
  INV_X1 U664 ( .A(n588), .ZN(n589) );
  NAND2_X1 U665 ( .A1(n688), .A2(n589), .ZN(n590) );
  XNOR2_X1 U666 ( .A(KEYINPUT43), .B(n590), .ZN(n592) );
  AND2_X1 U667 ( .A1(n591), .A2(n592), .ZN(n641) );
  NOR2_X1 U668 ( .A1(n668), .A2(n641), .ZN(n593) );
  NAND2_X1 U669 ( .A1(n594), .A2(n593), .ZN(n739) );
  NOR2_X1 U670 ( .A1(n730), .A2(n739), .ZN(n603) );
  AND2_X1 U671 ( .A1(n596), .A2(KEYINPUT86), .ZN(n595) );
  NAND2_X1 U672 ( .A1(n603), .A2(n595), .ZN(n601) );
  INV_X1 U673 ( .A(n730), .ZN(n597) );
  NAND2_X1 U674 ( .A1(n597), .A2(n596), .ZN(n599) );
  NOR2_X1 U675 ( .A1(n739), .A2(KEYINPUT86), .ZN(n598) );
  NAND2_X1 U676 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U677 ( .A1(n600), .A2(n601), .ZN(n602) );
  XNOR2_X1 U678 ( .A(n602), .B(KEYINPUT85), .ZN(n605) );
  AND2_X1 U679 ( .A1(n669), .A2(KEYINPUT2), .ZN(n604) );
  OR2_X2 U680 ( .A1(n605), .A2(n604), .ZN(n611) );
  INV_X1 U681 ( .A(n669), .ZN(n609) );
  XNOR2_X1 U682 ( .A(n606), .B(KEYINPUT87), .ZN(n607) );
  AND2_X1 U683 ( .A1(n607), .A2(KEYINPUT2), .ZN(n608) );
  NAND2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X2 U685 ( .A1(n611), .A2(n610), .ZN(n716) );
  NAND2_X1 U686 ( .A1(n716), .A2(G472), .ZN(n614) );
  XNOR2_X1 U687 ( .A(n614), .B(n613), .ZN(n616) );
  NOR2_X1 U688 ( .A1(n743), .A2(G952), .ZN(n615) );
  NAND2_X1 U689 ( .A1(n616), .A2(n721), .ZN(n618) );
  XOR2_X1 U690 ( .A(KEYINPUT63), .B(KEYINPUT89), .Z(n617) );
  XNOR2_X1 U691 ( .A(n618), .B(n617), .ZN(G57) );
  NAND2_X1 U692 ( .A1(n716), .A2(G210), .ZN(n623) );
  XNOR2_X1 U693 ( .A(KEYINPUT90), .B(KEYINPUT54), .ZN(n619) );
  XNOR2_X1 U694 ( .A(n619), .B(KEYINPUT55), .ZN(n620) );
  XNOR2_X1 U695 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U696 ( .A(n623), .B(n622), .ZN(n624) );
  NAND2_X1 U697 ( .A1(n624), .A2(n721), .ZN(n626) );
  INV_X1 U698 ( .A(KEYINPUT56), .ZN(n625) );
  XNOR2_X1 U699 ( .A(n626), .B(n625), .ZN(G51) );
  NAND2_X1 U700 ( .A1(n716), .A2(G475), .ZN(n630) );
  XNOR2_X1 U701 ( .A(KEYINPUT121), .B(KEYINPUT59), .ZN(n627) );
  XNOR2_X1 U702 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U703 ( .A(n630), .B(n629), .ZN(n631) );
  NAND2_X1 U704 ( .A1(n631), .A2(n721), .ZN(n633) );
  INV_X1 U705 ( .A(KEYINPUT60), .ZN(n632) );
  XNOR2_X1 U706 ( .A(n633), .B(n632), .ZN(G60) );
  NAND2_X1 U707 ( .A1(n716), .A2(G217), .ZN(n636) );
  XNOR2_X1 U708 ( .A(n636), .B(n635), .ZN(n637) );
  NAND2_X1 U709 ( .A1(n637), .A2(n721), .ZN(n638) );
  XNOR2_X1 U710 ( .A(n638), .B(KEYINPUT123), .ZN(G66) );
  XOR2_X1 U711 ( .A(G110), .B(n639), .Z(G12) );
  XNOR2_X1 U712 ( .A(G140), .B(KEYINPUT116), .ZN(n640) );
  XOR2_X1 U713 ( .A(n641), .B(n640), .Z(G42) );
  XOR2_X1 U714 ( .A(G143), .B(n642), .Z(G45) );
  XOR2_X1 U715 ( .A(n643), .B(G122), .Z(G24) );
  XOR2_X1 U716 ( .A(G101), .B(KEYINPUT109), .Z(n644) );
  XNOR2_X1 U717 ( .A(n645), .B(n644), .ZN(G3) );
  NOR2_X1 U718 ( .A1(n648), .A2(n660), .ZN(n646) );
  XOR2_X1 U719 ( .A(KEYINPUT110), .B(n646), .Z(n647) );
  XNOR2_X1 U720 ( .A(G104), .B(n647), .ZN(G6) );
  NOR2_X1 U721 ( .A1(n648), .A2(n663), .ZN(n653) );
  XOR2_X1 U722 ( .A(KEYINPUT27), .B(KEYINPUT112), .Z(n650) );
  XNOR2_X1 U723 ( .A(G107), .B(KEYINPUT111), .ZN(n649) );
  XNOR2_X1 U724 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U725 ( .A(KEYINPUT26), .B(n651), .ZN(n652) );
  XNOR2_X1 U726 ( .A(n653), .B(n652), .ZN(G9) );
  NOR2_X1 U727 ( .A1(n657), .A2(n663), .ZN(n655) );
  XNOR2_X1 U728 ( .A(KEYINPUT113), .B(KEYINPUT29), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n655), .B(n654), .ZN(n656) );
  XOR2_X1 U730 ( .A(n357), .B(n656), .Z(G30) );
  NOR2_X1 U731 ( .A1(n657), .A2(n660), .ZN(n658) );
  XOR2_X1 U732 ( .A(KEYINPUT114), .B(n658), .Z(n659) );
  XNOR2_X1 U733 ( .A(G146), .B(n659), .ZN(G48) );
  NOR2_X1 U734 ( .A1(n660), .A2(n662), .ZN(n661) );
  XOR2_X1 U735 ( .A(G113), .B(n661), .Z(G15) );
  NOR2_X1 U736 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U737 ( .A(G116), .B(n664), .Z(G18) );
  XOR2_X1 U738 ( .A(KEYINPUT37), .B(KEYINPUT115), .Z(n667) );
  XNOR2_X1 U739 ( .A(G125), .B(n665), .ZN(n666) );
  XNOR2_X1 U740 ( .A(n667), .B(n666), .ZN(G27) );
  XOR2_X1 U741 ( .A(G134), .B(n668), .Z(G36) );
  XOR2_X1 U742 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n715) );
  NOR2_X1 U743 ( .A1(n669), .A2(KEYINPUT81), .ZN(n673) );
  INV_X1 U744 ( .A(n673), .ZN(n671) );
  NAND2_X1 U745 ( .A1(n669), .A2(KEYINPUT81), .ZN(n670) );
  NAND2_X1 U746 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U747 ( .A1(KEYINPUT2), .A2(n672), .ZN(n708) );
  NAND2_X1 U748 ( .A1(n673), .A2(KEYINPUT2), .ZN(n706) );
  NOR2_X1 U749 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U750 ( .A1(n677), .A2(n676), .ZN(n681) );
  NOR2_X1 U751 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U752 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U753 ( .A1(n682), .A2(n709), .ZN(n699) );
  NAND2_X1 U754 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U755 ( .A(n685), .B(KEYINPUT117), .ZN(n686) );
  XNOR2_X1 U756 ( .A(KEYINPUT49), .B(n686), .ZN(n693) );
  XOR2_X1 U757 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n690) );
  NAND2_X1 U758 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U759 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X1 U760 ( .A1(n691), .A2(n542), .ZN(n692) );
  NAND2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U762 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U763 ( .A(KEYINPUT51), .B(n696), .ZN(n697) );
  NOR2_X1 U764 ( .A1(n710), .A2(n697), .ZN(n698) );
  NOR2_X1 U765 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U766 ( .A(n700), .B(KEYINPUT119), .Z(n701) );
  XNOR2_X1 U767 ( .A(KEYINPUT52), .B(n701), .ZN(n702) );
  NOR2_X1 U768 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U769 ( .A1(n704), .A2(G952), .ZN(n705) );
  NAND2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U771 ( .A1(n708), .A2(n707), .ZN(n713) );
  NOR2_X1 U772 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U773 ( .A1(G953), .A2(n711), .ZN(n712) );
  NAND2_X1 U774 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U775 ( .A(n715), .B(n714), .ZN(G75) );
  NAND2_X1 U776 ( .A1(n723), .A2(G469), .ZN(n720) );
  XOR2_X1 U777 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n717) );
  INV_X1 U778 ( .A(n721), .ZN(n726) );
  NOR2_X1 U779 ( .A1(n722), .A2(n726), .ZN(G54) );
  NAND2_X1 U780 ( .A1(n723), .A2(G478), .ZN(n725) );
  XNOR2_X1 U781 ( .A(n727), .B(G110), .ZN(n729) );
  NOR2_X1 U782 ( .A1(n729), .A2(n728), .ZN(n738) );
  NOR2_X1 U783 ( .A1(n730), .A2(G953), .ZN(n731) );
  XNOR2_X1 U784 ( .A(n731), .B(KEYINPUT125), .ZN(n736) );
  NAND2_X1 U785 ( .A1(G953), .A2(G224), .ZN(n732) );
  XNOR2_X1 U786 ( .A(KEYINPUT61), .B(n732), .ZN(n733) );
  NAND2_X1 U787 ( .A1(n733), .A2(G898), .ZN(n734) );
  XNOR2_X1 U788 ( .A(KEYINPUT124), .B(n734), .ZN(n735) );
  NAND2_X1 U789 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U790 ( .A(n738), .B(n737), .ZN(G69) );
  XOR2_X1 U791 ( .A(n740), .B(KEYINPUT126), .Z(n741) );
  XNOR2_X1 U792 ( .A(n742), .B(n741), .ZN(n745) );
  XNOR2_X1 U793 ( .A(n355), .B(n745), .ZN(n744) );
  NAND2_X1 U794 ( .A1(n744), .A2(n743), .ZN(n750) );
  XNOR2_X1 U795 ( .A(G227), .B(n745), .ZN(n746) );
  NAND2_X1 U796 ( .A1(n746), .A2(G900), .ZN(n747) );
  XOR2_X1 U797 ( .A(KEYINPUT127), .B(n747), .Z(n748) );
  NAND2_X1 U798 ( .A1(G953), .A2(n748), .ZN(n749) );
  NAND2_X1 U799 ( .A1(n750), .A2(n749), .ZN(G72) );
  BUF_X1 U800 ( .A(n751), .Z(n752) );
  XOR2_X1 U801 ( .A(G131), .B(n752), .Z(G33) );
  XOR2_X1 U802 ( .A(G137), .B(n753), .Z(G39) );
  XOR2_X1 U803 ( .A(G119), .B(n754), .Z(G21) );
endmodule

