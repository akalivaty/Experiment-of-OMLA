//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G211gat), .B(G218gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT69), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT69), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G218gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT22), .B1(new_n212), .B2(G211gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(G197gat), .B(G204gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n207), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G211gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n217), .B1(new_n209), .B2(new_n211), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n214), .B(new_n206), .C1(new_n218), .C2(KEYINPUT22), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n222));
  INV_X1    g021(.A(G183gat), .ZN(new_n223));
  INV_X1    g022(.A(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G169gat), .ZN(new_n230));
  INV_X1    g029(.A(G176gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT23), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT23), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(G169gat), .B2(G176gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n222), .B1(new_n229), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n238));
  NOR3_X1   g037(.A1(new_n233), .A2(G169gat), .A3(G176gat), .ZN(new_n239));
  INV_X1    g038(.A(new_n235), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n232), .A2(KEYINPUT65), .A3(new_n235), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n234), .A2(KEYINPUT25), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n247));
  NOR3_X1   g046(.A1(new_n246), .A2(new_n247), .A3(new_n227), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n237), .B1(new_n244), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(G226gat), .A2(G233gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n230), .A2(new_n231), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n251), .A2(KEYINPUT26), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n251), .B1(new_n240), .B2(KEYINPUT26), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n252), .A2(new_n253), .B1(G183gat), .B2(G190gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT28), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT27), .B(G183gat), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n255), .B1(new_n256), .B2(new_n224), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n256), .A2(new_n255), .A3(new_n224), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n254), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n249), .A2(new_n250), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n262), .B1(new_n249), .B2(new_n260), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n221), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n249), .A2(new_n250), .A3(new_n260), .ZN(new_n265));
  OR2_X1    g064(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n266), .A2(new_n245), .A3(new_n225), .A4(new_n226), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n267), .A2(new_n242), .A3(new_n241), .A4(new_n243), .ZN(new_n268));
  INV_X1    g067(.A(new_n259), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n269), .A2(new_n257), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n268), .A2(new_n237), .B1(new_n270), .B2(new_n254), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n265), .B(new_n220), .C1(new_n271), .C2(new_n262), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n264), .A2(KEYINPUT70), .A3(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n274), .B(new_n221), .C1(new_n261), .C2(new_n263), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n205), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G113gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n278), .A2(KEYINPUT67), .A3(G120gat), .ZN(new_n279));
  INV_X1    g078(.A(G134gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(G127gat), .ZN(new_n281));
  INV_X1    g080(.A(G127gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G134gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n279), .A2(new_n281), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G120gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G113gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n278), .A2(G120gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT67), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n288), .A2(new_n289), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(new_n284), .ZN(new_n293));
  XNOR2_X1  g092(.A(G127gat), .B(G134gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n286), .A2(new_n291), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G141gat), .B(G148gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G155gat), .ZN(new_n302));
  INV_X1    g101(.A(G162gat), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT2), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OR2_X1    g103(.A1(KEYINPUT72), .A2(KEYINPUT2), .ZN(new_n305));
  OR2_X1    g104(.A1(G141gat), .A2(G148gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(KEYINPUT72), .A2(KEYINPUT2), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n305), .A2(new_n306), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n301), .A2(new_n304), .B1(new_n299), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT73), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n296), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n309), .A2(new_n299), .ZN(new_n313));
  XNOR2_X1  g112(.A(G155gat), .B(G162gat), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n314), .A2(new_n306), .A3(new_n304), .A4(new_n307), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT1), .B1(new_n288), .B2(new_n289), .ZN(new_n318));
  OAI22_X1  g117(.A1(new_n317), .A2(new_n285), .B1(new_n318), .B2(new_n294), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT73), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT4), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n312), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G225gat), .A2(G233gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n316), .A2(new_n319), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT4), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n316), .A2(KEYINPUT3), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(new_n319), .A3(new_n328), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n322), .A2(new_n323), .A3(new_n325), .A4(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT5), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n319), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n312), .A2(new_n320), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n323), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n331), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n330), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI211_X1 g136(.A(KEYINPUT74), .B(new_n331), .C1(new_n333), .C2(new_n334), .ZN(new_n338));
  OR2_X1    g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n311), .B1(new_n296), .B2(new_n310), .ZN(new_n340));
  NOR3_X1   g139(.A1(new_n316), .A2(new_n319), .A3(KEYINPUT73), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT4), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT75), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n324), .A2(KEYINPUT4), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n321), .B1(new_n312), .B2(new_n320), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT75), .B1(new_n347), .B2(new_n344), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n329), .A2(new_n331), .A3(new_n323), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT76), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n353));
  AOI211_X1 g152(.A(new_n353), .B(new_n350), .C1(new_n346), .C2(new_n348), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n339), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G1gat), .B(G29gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(KEYINPUT0), .ZN(new_n357));
  XNOR2_X1  g156(.A(G57gat), .B(G85gat), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n357), .B(new_n358), .Z(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n355), .A2(KEYINPUT6), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n273), .A2(new_n275), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT37), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n205), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n363), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT84), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT84), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n362), .A2(new_n367), .A3(new_n363), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n364), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT38), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n277), .B(new_n361), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT82), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT6), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n337), .A2(new_n338), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n343), .B1(new_n342), .B2(new_n345), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n347), .A2(KEYINPUT75), .A3(new_n344), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n351), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(new_n353), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n349), .A2(KEYINPUT76), .A3(new_n351), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n375), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n374), .B1(new_n381), .B2(new_n359), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n339), .B(new_n359), .C1(new_n352), .C2(new_n354), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n373), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n355), .A2(new_n360), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n386), .A2(KEYINPUT82), .A3(new_n374), .A4(new_n383), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n205), .A2(new_n370), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n264), .A2(KEYINPUT83), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT83), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n390), .B(new_n221), .C1(new_n261), .C2(new_n263), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n272), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n388), .B1(new_n392), .B2(KEYINPUT37), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n367), .B1(new_n362), .B2(new_n363), .ZN(new_n394));
  AOI211_X1 g193(.A(KEYINPUT84), .B(KEYINPUT37), .C1(new_n273), .C2(new_n275), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT85), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT85), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n398), .B(new_n393), .C1(new_n394), .C2(new_n395), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n372), .A2(new_n385), .A3(new_n387), .A4(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n329), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n402), .B1(new_n346), .B2(new_n348), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT39), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n405), .A3(new_n334), .ZN(new_n406));
  OR2_X1    g205(.A1(new_n333), .A2(new_n334), .ZN(new_n407));
  OAI211_X1 g206(.A(KEYINPUT39), .B(new_n407), .C1(new_n403), .C2(new_n323), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n359), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT40), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n406), .A2(new_n408), .A3(KEYINPUT40), .A4(new_n359), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AND2_X1   g212(.A1(KEYINPUT71), .A2(KEYINPUT30), .ZN(new_n414));
  NOR2_X1   g213(.A1(KEYINPUT71), .A2(KEYINPUT30), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n276), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n273), .A2(new_n275), .A3(new_n205), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n414), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n417), .B1(new_n419), .B2(new_n276), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n386), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT81), .B1(new_n413), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n420), .B1(new_n360), .B2(new_n355), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT81), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n424), .A2(new_n425), .A3(new_n412), .A4(new_n411), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  XOR2_X1   g226(.A(G78gat), .B(G106gat), .Z(new_n428));
  XNOR2_X1  g227(.A(KEYINPUT31), .B(G50gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT80), .ZN(new_n431));
  INV_X1    g230(.A(G228gat), .ZN(new_n432));
  INV_X1    g231(.A(G233gat), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT29), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n327), .A2(new_n435), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n436), .A2(new_n221), .B1(KEYINPUT3), .B2(new_n316), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT29), .B1(new_n216), .B2(new_n219), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n316), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n434), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n219), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT22), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT69), .B(G218gat), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n442), .B1(new_n443), .B2(new_n217), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n206), .B1(new_n444), .B2(new_n214), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n435), .B1(new_n441), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT3), .B1(new_n446), .B2(KEYINPUT77), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT77), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n220), .A2(new_n448), .A3(new_n435), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n310), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT29), .B1(new_n310), .B2(new_n326), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n434), .B1(new_n451), .B2(new_n220), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT78), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n326), .B1(new_n438), .B2(new_n448), .ZN(new_n454));
  AOI211_X1 g253(.A(KEYINPUT77), .B(KEYINPUT29), .C1(new_n216), .C2(new_n219), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n316), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n452), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT78), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n440), .B1(new_n453), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(G22gat), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n431), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n440), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n446), .A2(KEYINPUT77), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n464), .A2(new_n326), .A3(new_n449), .ZN(new_n465));
  AOI211_X1 g264(.A(KEYINPUT78), .B(new_n452), .C1(new_n465), .C2(new_n316), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n458), .B1(new_n456), .B2(new_n457), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n468), .A2(KEYINPUT80), .A3(G22gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n462), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n461), .B(new_n463), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT79), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n453), .A2(new_n459), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n474), .A2(KEYINPUT79), .A3(new_n461), .A4(new_n463), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n430), .B1(new_n470), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n430), .B1(new_n468), .B2(G22gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n471), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n401), .A2(new_n427), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT36), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n249), .A2(new_n260), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n296), .ZN(new_n484));
  NAND2_X1  g283(.A1(G227gat), .A2(G233gat), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n249), .A2(new_n319), .A3(new_n260), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT33), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XOR2_X1   g289(.A(G15gat), .B(G43gat), .Z(new_n491));
  XNOR2_X1  g290(.A(G71gat), .B(G99gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n484), .A2(new_n487), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n485), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT34), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT34), .ZN(new_n498));
  INV_X1    g297(.A(new_n487), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n319), .B1(new_n249), .B2(new_n260), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n498), .B(new_n485), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n494), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n501), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n498), .B1(new_n495), .B2(new_n485), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n490), .B(new_n493), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n488), .A2(KEYINPUT32), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n502), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n507), .B1(new_n502), .B2(new_n505), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n482), .B1(new_n510), .B2(KEYINPUT68), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT68), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n512), .B(KEYINPUT36), .C1(new_n508), .C2(new_n509), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n477), .A2(new_n479), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n386), .A2(new_n374), .A3(new_n383), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n421), .B1(new_n516), .B2(new_n361), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n514), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n481), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n480), .A2(new_n517), .A3(new_n510), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT35), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n385), .A2(new_n387), .A3(new_n361), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n502), .A2(new_n505), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n506), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n502), .A2(new_n505), .A3(new_n507), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n527), .A2(new_n421), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT35), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n523), .A2(new_n528), .A3(new_n480), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n522), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n520), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(G43gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(G50gat), .ZN(new_n534));
  INV_X1    g333(.A(G50gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(G43gat), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n534), .A2(new_n536), .A3(KEYINPUT15), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(KEYINPUT86), .B(KEYINPUT15), .Z(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT87), .B(G50gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n533), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n541), .A2(KEYINPUT88), .B1(G43gat), .B2(new_n535), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT88), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n540), .A2(new_n543), .A3(new_n533), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n539), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(KEYINPUT14), .B(G29gat), .Z(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(G36gat), .ZN(new_n547));
  INV_X1    g346(.A(G29gat), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n548), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n538), .B1(new_n545), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT17), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n537), .B1(new_n547), .B2(new_n549), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT89), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n551), .A2(KEYINPUT89), .A3(new_n552), .A4(new_n553), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G15gat), .B(G22gat), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n559), .A2(G1gat), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT16), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n559), .B1(new_n561), .B2(G1gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(G8gat), .ZN(new_n564));
  INV_X1    g363(.A(G8gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n560), .A2(new_n565), .A3(new_n562), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT90), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n564), .A2(KEYINPUT90), .A3(new_n566), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n551), .A2(new_n553), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n571), .B1(KEYINPUT17), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G229gat), .A2(G233gat), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n551), .A2(new_n553), .A3(new_n567), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT18), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n574), .A2(KEYINPUT18), .A3(new_n575), .A4(new_n576), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n575), .B(KEYINPUT13), .Z(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n567), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n572), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n582), .B1(new_n584), .B2(new_n576), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT91), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n579), .A2(new_n580), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G113gat), .B(G141gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(G197gat), .ZN(new_n589));
  XOR2_X1   g388(.A(KEYINPUT11), .B(G169gat), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n591), .B(KEYINPUT12), .Z(new_n592));
  NAND2_X1  g391(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n592), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n579), .A2(new_n594), .A3(new_n580), .A4(new_n586), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G232gat), .A2(G233gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n597), .B(KEYINPUT94), .Z(new_n598));
  INV_X1    g397(.A(KEYINPUT41), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G134gat), .B(G162gat), .Z(new_n601));
  XOR2_X1   g400(.A(new_n600), .B(new_n601), .Z(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G85gat), .A2(G92gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT7), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  INV_X1    g405(.A(G85gat), .ZN(new_n607));
  INV_X1    g406(.A(G92gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G99gat), .B(G106gat), .Z(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n611), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n613), .A2(new_n605), .A3(new_n609), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  OAI22_X1  g414(.A1(new_n572), .A2(new_n615), .B1(new_n599), .B2(new_n598), .ZN(new_n616));
  INV_X1    g415(.A(new_n615), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n617), .B1(new_n572), .B2(KEYINPUT17), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n616), .B1(new_n558), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G190gat), .B(G218gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT95), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n619), .A2(new_n620), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n603), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AND2_X1   g424(.A1(G71gat), .A2(G78gat), .ZN(new_n626));
  NOR2_X1   g425(.A1(G71gat), .A2(G78gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(G57gat), .B(G64gat), .Z(new_n629));
  INV_X1    g428(.A(KEYINPUT92), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n629), .B1(KEYINPUT9), .B2(new_n626), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI221_X1 g432(.A(new_n629), .B1(KEYINPUT9), .B2(new_n626), .C1(new_n628), .C2(new_n630), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT93), .B(KEYINPUT21), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(G231gat), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n433), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n635), .B(new_n636), .C1(new_n638), .C2(new_n433), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(G127gat), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n640), .A2(new_n282), .A3(new_n641), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n633), .A2(new_n634), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n567), .B1(KEYINPUT21), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n647), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n643), .A2(new_n649), .A3(new_n644), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(new_n302), .ZN(new_n653));
  XNOR2_X1  g452(.A(G183gat), .B(G211gat), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n653), .B(new_n654), .Z(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n648), .A2(new_n650), .A3(new_n655), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(KEYINPUT95), .B1(new_n619), .B2(new_n620), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n660), .B(new_n602), .C1(new_n619), .C2(new_n620), .ZN(new_n661));
  NAND2_X1  g460(.A1(G230gat), .A2(G233gat), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT96), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n614), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n646), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n617), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n646), .A2(new_n615), .A3(new_n664), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT10), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n617), .A2(KEYINPUT10), .A3(new_n646), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n662), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n666), .A2(new_n667), .ZN(new_n672));
  INV_X1    g471(.A(new_n662), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(G120gat), .B(G148gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(G176gat), .B(G204gat), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n675), .B(new_n676), .Z(new_n677));
  NAND3_X1  g476(.A1(new_n671), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n677), .B1(new_n671), .B2(new_n674), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n625), .A2(new_n659), .A3(new_n661), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT97), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n532), .A2(new_n596), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n516), .A2(new_n361), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT98), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g488(.A1(new_n684), .A2(new_n420), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT16), .B(G8gat), .Z(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(new_n565), .B2(new_n690), .ZN(new_n693));
  MUX2_X1   g492(.A(new_n692), .B(new_n693), .S(KEYINPUT42), .Z(G1325gat));
  AOI21_X1  g493(.A(KEYINPUT36), .B1(new_n527), .B2(new_n512), .ZN(new_n695));
  INV_X1    g494(.A(new_n513), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G15gat), .B1(new_n684), .B2(new_n697), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n527), .A2(G15gat), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n698), .B1(new_n684), .B2(new_n699), .ZN(G1326gat));
  NOR2_X1   g499(.A1(new_n684), .A2(new_n480), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT43), .B(G22gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1327gat));
  NAND2_X1  g502(.A1(new_n625), .A2(new_n661), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n532), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n596), .ZN(new_n707));
  INV_X1    g506(.A(new_n681), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n707), .A2(new_n659), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n711), .A2(new_n548), .A3(new_n686), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT45), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714));
  AOI22_X1  g513(.A1(new_n481), .A2(new_n519), .B1(new_n522), .B2(new_n530), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n625), .A2(new_n661), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n697), .B1(new_n480), .B2(new_n517), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n397), .A2(new_n399), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(new_n371), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n385), .A2(new_n387), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n515), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n718), .B1(new_n722), .B2(new_n427), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n523), .A2(new_n529), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n480), .A2(new_n528), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n724), .A2(new_n725), .B1(KEYINPUT35), .B2(new_n521), .ZN(new_n726));
  OAI211_X1 g525(.A(KEYINPUT44), .B(new_n704), .C1(new_n723), .C2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n717), .A2(new_n709), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT99), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n717), .A2(new_n727), .A3(KEYINPUT99), .A4(new_n709), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n730), .A2(new_n686), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n713), .B1(new_n548), .B2(new_n732), .ZN(G1328gat));
  NOR3_X1   g532(.A1(new_n710), .A2(G36gat), .A3(new_n420), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT46), .ZN(new_n735));
  INV_X1    g534(.A(G36gat), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n730), .A2(new_n421), .A3(new_n731), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(G1329gat));
  NOR3_X1   g537(.A1(new_n710), .A2(G43gat), .A3(new_n527), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(G43gat), .B1(new_n728), .B2(new_n697), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n740), .A2(KEYINPUT47), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n730), .A2(new_n514), .A3(new_n731), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT100), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n743), .A2(new_n744), .A3(G43gat), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n744), .B1(new_n743), .B2(G43gat), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n745), .A2(new_n746), .A3(new_n739), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n742), .B1(new_n747), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g547(.A1(new_n710), .A2(new_n480), .A3(new_n540), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n540), .B1(new_n728), .B2(new_n480), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n750), .A2(KEYINPUT48), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n730), .A2(new_n515), .A3(new_n731), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n540), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n750), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT48), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT101), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n749), .B1(new_n753), .B2(new_n540), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT101), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n758), .A2(new_n759), .A3(KEYINPUT48), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n752), .B1(new_n757), .B2(new_n760), .ZN(G1331gat));
  NAND4_X1  g560(.A1(new_n707), .A2(new_n659), .A3(new_n716), .A4(new_n708), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n715), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n686), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n763), .A2(new_n421), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1333gat));
  INV_X1    g570(.A(G71gat), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n763), .A2(new_n772), .A3(new_n510), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n715), .A2(new_n697), .A3(new_n762), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(new_n772), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n775), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g575(.A1(new_n763), .A2(new_n515), .ZN(new_n777));
  XNOR2_X1  g576(.A(KEYINPUT104), .B(G78gat), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n777), .B(new_n778), .ZN(G1335gat));
  NOR2_X1   g578(.A1(new_n596), .A2(new_n659), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n705), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n782), .B1(KEYINPUT107), .B2(KEYINPUT51), .ZN(new_n783));
  OR2_X1    g582(.A1(KEYINPUT107), .A2(KEYINPUT51), .ZN(new_n784));
  XOR2_X1   g583(.A(new_n783), .B(new_n784), .Z(new_n785));
  NAND4_X1  g584(.A1(new_n785), .A2(new_n607), .A3(new_n708), .A4(new_n686), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n780), .A2(new_n708), .ZN(new_n787));
  XOR2_X1   g586(.A(new_n787), .B(KEYINPUT105), .Z(new_n788));
  NAND3_X1  g587(.A1(new_n717), .A2(new_n727), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT106), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n717), .A2(new_n727), .A3(new_n788), .A4(KEYINPUT106), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(new_n686), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G85gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n786), .A2(new_n794), .ZN(G1336gat));
  OR2_X1    g594(.A1(new_n783), .A2(new_n784), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n783), .A2(new_n784), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n421), .A2(new_n608), .A3(new_n708), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT108), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n796), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801));
  OAI21_X1  g600(.A(G92gat), .B1(new_n789), .B2(new_n420), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT51), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT109), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n782), .B2(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(KEYINPUT109), .B(KEYINPUT51), .C1(new_n705), .C2(new_n781), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n791), .A2(new_n421), .A3(new_n792), .ZN(new_n809));
  AOI22_X1  g608(.A1(new_n808), .A2(new_n799), .B1(new_n809), .B2(G92gat), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n803), .B1(new_n801), .B2(new_n810), .ZN(G1337gat));
  NOR3_X1   g610(.A1(new_n527), .A2(G99gat), .A3(new_n681), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n785), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n791), .A2(new_n514), .A3(new_n792), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G99gat), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(G1338gat));
  NOR3_X1   g615(.A1(new_n480), .A2(G106gat), .A3(new_n681), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n806), .A2(new_n807), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT111), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n806), .A2(new_n807), .A3(new_n820), .A4(new_n817), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n791), .A2(new_n515), .A3(new_n792), .ZN(new_n823));
  XNOR2_X1  g622(.A(KEYINPUT110), .B(G106gat), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT53), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n796), .A2(new_n797), .A3(new_n817), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n824), .B1(new_n789), .B2(new_n480), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n826), .A2(new_n830), .ZN(G1339gat));
  INV_X1    g630(.A(KEYINPUT114), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n671), .A2(KEYINPUT54), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT112), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n669), .B1(new_n672), .B2(KEYINPUT10), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(new_n662), .ZN(new_n837));
  NOR4_X1   g636(.A1(new_n668), .A2(new_n670), .A3(new_n835), .A4(new_n662), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n834), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n677), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n841), .B1(new_n671), .B2(KEYINPUT54), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n833), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n842), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n668), .A2(new_n670), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT112), .B1(new_n845), .B2(new_n673), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n838), .ZN(new_n847));
  OAI211_X1 g646(.A(KEYINPUT55), .B(new_n844), .C1(new_n847), .C2(new_n834), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n843), .A2(new_n678), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n849), .B1(new_n593), .B2(new_n595), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n584), .A2(new_n576), .A3(new_n582), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT113), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n575), .B1(new_n574), .B2(new_n576), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n591), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n595), .A2(new_n708), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n832), .B1(new_n850), .B2(new_n855), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n843), .A2(new_n678), .A3(new_n848), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n596), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n855), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n858), .A2(new_n859), .A3(KEYINPUT114), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n856), .A2(new_n716), .A3(new_n860), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n595), .A2(new_n854), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n857), .A2(new_n862), .A3(new_n704), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n659), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n596), .A2(new_n682), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n687), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n725), .ZN(new_n868));
  OAI21_X1  g667(.A(G113gat), .B1(new_n868), .B2(new_n707), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n596), .A2(new_n278), .ZN(new_n870));
  XOR2_X1   g669(.A(new_n870), .B(KEYINPUT115), .Z(new_n871));
  OAI21_X1  g670(.A(new_n869), .B1(new_n868), .B2(new_n871), .ZN(G1340gat));
  NOR2_X1   g671(.A1(new_n868), .A2(new_n681), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(new_n287), .ZN(G1341gat));
  INV_X1    g673(.A(new_n659), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(new_n282), .ZN(G1342gat));
  NAND2_X1  g676(.A1(new_n480), .A2(new_n510), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n704), .A2(new_n420), .ZN(new_n880));
  XOR2_X1   g679(.A(new_n880), .B(KEYINPUT116), .Z(new_n881));
  NAND4_X1  g680(.A1(new_n867), .A2(new_n280), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n882), .B(KEYINPUT56), .Z(new_n883));
  OAI21_X1  g682(.A(G134gat), .B1(new_n868), .B2(new_n716), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(G1343gat));
  NOR2_X1   g684(.A1(new_n866), .A2(new_n480), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n686), .A2(new_n697), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n887), .A2(new_n421), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(G141gat), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n596), .A2(new_n891), .ZN(new_n892));
  XOR2_X1   g691(.A(new_n892), .B(KEYINPUT119), .Z(new_n893));
  AOI21_X1  g692(.A(KEYINPUT120), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n888), .ZN(new_n895));
  XNOR2_X1  g694(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n896), .B1(new_n866), .B2(new_n480), .ZN(new_n897));
  INV_X1    g696(.A(new_n865), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n704), .B1(new_n858), .B2(new_n859), .ZN(new_n899));
  INV_X1    g698(.A(new_n863), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n875), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n898), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n855), .B1(new_n596), .B2(new_n857), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n863), .B1(new_n904), .B2(new_n704), .ZN(new_n905));
  AOI21_X1  g704(.A(KEYINPUT118), .B1(new_n905), .B2(new_n875), .ZN(new_n906));
  OAI211_X1 g705(.A(KEYINPUT57), .B(new_n515), .C1(new_n903), .C2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n895), .B1(new_n897), .B2(new_n907), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n908), .A2(new_n596), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n894), .B1(new_n909), .B2(new_n891), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT58), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT58), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n912), .B(new_n894), .C1(new_n909), .C2(new_n891), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1344gat));
  INV_X1    g713(.A(KEYINPUT59), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n908), .A2(new_n915), .A3(new_n708), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT57), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n716), .A2(KEYINPUT97), .A3(new_n659), .A4(new_n681), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT97), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n682), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n918), .A2(new_n707), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT121), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n918), .A2(new_n923), .A3(new_n707), .A4(new_n920), .ZN(new_n924));
  AOI22_X1  g723(.A1(new_n922), .A2(new_n924), .B1(new_n905), .B2(new_n875), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n515), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n923), .B1(new_n683), .B2(new_n707), .ZN(new_n928));
  INV_X1    g727(.A(new_n924), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n901), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n930), .A2(KEYINPUT122), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n917), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n896), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n515), .B(new_n933), .C1(new_n864), .C2(new_n865), .ZN(new_n934));
  AOI211_X1 g733(.A(new_n681), .B(new_n895), .C1(new_n932), .C2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n915), .B1(new_n890), .B2(new_n708), .ZN(new_n937));
  OAI221_X1 g736(.A(new_n916), .B1(new_n935), .B2(new_n936), .C1(new_n937), .C2(G148gat), .ZN(G1345gat));
  NAND3_X1  g737(.A1(new_n890), .A2(new_n302), .A3(new_n659), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n908), .A2(new_n659), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(new_n302), .ZN(G1346gat));
  INV_X1    g740(.A(new_n887), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n886), .A2(new_n303), .A3(new_n881), .A4(new_n942), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n908), .A2(new_n704), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n944), .B2(new_n303), .ZN(G1347gat));
  AOI21_X1  g744(.A(new_n704), .B1(new_n904), .B2(KEYINPUT114), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n900), .B1(new_n946), .B2(new_n856), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n898), .B1(new_n947), .B2(new_n659), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n686), .A2(new_n420), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n879), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n951), .A2(new_n707), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(new_n230), .ZN(G1348gat));
  NOR2_X1   g752(.A1(new_n951), .A2(new_n681), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(new_n231), .ZN(G1349gat));
  OR3_X1    g754(.A1(new_n951), .A2(new_n256), .A3(new_n875), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n223), .B1(new_n951), .B2(new_n875), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT60), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n958), .B(new_n959), .ZN(G1350gat));
  OAI22_X1  g759(.A1(new_n951), .A2(new_n716), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n961));
  NAND2_X1  g760(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n961), .B(new_n962), .ZN(G1351gat));
  INV_X1    g762(.A(G197gat), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n932), .A2(new_n934), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n697), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n965), .A2(new_n596), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n964), .B1(new_n968), .B2(KEYINPUT123), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n969), .B1(KEYINPUT123), .B2(new_n968), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n514), .A2(new_n480), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n948), .A2(new_n949), .A3(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n973), .A2(new_n964), .A3(new_n596), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n970), .A2(new_n974), .ZN(G1352gat));
  OR3_X1    g774(.A1(new_n972), .A2(G204gat), .A3(new_n681), .ZN(new_n976));
  OR2_X1    g775(.A1(new_n976), .A2(KEYINPUT124), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(KEYINPUT124), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT62), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n965), .A2(new_n708), .A3(new_n967), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(G204gat), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n977), .A2(KEYINPUT62), .A3(new_n978), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(G1353gat));
  NAND3_X1  g784(.A1(new_n973), .A2(new_n217), .A3(new_n659), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n965), .A2(new_n659), .A3(new_n967), .ZN(new_n987));
  AND3_X1   g786(.A1(new_n987), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n988));
  AOI21_X1  g787(.A(KEYINPUT63), .B1(new_n987), .B2(G211gat), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(G1354gat));
  NAND4_X1  g789(.A1(new_n948), .A2(new_n704), .A3(new_n949), .A4(new_n971), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n991), .A2(new_n208), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT125), .ZN(new_n993));
  XNOR2_X1  g792(.A(new_n992), .B(new_n993), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n480), .B1(new_n930), .B2(KEYINPUT122), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n925), .A2(new_n926), .ZN(new_n996));
  AOI21_X1  g795(.A(KEYINPUT57), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(new_n934), .ZN(new_n998));
  OAI211_X1 g797(.A(KEYINPUT126), .B(new_n967), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  NOR2_X1   g798(.A1(new_n716), .A2(new_n443), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g800(.A(KEYINPUT126), .B1(new_n965), .B2(new_n967), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n994), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(KEYINPUT127), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT127), .ZN(new_n1005));
  OAI211_X1 g804(.A(new_n994), .B(new_n1005), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1004), .A2(new_n1006), .ZN(G1355gat));
endmodule


