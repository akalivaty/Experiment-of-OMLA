

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(G651), .A2(n573), .ZN(n795) );
  AND2_X1 U550 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U551 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  NOR2_X2 U552 ( .A1(n674), .A2(n673), .ZN(n677) );
  OR2_X1 U553 ( .A1(KEYINPUT33), .A2(n685), .ZN(n727) );
  NAND2_X1 U554 ( .A1(n607), .A2(n606), .ZN(n1005) );
  XNOR2_X2 U555 ( .A(n661), .B(KEYINPUT95), .ZN(n672) );
  NOR2_X2 U556 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X2 U557 ( .A1(n650), .A2(n649), .ZN(n660) );
  AND2_X2 U558 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U559 ( .A(n610), .B(n609), .ZN(n690) );
  INV_X1 U560 ( .A(KEYINPUT17), .ZN(n518) );
  XNOR2_X1 U561 ( .A(n514), .B(n513), .ZN(n517) );
  INV_X1 U562 ( .A(KEYINPUT23), .ZN(n513) );
  NOR2_X1 U563 ( .A1(n523), .A2(n522), .ZN(n608) );
  XOR2_X1 U564 ( .A(KEYINPUT12), .B(n599), .Z(n512) );
  NOR2_X1 U565 ( .A1(n1005), .A2(n619), .ZN(n621) );
  INV_X1 U566 ( .A(KEYINPUT92), .ZN(n629) );
  INV_X1 U567 ( .A(KEYINPUT93), .ZN(n638) );
  XNOR2_X1 U568 ( .A(n653), .B(KEYINPUT30), .ZN(n654) );
  XNOR2_X1 U569 ( .A(KEYINPUT31), .B(KEYINPUT94), .ZN(n657) );
  XNOR2_X1 U570 ( .A(n658), .B(n657), .ZN(n659) );
  NAND2_X1 U571 ( .A1(n691), .A2(n611), .ZN(n624) );
  BUF_X1 U572 ( .A(n624), .Z(n662) );
  NAND2_X1 U573 ( .A1(G8), .A2(n662), .ZN(n739) );
  NAND2_X1 U574 ( .A1(n608), .A2(G40), .ZN(n610) );
  INV_X1 U575 ( .A(G651), .ZN(n533) );
  NAND2_X1 U576 ( .A1(n746), .A2(n745), .ZN(n748) );
  BUF_X1 U577 ( .A(n608), .Z(G160) );
  XNOR2_X2 U578 ( .A(G2104), .B(KEYINPUT65), .ZN(n515) );
  NOR2_X2 U579 ( .A1(n515), .A2(G2105), .ZN(n542) );
  NAND2_X1 U580 ( .A1(n542), .A2(G101), .ZN(n514) );
  AND2_X1 U581 ( .A1(n515), .A2(G2105), .ZN(n692) );
  NAND2_X1 U582 ( .A1(n692), .A2(G125), .ZN(n516) );
  NAND2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n523) );
  XNOR2_X2 U584 ( .A(n519), .B(n518), .ZN(n695) );
  NAND2_X1 U585 ( .A1(G137), .A2(n695), .ZN(n521) );
  AND2_X1 U586 ( .A1(G2105), .A2(G2104), .ZN(n895) );
  NAND2_X1 U587 ( .A1(G113), .A2(n895), .ZN(n520) );
  NAND2_X1 U588 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U589 ( .A1(G543), .A2(n533), .ZN(n524) );
  XOR2_X1 U590 ( .A(KEYINPUT66), .B(n524), .Z(n525) );
  XNOR2_X2 U591 ( .A(KEYINPUT1), .B(n525), .ZN(n791) );
  NAND2_X1 U592 ( .A1(G63), .A2(n791), .ZN(n526) );
  XNOR2_X1 U593 ( .A(KEYINPUT75), .B(n526), .ZN(n529) );
  XOR2_X1 U594 ( .A(KEYINPUT0), .B(G543), .Z(n573) );
  NAND2_X1 U595 ( .A1(n795), .A2(G51), .ZN(n527) );
  XOR2_X1 U596 ( .A(KEYINPUT76), .B(n527), .Z(n528) );
  NOR2_X1 U597 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n530), .B(KEYINPUT6), .ZN(n538) );
  NOR2_X2 U599 ( .A1(G651), .A2(G543), .ZN(n794) );
  NAND2_X1 U600 ( .A1(G89), .A2(n794), .ZN(n531) );
  XNOR2_X1 U601 ( .A(n531), .B(KEYINPUT4), .ZN(n532) );
  XNOR2_X1 U602 ( .A(n532), .B(KEYINPUT74), .ZN(n535) );
  NOR2_X2 U603 ( .A1(n573), .A2(n533), .ZN(n790) );
  NAND2_X1 U604 ( .A1(G76), .A2(n790), .ZN(n534) );
  NAND2_X1 U605 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U606 ( .A(KEYINPUT5), .B(n536), .ZN(n537) );
  NAND2_X1 U607 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n539), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U609 ( .A1(G126), .A2(n692), .ZN(n541) );
  NAND2_X1 U610 ( .A1(G138), .A2(n695), .ZN(n540) );
  NAND2_X1 U611 ( .A1(n541), .A2(n540), .ZN(n546) );
  BUF_X2 U612 ( .A(n542), .Z(n898) );
  NAND2_X1 U613 ( .A1(G102), .A2(n898), .ZN(n544) );
  NAND2_X1 U614 ( .A1(G114), .A2(n895), .ZN(n543) );
  NAND2_X1 U615 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U616 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U617 ( .A(n547), .B(KEYINPUT82), .ZN(G164) );
  NAND2_X1 U618 ( .A1(n795), .A2(G53), .ZN(n549) );
  NAND2_X1 U619 ( .A1(G65), .A2(n791), .ZN(n548) );
  NAND2_X1 U620 ( .A1(n549), .A2(n548), .ZN(n555) );
  NAND2_X1 U621 ( .A1(n794), .A2(G91), .ZN(n550) );
  XOR2_X1 U622 ( .A(KEYINPUT69), .B(n550), .Z(n552) );
  NAND2_X1 U623 ( .A1(n790), .A2(G78), .ZN(n551) );
  NAND2_X1 U624 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U625 ( .A(KEYINPUT70), .B(n553), .ZN(n554) );
  NOR2_X1 U626 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U627 ( .A(n556), .B(KEYINPUT71), .ZN(G299) );
  NAND2_X1 U628 ( .A1(G64), .A2(n791), .ZN(n557) );
  XNOR2_X1 U629 ( .A(KEYINPUT67), .B(n557), .ZN(n563) );
  NAND2_X1 U630 ( .A1(G77), .A2(n790), .ZN(n559) );
  NAND2_X1 U631 ( .A1(G90), .A2(n794), .ZN(n558) );
  NAND2_X1 U632 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U633 ( .A(KEYINPUT68), .B(n560), .Z(n561) );
  XNOR2_X1 U634 ( .A(KEYINPUT9), .B(n561), .ZN(n562) );
  NOR2_X1 U635 ( .A1(n563), .A2(n562), .ZN(n565) );
  NAND2_X1 U636 ( .A1(n795), .A2(G52), .ZN(n564) );
  NAND2_X1 U637 ( .A1(n565), .A2(n564), .ZN(G301) );
  XOR2_X1 U638 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U639 ( .A1(G75), .A2(n790), .ZN(n566) );
  XNOR2_X1 U640 ( .A(n566), .B(KEYINPUT80), .ZN(n568) );
  NAND2_X1 U641 ( .A1(G62), .A2(n791), .ZN(n567) );
  NAND2_X1 U642 ( .A1(n568), .A2(n567), .ZN(n572) );
  NAND2_X1 U643 ( .A1(G88), .A2(n794), .ZN(n570) );
  NAND2_X1 U644 ( .A1(G50), .A2(n795), .ZN(n569) );
  NAND2_X1 U645 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U646 ( .A1(n572), .A2(n571), .ZN(G166) );
  INV_X1 U647 ( .A(G166), .ZN(G303) );
  NAND2_X1 U648 ( .A1(G87), .A2(n573), .ZN(n575) );
  NAND2_X1 U649 ( .A1(G74), .A2(G651), .ZN(n574) );
  NAND2_X1 U650 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U651 ( .A1(n791), .A2(n576), .ZN(n578) );
  NAND2_X1 U652 ( .A1(n795), .A2(G49), .ZN(n577) );
  NAND2_X1 U653 ( .A1(n578), .A2(n577), .ZN(G288) );
  NAND2_X1 U654 ( .A1(n794), .A2(G86), .ZN(n580) );
  NAND2_X1 U655 ( .A1(G61), .A2(n791), .ZN(n579) );
  NAND2_X1 U656 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n790), .A2(G73), .ZN(n581) );
  XOR2_X1 U658 ( .A(KEYINPUT2), .B(n581), .Z(n582) );
  NOR2_X1 U659 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U660 ( .A1(n795), .A2(G48), .ZN(n584) );
  NAND2_X1 U661 ( .A1(n585), .A2(n584), .ZN(G305) );
  AND2_X1 U662 ( .A1(G60), .A2(n791), .ZN(n589) );
  NAND2_X1 U663 ( .A1(G72), .A2(n790), .ZN(n587) );
  NAND2_X1 U664 ( .A1(G85), .A2(n794), .ZN(n586) );
  NAND2_X1 U665 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U666 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n795), .A2(G47), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(G290) );
  NAND2_X1 U669 ( .A1(n790), .A2(G79), .ZN(n593) );
  NAND2_X1 U670 ( .A1(G66), .A2(n791), .ZN(n592) );
  NAND2_X1 U671 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U672 ( .A1(G92), .A2(n794), .ZN(n595) );
  NAND2_X1 U673 ( .A1(G54), .A2(n795), .ZN(n594) );
  NAND2_X1 U674 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U675 ( .A1(n597), .A2(n596), .ZN(n618) );
  XOR2_X1 U676 ( .A(KEYINPUT15), .B(n618), .Z(n1018) );
  NAND2_X1 U677 ( .A1(n790), .A2(G68), .ZN(n598) );
  XNOR2_X1 U678 ( .A(KEYINPUT73), .B(n598), .ZN(n600) );
  NAND2_X1 U679 ( .A1(n794), .A2(G81), .ZN(n599) );
  NOR2_X1 U680 ( .A1(n600), .A2(n512), .ZN(n601) );
  XNOR2_X1 U681 ( .A(n601), .B(KEYINPUT13), .ZN(n605) );
  XOR2_X1 U682 ( .A(KEYINPUT14), .B(KEYINPUT72), .Z(n603) );
  NAND2_X1 U683 ( .A1(G56), .A2(n791), .ZN(n602) );
  XNOR2_X1 U684 ( .A(n603), .B(n602), .ZN(n604) );
  NOR2_X1 U685 ( .A1(n605), .A2(n604), .ZN(n607) );
  NAND2_X1 U686 ( .A1(n795), .A2(G43), .ZN(n606) );
  NOR2_X1 U687 ( .A1(G1384), .A2(G164), .ZN(n691) );
  INV_X1 U688 ( .A(KEYINPUT83), .ZN(n609) );
  XNOR2_X1 U689 ( .A(KEYINPUT89), .B(n690), .ZN(n611) );
  XNOR2_X1 U690 ( .A(G1996), .B(KEYINPUT91), .ZN(n925) );
  NOR2_X1 U691 ( .A1(n624), .A2(n925), .ZN(n613) );
  INV_X1 U692 ( .A(KEYINPUT26), .ZN(n612) );
  NAND2_X1 U693 ( .A1(n613), .A2(n612), .ZN(n615) );
  OR2_X1 U694 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n623) );
  NAND2_X1 U696 ( .A1(n624), .A2(G1341), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n623), .A2(n620), .ZN(n616) );
  NOR2_X1 U698 ( .A1(n1005), .A2(n616), .ZN(n617) );
  NOR2_X1 U699 ( .A1(n1018), .A2(n617), .ZN(n632) );
  XNOR2_X1 U700 ( .A(KEYINPUT15), .B(n618), .ZN(n619) );
  AND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n628) );
  INV_X1 U703 ( .A(n624), .ZN(n645) );
  NOR2_X1 U704 ( .A1(n645), .A2(G1348), .ZN(n626) );
  NOR2_X1 U705 ( .A1(G2067), .A2(n662), .ZN(n625) );
  NOR2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n630) );
  XNOR2_X1 U708 ( .A(n630), .B(n629), .ZN(n631) );
  NOR2_X1 U709 ( .A1(n632), .A2(n631), .ZN(n637) );
  NAND2_X1 U710 ( .A1(n645), .A2(G2072), .ZN(n633) );
  XOR2_X1 U711 ( .A(KEYINPUT27), .B(n633), .Z(n635) );
  NAND2_X1 U712 ( .A1(G1956), .A2(n662), .ZN(n634) );
  NAND2_X1 U713 ( .A1(n635), .A2(n634), .ZN(n640) );
  NOR2_X1 U714 ( .A1(G299), .A2(n640), .ZN(n636) );
  NOR2_X1 U715 ( .A1(n637), .A2(n636), .ZN(n639) );
  XNOR2_X1 U716 ( .A(n639), .B(n638), .ZN(n643) );
  NAND2_X1 U717 ( .A1(G299), .A2(n640), .ZN(n641) );
  XOR2_X1 U718 ( .A(KEYINPUT28), .B(n641), .Z(n642) );
  NOR2_X1 U719 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U720 ( .A(n644), .B(KEYINPUT29), .ZN(n650) );
  NAND2_X1 U721 ( .A1(G1961), .A2(n662), .ZN(n647) );
  XOR2_X1 U722 ( .A(KEYINPUT25), .B(G2078), .Z(n931) );
  NAND2_X1 U723 ( .A1(n645), .A2(n931), .ZN(n646) );
  NAND2_X1 U724 ( .A1(n647), .A2(n646), .ZN(n651) );
  NOR2_X1 U725 ( .A1(G301), .A2(n651), .ZN(n648) );
  XOR2_X1 U726 ( .A(KEYINPUT90), .B(n648), .Z(n649) );
  AND2_X1 U727 ( .A1(G301), .A2(n651), .ZN(n656) );
  NOR2_X1 U728 ( .A1(G1966), .A2(n739), .ZN(n673) );
  NOR2_X1 U729 ( .A1(G2084), .A2(n662), .ZN(n675) );
  NOR2_X1 U730 ( .A1(n673), .A2(n675), .ZN(n652) );
  NAND2_X1 U731 ( .A1(G8), .A2(n652), .ZN(n653) );
  NOR2_X1 U732 ( .A1(n654), .A2(G168), .ZN(n655) );
  NOR2_X1 U733 ( .A1(n656), .A2(n655), .ZN(n658) );
  NAND2_X1 U734 ( .A1(n672), .A2(G286), .ZN(n670) );
  INV_X1 U735 ( .A(G8), .ZN(n668) );
  NOR2_X1 U736 ( .A1(G2090), .A2(n662), .ZN(n663) );
  XNOR2_X1 U737 ( .A(n663), .B(KEYINPUT96), .ZN(n665) );
  NOR2_X1 U738 ( .A1(n739), .A2(G1971), .ZN(n664) );
  NOR2_X1 U739 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U740 ( .A1(n666), .A2(G303), .ZN(n667) );
  OR2_X1 U741 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X2 U742 ( .A(n671), .B(KEYINPUT32), .ZN(n730) );
  INV_X1 U743 ( .A(n672), .ZN(n674) );
  NAND2_X1 U744 ( .A1(G8), .A2(n675), .ZN(n676) );
  NAND2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n728) );
  NAND2_X1 U746 ( .A1(G1976), .A2(G288), .ZN(n1017) );
  INV_X1 U747 ( .A(n739), .ZN(n733) );
  NAND2_X1 U748 ( .A1(n1017), .A2(n733), .ZN(n681) );
  INV_X1 U749 ( .A(n681), .ZN(n678) );
  AND2_X1 U750 ( .A1(n728), .A2(n678), .ZN(n679) );
  NAND2_X1 U751 ( .A1(n730), .A2(n679), .ZN(n683) );
  NOR2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n686) );
  NOR2_X1 U753 ( .A1(G1971), .A2(G303), .ZN(n680) );
  NOR2_X1 U754 ( .A1(n686), .A2(n680), .ZN(n1012) );
  OR2_X1 U755 ( .A1(n681), .A2(n1012), .ZN(n682) );
  NAND2_X1 U756 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U757 ( .A(n684), .B(KEYINPUT64), .ZN(n685) );
  NAND2_X1 U758 ( .A1(n686), .A2(KEYINPUT33), .ZN(n687) );
  NOR2_X1 U759 ( .A1(n687), .A2(n739), .ZN(n689) );
  XOR2_X1 U760 ( .A(G1981), .B(G305), .Z(n1002) );
  INV_X1 U761 ( .A(n1002), .ZN(n688) );
  NOR2_X1 U762 ( .A1(n689), .A2(n688), .ZN(n725) );
  NOR2_X1 U763 ( .A1(n691), .A2(n690), .ZN(n761) );
  NAND2_X1 U764 ( .A1(G119), .A2(n692), .ZN(n694) );
  NAND2_X1 U765 ( .A1(G95), .A2(n898), .ZN(n693) );
  NAND2_X1 U766 ( .A1(n694), .A2(n693), .ZN(n699) );
  NAND2_X1 U767 ( .A1(G131), .A2(n695), .ZN(n697) );
  NAND2_X1 U768 ( .A1(G107), .A2(n895), .ZN(n696) );
  NAND2_X1 U769 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U770 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U771 ( .A(KEYINPUT86), .B(n700), .Z(n907) );
  NAND2_X1 U772 ( .A1(G1991), .A2(n907), .ZN(n709) );
  NAND2_X1 U773 ( .A1(G141), .A2(n695), .ZN(n702) );
  NAND2_X1 U774 ( .A1(G117), .A2(n895), .ZN(n701) );
  NAND2_X1 U775 ( .A1(n702), .A2(n701), .ZN(n705) );
  NAND2_X1 U776 ( .A1(n898), .A2(G105), .ZN(n703) );
  XOR2_X1 U777 ( .A(KEYINPUT38), .B(n703), .Z(n704) );
  NOR2_X1 U778 ( .A1(n705), .A2(n704), .ZN(n707) );
  NAND2_X1 U779 ( .A1(n692), .A2(G129), .ZN(n706) );
  NAND2_X1 U780 ( .A1(n707), .A2(n706), .ZN(n882) );
  NAND2_X1 U781 ( .A1(G1996), .A2(n882), .ZN(n708) );
  NAND2_X1 U782 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U783 ( .A(KEYINPUT87), .B(n710), .Z(n987) );
  NAND2_X1 U784 ( .A1(n761), .A2(n987), .ZN(n749) );
  NAND2_X1 U785 ( .A1(G104), .A2(n898), .ZN(n712) );
  NAND2_X1 U786 ( .A1(G140), .A2(n695), .ZN(n711) );
  NAND2_X1 U787 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U788 ( .A(KEYINPUT34), .B(n713), .ZN(n719) );
  NAND2_X1 U789 ( .A1(G128), .A2(n692), .ZN(n715) );
  NAND2_X1 U790 ( .A1(G116), .A2(n895), .ZN(n714) );
  NAND2_X1 U791 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U792 ( .A(KEYINPUT35), .B(n716), .ZN(n717) );
  XNOR2_X1 U793 ( .A(KEYINPUT85), .B(n717), .ZN(n718) );
  NOR2_X1 U794 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U795 ( .A(KEYINPUT36), .B(n720), .ZN(n908) );
  XNOR2_X1 U796 ( .A(G2067), .B(KEYINPUT37), .ZN(n758) );
  NOR2_X1 U797 ( .A1(n908), .A2(n758), .ZN(n978) );
  NAND2_X1 U798 ( .A1(n761), .A2(n978), .ZN(n756) );
  NAND2_X1 U799 ( .A1(n749), .A2(n756), .ZN(n721) );
  XNOR2_X1 U800 ( .A(n721), .B(KEYINPUT88), .ZN(n724) );
  XNOR2_X1 U801 ( .A(G1986), .B(G290), .ZN(n1010) );
  NAND2_X1 U802 ( .A1(n761), .A2(n1010), .ZN(n722) );
  XOR2_X1 U803 ( .A(KEYINPUT84), .B(n722), .Z(n723) );
  NOR2_X1 U804 ( .A1(n724), .A2(n723), .ZN(n742) );
  AND2_X1 U805 ( .A1(n725), .A2(n742), .ZN(n726) );
  NAND2_X1 U806 ( .A1(n727), .A2(n726), .ZN(n746) );
  AND2_X1 U807 ( .A1(n728), .A2(n739), .ZN(n729) );
  NAND2_X1 U808 ( .A1(n730), .A2(n729), .ZN(n735) );
  NOR2_X1 U809 ( .A1(G2090), .A2(G303), .ZN(n731) );
  NAND2_X1 U810 ( .A1(G8), .A2(n731), .ZN(n732) );
  OR2_X1 U811 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U812 ( .A(n736), .B(KEYINPUT97), .ZN(n741) );
  NOR2_X1 U813 ( .A1(G1981), .A2(G305), .ZN(n737) );
  XOR2_X1 U814 ( .A(n737), .B(KEYINPUT24), .Z(n738) );
  NOR2_X1 U815 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U816 ( .A1(n741), .A2(n740), .ZN(n744) );
  INV_X1 U817 ( .A(n742), .ZN(n743) );
  OR2_X2 U818 ( .A1(n744), .A2(n743), .ZN(n745) );
  INV_X1 U819 ( .A(KEYINPUT98), .ZN(n747) );
  XNOR2_X1 U820 ( .A(n748), .B(n747), .ZN(n763) );
  NOR2_X1 U821 ( .A1(G1996), .A2(n882), .ZN(n990) );
  INV_X1 U822 ( .A(n749), .ZN(n753) );
  NOR2_X1 U823 ( .A1(G1991), .A2(n907), .ZN(n983) );
  NOR2_X1 U824 ( .A1(G1986), .A2(G290), .ZN(n750) );
  XOR2_X1 U825 ( .A(n750), .B(KEYINPUT99), .Z(n751) );
  NOR2_X1 U826 ( .A1(n983), .A2(n751), .ZN(n752) );
  NOR2_X1 U827 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U828 ( .A1(n990), .A2(n754), .ZN(n755) );
  XNOR2_X1 U829 ( .A(n755), .B(KEYINPUT39), .ZN(n757) );
  NAND2_X1 U830 ( .A1(n757), .A2(n756), .ZN(n759) );
  NAND2_X1 U831 ( .A1(n908), .A2(n758), .ZN(n977) );
  NAND2_X1 U832 ( .A1(n759), .A2(n977), .ZN(n760) );
  NAND2_X1 U833 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U834 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U835 ( .A(n764), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U836 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U837 ( .A1(G123), .A2(n692), .ZN(n765) );
  XNOR2_X1 U838 ( .A(n765), .B(KEYINPUT18), .ZN(n772) );
  NAND2_X1 U839 ( .A1(G99), .A2(n898), .ZN(n767) );
  NAND2_X1 U840 ( .A1(G135), .A2(n695), .ZN(n766) );
  NAND2_X1 U841 ( .A1(n767), .A2(n766), .ZN(n770) );
  NAND2_X1 U842 ( .A1(G111), .A2(n895), .ZN(n768) );
  XNOR2_X1 U843 ( .A(KEYINPUT79), .B(n768), .ZN(n769) );
  NOR2_X1 U844 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U845 ( .A1(n772), .A2(n771), .ZN(n984) );
  XNOR2_X1 U846 ( .A(G2096), .B(n984), .ZN(n773) );
  OR2_X1 U847 ( .A1(G2100), .A2(n773), .ZN(G156) );
  INV_X1 U848 ( .A(G57), .ZN(G237) );
  INV_X1 U849 ( .A(G132), .ZN(G219) );
  INV_X1 U850 ( .A(G82), .ZN(G220) );
  NAND2_X1 U851 ( .A1(G7), .A2(G661), .ZN(n774) );
  XNOR2_X1 U852 ( .A(n774), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U853 ( .A(G223), .ZN(n836) );
  NAND2_X1 U854 ( .A1(n836), .A2(G567), .ZN(n775) );
  XOR2_X1 U855 ( .A(KEYINPUT11), .B(n775), .Z(G234) );
  INV_X1 U856 ( .A(G860), .ZN(n789) );
  OR2_X1 U857 ( .A1(n1005), .A2(n789), .ZN(G153) );
  NAND2_X1 U858 ( .A1(G868), .A2(G301), .ZN(n777) );
  OR2_X1 U859 ( .A1(n1018), .A2(G868), .ZN(n776) );
  NAND2_X1 U860 ( .A1(n777), .A2(n776), .ZN(G284) );
  INV_X1 U861 ( .A(G868), .ZN(n778) );
  NOR2_X1 U862 ( .A1(G286), .A2(n778), .ZN(n779) );
  XOR2_X1 U863 ( .A(KEYINPUT77), .B(n779), .Z(n781) );
  NOR2_X1 U864 ( .A1(G868), .A2(G299), .ZN(n780) );
  NOR2_X1 U865 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U866 ( .A(KEYINPUT78), .B(n782), .ZN(G297) );
  NAND2_X1 U867 ( .A1(n789), .A2(G559), .ZN(n783) );
  NAND2_X1 U868 ( .A1(n783), .A2(n1018), .ZN(n784) );
  XNOR2_X1 U869 ( .A(n784), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U870 ( .A1(G868), .A2(n1005), .ZN(n787) );
  NAND2_X1 U871 ( .A1(G868), .A2(n1018), .ZN(n785) );
  NOR2_X1 U872 ( .A1(G559), .A2(n785), .ZN(n786) );
  NOR2_X1 U873 ( .A1(n787), .A2(n786), .ZN(G282) );
  NAND2_X1 U874 ( .A1(G559), .A2(n1018), .ZN(n788) );
  XOR2_X1 U875 ( .A(n1005), .B(n788), .Z(n806) );
  NAND2_X1 U876 ( .A1(n789), .A2(n806), .ZN(n800) );
  NAND2_X1 U877 ( .A1(n790), .A2(G80), .ZN(n793) );
  NAND2_X1 U878 ( .A1(G67), .A2(n791), .ZN(n792) );
  NAND2_X1 U879 ( .A1(n793), .A2(n792), .ZN(n799) );
  NAND2_X1 U880 ( .A1(G93), .A2(n794), .ZN(n797) );
  NAND2_X1 U881 ( .A1(G55), .A2(n795), .ZN(n796) );
  NAND2_X1 U882 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U883 ( .A1(n799), .A2(n798), .ZN(n808) );
  XOR2_X1 U884 ( .A(n800), .B(n808), .Z(G145) );
  XNOR2_X1 U885 ( .A(KEYINPUT19), .B(G288), .ZN(n805) );
  XNOR2_X1 U886 ( .A(G166), .B(G305), .ZN(n801) );
  XNOR2_X1 U887 ( .A(n801), .B(G299), .ZN(n802) );
  XNOR2_X1 U888 ( .A(n808), .B(n802), .ZN(n803) );
  XNOR2_X1 U889 ( .A(n803), .B(G290), .ZN(n804) );
  XNOR2_X1 U890 ( .A(n805), .B(n804), .ZN(n848) );
  XNOR2_X1 U891 ( .A(n806), .B(n848), .ZN(n807) );
  NAND2_X1 U892 ( .A1(n807), .A2(G868), .ZN(n810) );
  OR2_X1 U893 ( .A1(G868), .A2(n808), .ZN(n809) );
  NAND2_X1 U894 ( .A1(n810), .A2(n809), .ZN(G295) );
  NAND2_X1 U895 ( .A1(G2084), .A2(G2078), .ZN(n811) );
  XOR2_X1 U896 ( .A(KEYINPUT20), .B(n811), .Z(n812) );
  NAND2_X1 U897 ( .A1(G2090), .A2(n812), .ZN(n813) );
  XNOR2_X1 U898 ( .A(KEYINPUT21), .B(n813), .ZN(n814) );
  NAND2_X1 U899 ( .A1(n814), .A2(G2072), .ZN(G158) );
  XOR2_X1 U900 ( .A(KEYINPUT81), .B(G44), .Z(n815) );
  XNOR2_X1 U901 ( .A(KEYINPUT3), .B(n815), .ZN(G218) );
  NOR2_X1 U902 ( .A1(G220), .A2(G219), .ZN(n816) );
  XOR2_X1 U903 ( .A(KEYINPUT22), .B(n816), .Z(n817) );
  NOR2_X1 U904 ( .A1(G218), .A2(n817), .ZN(n818) );
  NAND2_X1 U905 ( .A1(G96), .A2(n818), .ZN(n844) );
  NAND2_X1 U906 ( .A1(G2106), .A2(n844), .ZN(n822) );
  NAND2_X1 U907 ( .A1(G120), .A2(G69), .ZN(n819) );
  NOR2_X1 U908 ( .A1(G237), .A2(n819), .ZN(n820) );
  NAND2_X1 U909 ( .A1(G108), .A2(n820), .ZN(n843) );
  NAND2_X1 U910 ( .A1(G567), .A2(n843), .ZN(n821) );
  NAND2_X1 U911 ( .A1(n822), .A2(n821), .ZN(n914) );
  NAND2_X1 U912 ( .A1(G483), .A2(G661), .ZN(n823) );
  NOR2_X1 U913 ( .A1(n914), .A2(n823), .ZN(n841) );
  NAND2_X1 U914 ( .A1(n841), .A2(G36), .ZN(G176) );
  XNOR2_X1 U915 ( .A(G1341), .B(G1348), .ZN(n824) );
  XNOR2_X1 U916 ( .A(n824), .B(G2427), .ZN(n834) );
  XOR2_X1 U917 ( .A(G2446), .B(KEYINPUT100), .Z(n826) );
  XNOR2_X1 U918 ( .A(G2430), .B(G2451), .ZN(n825) );
  XNOR2_X1 U919 ( .A(n826), .B(n825), .ZN(n830) );
  XOR2_X1 U920 ( .A(G2435), .B(KEYINPUT101), .Z(n828) );
  XNOR2_X1 U921 ( .A(G2438), .B(G2454), .ZN(n827) );
  XNOR2_X1 U922 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U923 ( .A(n830), .B(n829), .Z(n832) );
  XNOR2_X1 U924 ( .A(KEYINPUT102), .B(G2443), .ZN(n831) );
  XNOR2_X1 U925 ( .A(n832), .B(n831), .ZN(n833) );
  XNOR2_X1 U926 ( .A(n834), .B(n833), .ZN(n835) );
  NAND2_X1 U927 ( .A1(n835), .A2(G14), .ZN(n917) );
  XNOR2_X1 U928 ( .A(KEYINPUT103), .B(n917), .ZN(G401) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n836), .ZN(G217) );
  NAND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n837) );
  XOR2_X1 U931 ( .A(KEYINPUT104), .B(n837), .Z(n838) );
  NAND2_X1 U932 ( .A1(n838), .A2(G661), .ZN(n839) );
  XOR2_X1 U933 ( .A(KEYINPUT105), .B(n839), .Z(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n840) );
  XNOR2_X1 U935 ( .A(KEYINPUT106), .B(n840), .ZN(n842) );
  NAND2_X1 U936 ( .A1(n842), .A2(n841), .ZN(G188) );
  XNOR2_X1 U937 ( .A(G96), .B(KEYINPUT107), .ZN(G221) );
  XOR2_X1 U938 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  INV_X1 U940 ( .A(G120), .ZN(G236) );
  NOR2_X1 U941 ( .A1(n844), .A2(n843), .ZN(n845) );
  XNOR2_X1 U942 ( .A(n845), .B(KEYINPUT109), .ZN(G261) );
  INV_X1 U943 ( .A(G261), .ZN(G325) );
  INV_X1 U944 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U945 ( .A(n1005), .B(KEYINPUT119), .ZN(n847) );
  XNOR2_X1 U946 ( .A(G171), .B(n1018), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n850) );
  XOR2_X1 U948 ( .A(G286), .B(n848), .Z(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n851) );
  NOR2_X1 U950 ( .A1(G37), .A2(n851), .ZN(G397) );
  XOR2_X1 U951 ( .A(G2096), .B(G2090), .Z(n853) );
  XNOR2_X1 U952 ( .A(G2067), .B(G2072), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n863) );
  XOR2_X1 U954 ( .A(KEYINPUT42), .B(KEYINPUT43), .Z(n855) );
  XNOR2_X1 U955 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U957 ( .A(G2100), .B(G2678), .Z(n857) );
  XNOR2_X1 U958 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U960 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U961 ( .A(G2084), .B(G2078), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U963 ( .A(n863), .B(n862), .Z(G227) );
  XOR2_X1 U964 ( .A(G1961), .B(G1971), .Z(n865) );
  XNOR2_X1 U965 ( .A(G1986), .B(G1976), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U967 ( .A(n866), .B(G2474), .Z(n868) );
  XNOR2_X1 U968 ( .A(G1981), .B(G1966), .ZN(n867) );
  XNOR2_X1 U969 ( .A(n868), .B(n867), .ZN(n872) );
  XOR2_X1 U970 ( .A(KEYINPUT41), .B(G1956), .Z(n870) );
  XNOR2_X1 U971 ( .A(G1996), .B(G1991), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U973 ( .A(n872), .B(n871), .ZN(G229) );
  NAND2_X1 U974 ( .A1(G100), .A2(n898), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G112), .A2(n895), .ZN(n873) );
  NAND2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n881) );
  NAND2_X1 U977 ( .A1(n695), .A2(G136), .ZN(n875) );
  XNOR2_X1 U978 ( .A(KEYINPUT115), .B(n875), .ZN(n878) );
  NAND2_X1 U979 ( .A1(n692), .A2(G124), .ZN(n876) );
  XOR2_X1 U980 ( .A(KEYINPUT44), .B(n876), .Z(n877) );
  NOR2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U982 ( .A(KEYINPUT116), .B(n879), .Z(n880) );
  NOR2_X1 U983 ( .A1(n881), .A2(n880), .ZN(G162) );
  XNOR2_X1 U984 ( .A(G160), .B(n882), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n883), .B(n984), .ZN(n887) );
  XOR2_X1 U986 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n885) );
  XNOR2_X1 U987 ( .A(KEYINPUT118), .B(KEYINPUT117), .ZN(n884) );
  XNOR2_X1 U988 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U989 ( .A(n887), .B(n886), .Z(n906) );
  NAND2_X1 U990 ( .A1(G103), .A2(n898), .ZN(n889) );
  NAND2_X1 U991 ( .A1(G139), .A2(n695), .ZN(n888) );
  NAND2_X1 U992 ( .A1(n889), .A2(n888), .ZN(n894) );
  NAND2_X1 U993 ( .A1(G127), .A2(n692), .ZN(n891) );
  NAND2_X1 U994 ( .A1(G115), .A2(n895), .ZN(n890) );
  NAND2_X1 U995 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U996 ( .A(KEYINPUT47), .B(n892), .Z(n893) );
  NOR2_X1 U997 ( .A1(n894), .A2(n893), .ZN(n971) );
  NAND2_X1 U998 ( .A1(G130), .A2(n692), .ZN(n897) );
  NAND2_X1 U999 ( .A1(G118), .A2(n895), .ZN(n896) );
  NAND2_X1 U1000 ( .A1(n897), .A2(n896), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(G106), .A2(n898), .ZN(n900) );
  NAND2_X1 U1002 ( .A1(G142), .A2(n695), .ZN(n899) );
  NAND2_X1 U1003 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U1004 ( .A(KEYINPUT45), .B(n901), .Z(n902) );
  NOR2_X1 U1005 ( .A1(n903), .A2(n902), .ZN(n904) );
  XNOR2_X1 U1006 ( .A(n971), .B(n904), .ZN(n905) );
  XNOR2_X1 U1007 ( .A(n906), .B(n905), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n907), .B(G164), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(G162), .B(n910), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(n912), .B(n911), .ZN(n913) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n913), .ZN(G395) );
  XOR2_X1 U1013 ( .A(KEYINPUT110), .B(n914), .Z(G319) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n915) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n915), .ZN(n916) );
  NOR2_X1 U1016 ( .A1(G397), .A2(n916), .ZN(n921) );
  NAND2_X1 U1017 ( .A1(G319), .A2(n917), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(KEYINPUT120), .B(n918), .ZN(n919) );
  NOR2_X1 U1019 ( .A1(G395), .A2(n919), .ZN(n920) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1023 ( .A(G1991), .B(G25), .ZN(n923) );
  XNOR2_X1 U1024 ( .A(G33), .B(G2072), .ZN(n922) );
  NOR2_X1 U1025 ( .A1(n923), .A2(n922), .ZN(n930) );
  XOR2_X1 U1026 ( .A(G2067), .B(G26), .Z(n924) );
  NAND2_X1 U1027 ( .A1(n924), .A2(G28), .ZN(n928) );
  XOR2_X1 U1028 ( .A(G32), .B(n925), .Z(n926) );
  XNOR2_X1 U1029 ( .A(KEYINPUT124), .B(n926), .ZN(n927) );
  NOR2_X1 U1030 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(G27), .B(n931), .ZN(n932) );
  NOR2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1034 ( .A(KEYINPUT53), .B(n934), .Z(n937) );
  XOR2_X1 U1035 ( .A(G34), .B(KEYINPUT54), .Z(n935) );
  XNOR2_X1 U1036 ( .A(G2084), .B(n935), .ZN(n936) );
  NAND2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n939) );
  XNOR2_X1 U1038 ( .A(G35), .B(G2090), .ZN(n938) );
  NOR2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n964) );
  NAND2_X1 U1040 ( .A1(KEYINPUT55), .A2(n964), .ZN(n940) );
  NAND2_X1 U1041 ( .A1(G11), .A2(n940), .ZN(n970) );
  XOR2_X1 U1042 ( .A(G16), .B(KEYINPUT126), .Z(n963) );
  XOR2_X1 U1043 ( .A(G1348), .B(KEYINPUT59), .Z(n941) );
  XNOR2_X1 U1044 ( .A(G4), .B(n941), .ZN(n943) );
  XNOR2_X1 U1045 ( .A(G6), .B(G1981), .ZN(n942) );
  NOR2_X1 U1046 ( .A1(n943), .A2(n942), .ZN(n947) );
  XNOR2_X1 U1047 ( .A(G1341), .B(G19), .ZN(n945) );
  XNOR2_X1 U1048 ( .A(G20), .B(G1956), .ZN(n944) );
  NOR2_X1 U1049 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1050 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1051 ( .A(n948), .B(KEYINPUT60), .ZN(n949) );
  XNOR2_X1 U1052 ( .A(KEYINPUT127), .B(n949), .ZN(n953) );
  XNOR2_X1 U1053 ( .A(G1966), .B(G21), .ZN(n951) );
  XNOR2_X1 U1054 ( .A(G5), .B(G1961), .ZN(n950) );
  NOR2_X1 U1055 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1056 ( .A1(n953), .A2(n952), .ZN(n960) );
  XNOR2_X1 U1057 ( .A(G1976), .B(G23), .ZN(n955) );
  XNOR2_X1 U1058 ( .A(G1971), .B(G22), .ZN(n954) );
  NOR2_X1 U1059 ( .A1(n955), .A2(n954), .ZN(n957) );
  XOR2_X1 U1060 ( .A(G1986), .B(G24), .Z(n956) );
  NAND2_X1 U1061 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1062 ( .A(KEYINPUT58), .B(n958), .ZN(n959) );
  NOR2_X1 U1063 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1064 ( .A(n961), .B(KEYINPUT61), .ZN(n962) );
  NAND2_X1 U1065 ( .A1(n963), .A2(n962), .ZN(n968) );
  INV_X1 U1066 ( .A(n964), .ZN(n966) );
  NOR2_X1 U1067 ( .A1(G29), .A2(KEYINPUT55), .ZN(n965) );
  NAND2_X1 U1068 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1069 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1070 ( .A1(n970), .A2(n969), .ZN(n1001) );
  XOR2_X1 U1071 ( .A(G2072), .B(n971), .Z(n972) );
  XNOR2_X1 U1072 ( .A(KEYINPUT122), .B(n972), .ZN(n975) );
  XNOR2_X1 U1073 ( .A(G2078), .B(G164), .ZN(n973) );
  XNOR2_X1 U1074 ( .A(KEYINPUT123), .B(n973), .ZN(n974) );
  NOR2_X1 U1075 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1076 ( .A(KEYINPUT50), .B(n976), .ZN(n981) );
  INV_X1 U1077 ( .A(n977), .ZN(n979) );
  NOR2_X1 U1078 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1079 ( .A1(n981), .A2(n980), .ZN(n995) );
  XOR2_X1 U1080 ( .A(G160), .B(G2084), .Z(n982) );
  NOR2_X1 U1081 ( .A1(n983), .A2(n982), .ZN(n985) );
  NAND2_X1 U1082 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1083 ( .A1(n987), .A2(n986), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(G2090), .B(G162), .ZN(n988) );
  XNOR2_X1 U1085 ( .A(n988), .B(KEYINPUT121), .ZN(n989) );
  NOR2_X1 U1086 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1087 ( .A(KEYINPUT51), .B(n991), .Z(n992) );
  NAND2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1090 ( .A(KEYINPUT52), .B(n996), .ZN(n998) );
  INV_X1 U1091 ( .A(KEYINPUT55), .ZN(n997) );
  NAND2_X1 U1092 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1093 ( .A1(n999), .A2(G29), .ZN(n1000) );
  NAND2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1028) );
  XOR2_X1 U1095 ( .A(KEYINPUT56), .B(G16), .Z(n1026) );
  XNOR2_X1 U1096 ( .A(G1966), .B(G168), .ZN(n1003) );
  NAND2_X1 U1097 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1098 ( .A(n1004), .B(KEYINPUT57), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(n1005), .B(G1341), .ZN(n1007) );
  XNOR2_X1 U1100 ( .A(G299), .B(G1956), .ZN(n1006) );
  NOR2_X1 U1101 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1102 ( .A1(n1009), .A2(n1008), .ZN(n1024) );
  INV_X1 U1103 ( .A(n1010), .ZN(n1011) );
  NAND2_X1 U1104 ( .A1(n1012), .A2(n1011), .ZN(n1015) );
  XOR2_X1 U1105 ( .A(G1961), .B(G301), .Z(n1013) );
  XNOR2_X1 U1106 ( .A(KEYINPUT125), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1107 ( .A1(n1015), .A2(n1014), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(G1971), .A2(G303), .ZN(n1016) );
  NAND2_X1 U1109 ( .A1(n1017), .A2(n1016), .ZN(n1020) );
  XOR2_X1 U1110 ( .A(n1018), .B(G1348), .Z(n1019) );
  NOR2_X1 U1111 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1112 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1116 ( .A(n1029), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

