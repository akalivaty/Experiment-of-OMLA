//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT64), .B1(new_n188), .B2(G116), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n188), .A2(G116), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  XOR2_X1   g009(.A(KEYINPUT2), .B(G113), .Z(new_n196));
  XOR2_X1   g010(.A(new_n195), .B(new_n196), .Z(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G137), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT11), .A3(G134), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(G137), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n200), .A2(new_n202), .A3(new_n203), .A4(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n201), .A2(G134), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n199), .A2(G137), .ZN(new_n207));
  OAI21_X1  g021(.A(G131), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT1), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  AND4_X1   g028(.A1(new_n210), .A2(new_n212), .A3(new_n214), .A4(G128), .ZN(new_n215));
  XNOR2_X1  g029(.A(G143), .B(G146), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(G128), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n214), .A2(new_n210), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n209), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT0), .A4(G128), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT0), .B(G128), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n222), .B1(new_n216), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n200), .A2(new_n204), .A3(new_n202), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G131), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n224), .B1(new_n226), .B2(new_n205), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n221), .A2(new_n227), .A3(KEYINPUT30), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT30), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n209), .A2(KEYINPUT65), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n216), .A2(new_n210), .A3(G128), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n231), .B(new_n220), .C1(G128), .C2(new_n216), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n205), .A2(new_n208), .A3(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n230), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n224), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n226), .A2(new_n205), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n229), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n197), .B1(new_n228), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n235), .A2(new_n238), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(new_n197), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n244));
  INV_X1    g058(.A(G237), .ZN(new_n245));
  INV_X1    g059(.A(G953), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n246), .A3(G210), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n244), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G101), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n248), .B(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n240), .A2(new_n243), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT31), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n251), .A2(KEYINPUT67), .A3(KEYINPUT31), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT28), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n242), .B(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n197), .B1(new_n227), .B2(new_n221), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n250), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n232), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n238), .B(new_n229), .C1(new_n264), .C2(new_n209), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n205), .A2(new_n208), .A3(new_n233), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n233), .B1(new_n205), .B2(new_n208), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n227), .B1(new_n268), .B2(new_n232), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n265), .B1(new_n269), .B2(new_n229), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n242), .B1(new_n270), .B2(new_n197), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT31), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n271), .A2(KEYINPUT68), .A3(new_n272), .A4(new_n250), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n240), .A2(new_n243), .A3(new_n272), .A4(new_n250), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT68), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n256), .A2(new_n257), .A3(new_n263), .A4(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n254), .A2(new_n255), .B1(new_n276), .B2(new_n273), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n257), .B1(new_n280), .B2(new_n263), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n187), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT32), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n187), .ZN(new_n285));
  INV_X1    g099(.A(new_n255), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT67), .B1(new_n251), .B2(KEYINPUT31), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n277), .B(new_n263), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT69), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n285), .B1(new_n289), .B2(new_n278), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT32), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n261), .A2(new_n262), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n271), .A2(new_n250), .ZN(new_n293));
  NOR3_X1   g107(.A1(new_n292), .A2(KEYINPUT29), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT70), .B(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n241), .A2(new_n197), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n259), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n250), .A2(KEYINPUT29), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n296), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G472), .B1(new_n294), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n284), .A2(new_n291), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(G125), .B(G140), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT16), .ZN(new_n304));
  INV_X1    g118(.A(G140), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G125), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n304), .B(G146), .C1(KEYINPUT16), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n303), .A2(new_n211), .ZN(new_n308));
  XOR2_X1   g122(.A(KEYINPUT24), .B(G110), .Z(new_n309));
  INV_X1    g123(.A(G128), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(G119), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n188), .A2(G128), .ZN(new_n312));
  OR3_X1    g126(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT72), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT72), .B1(new_n311), .B2(new_n312), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n309), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT23), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n188), .B2(G128), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n310), .A2(KEYINPUT23), .A3(G119), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n317), .B(new_n318), .C1(G119), .C2(new_n310), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(G110), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n307), .B(new_n308), .C1(new_n315), .C2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n304), .B1(KEYINPUT16), .B2(new_n306), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(G146), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n313), .A2(new_n314), .A3(new_n309), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n319), .A2(KEYINPUT73), .A3(G110), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT73), .B1(new_n319), .B2(G110), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n321), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n246), .A2(G221), .A3(G234), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(KEYINPUT22), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n330), .B(G137), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT74), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n328), .A2(new_n334), .ZN(new_n335));
  OAI211_X1 g149(.A(KEYINPUT74), .B(new_n321), .C1(new_n323), .C2(new_n327), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n331), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n333), .B1(new_n337), .B2(KEYINPUT75), .ZN(new_n338));
  OR2_X1    g152(.A1(new_n333), .A2(KEYINPUT75), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI22_X1  g154(.A1(new_n340), .A2(new_n295), .B1(KEYINPUT76), .B2(KEYINPUT25), .ZN(new_n341));
  INV_X1    g155(.A(G234), .ZN(new_n342));
  OAI21_X1  g156(.A(G217), .B1(new_n295), .B2(new_n342), .ZN(new_n343));
  XOR2_X1   g157(.A(new_n343), .B(KEYINPUT71), .Z(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n338), .A2(new_n296), .A3(new_n339), .A4(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n341), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n345), .A2(G902), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n338), .A2(new_n349), .A3(new_n339), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n302), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(G110), .B(G140), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n246), .A2(G227), .ZN(new_n354));
  XOR2_X1   g168(.A(new_n353), .B(new_n354), .Z(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n357));
  AND2_X1   g171(.A1(KEYINPUT77), .A2(G107), .ZN(new_n358));
  NOR2_X1   g172(.A1(KEYINPUT77), .A2(G107), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n357), .B(G104), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G101), .ZN(new_n361));
  INV_X1    g175(.A(G107), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(G104), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(G104), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT3), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n360), .A2(new_n361), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT79), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n363), .B1(KEYINPUT3), .B2(new_n365), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n370), .A2(KEYINPUT79), .A3(new_n360), .A4(new_n361), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  OR2_X1    g186(.A1(KEYINPUT77), .A2(G107), .ZN(new_n373));
  INV_X1    g187(.A(G104), .ZN(new_n374));
  NAND2_X1  g188(.A1(KEYINPUT77), .A2(G107), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT81), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT81), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n373), .A2(new_n378), .A3(new_n374), .A4(new_n375), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n365), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G101), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n372), .A2(KEYINPUT82), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT82), .B1(new_n372), .B2(new_n381), .ZN(new_n383));
  OAI211_X1 g197(.A(KEYINPUT10), .B(new_n232), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n237), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n369), .A2(new_n371), .B1(new_n380), .B2(G101), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n232), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT10), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n370), .A2(new_n360), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G101), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT78), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n361), .B1(new_n370), .B2(new_n360), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT78), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n372), .A2(new_n392), .A3(new_n396), .ZN(new_n397));
  AND4_X1   g211(.A1(KEYINPUT80), .A2(new_n390), .A3(new_n393), .A4(G101), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT80), .B1(new_n394), .B2(new_n393), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n397), .A2(new_n400), .A3(new_n236), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n384), .A2(new_n385), .A3(new_n389), .A4(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n401), .A2(new_n389), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n385), .B1(new_n404), .B2(new_n384), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n356), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n372), .A2(new_n381), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT84), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n408), .A3(new_n264), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT84), .B1(new_n386), .B2(new_n232), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(new_n387), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(KEYINPUT83), .A3(new_n237), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT12), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT12), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n411), .A2(KEYINPUT83), .A3(new_n414), .A4(new_n237), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n413), .A2(new_n402), .A3(new_n415), .A4(new_n355), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n295), .B1(new_n406), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G469), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n413), .A2(new_n402), .A3(new_n415), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n356), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n402), .A2(new_n355), .ZN(new_n422));
  OR2_X1    g236(.A1(new_n422), .A2(new_n405), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(G469), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G902), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n418), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n419), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  XOR2_X1   g242(.A(KEYINPUT9), .B(G234), .Z(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n425), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n430), .A2(G221), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(G113), .B(G122), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(new_n374), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n245), .A2(new_n246), .A3(G214), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(new_n213), .ZN(new_n437));
  NAND2_X1  g251(.A1(KEYINPUT18), .A2(G131), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n303), .B(G146), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT88), .ZN(new_n441));
  OR2_X1    g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n441), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n439), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n437), .A2(G131), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n436), .B(G143), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n203), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n303), .A2(new_n449), .A3(KEYINPUT19), .ZN(new_n450));
  XOR2_X1   g264(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n451));
  OAI21_X1  g265(.A(new_n450), .B1(new_n303), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n211), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n448), .A2(new_n307), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n435), .B1(new_n444), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n437), .A2(KEYINPUT17), .A3(G131), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n323), .B(new_n457), .C1(KEYINPUT17), .C2(new_n448), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n435), .A3(new_n444), .ZN(new_n459));
  AOI21_X1  g273(.A(G475), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT20), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(new_n425), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n461), .B1(new_n460), .B2(new_n425), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n462), .B1(new_n463), .B2(KEYINPUT90), .ZN(new_n464));
  INV_X1    g278(.A(G475), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n458), .A2(new_n435), .A3(new_n444), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n465), .B(new_n425), .C1(new_n466), .C2(new_n455), .ZN(new_n467));
  OR3_X1    g281(.A1(new_n467), .A2(KEYINPUT90), .A3(KEYINPUT20), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n435), .B1(new_n458), .B2(new_n444), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n425), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n464), .A2(new_n468), .B1(G475), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G952), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(G953), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n473), .B1(new_n342), .B2(new_n245), .ZN(new_n474));
  AOI211_X1 g288(.A(new_n246), .B(new_n296), .C1(G234), .C2(G237), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  XOR2_X1   g290(.A(KEYINPUT21), .B(G898), .Z(new_n477));
  OAI21_X1  g291(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(KEYINPUT15), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n191), .A2(G122), .ZN(new_n482));
  INV_X1    g296(.A(G122), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G116), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n373), .A2(new_n375), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n213), .A2(G128), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n310), .A2(G143), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(new_n199), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n482), .A2(KEYINPUT14), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT92), .ZN(new_n493));
  OR2_X1    g307(.A1(new_n482), .A2(KEYINPUT14), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT92), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n482), .A2(new_n495), .A3(KEYINPUT14), .ZN(new_n496));
  AND4_X1   g310(.A1(new_n484), .A2(new_n493), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n487), .B(new_n491), .C1(new_n497), .C2(new_n362), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n485), .B(new_n486), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT13), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n488), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n489), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n488), .A2(new_n500), .ZN(new_n503));
  OAI21_X1  g317(.A(G134), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n490), .A2(new_n199), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT91), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n490), .A2(KEYINPUT91), .A3(new_n199), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n499), .A2(new_n504), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n498), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n429), .A2(G217), .A3(new_n246), .ZN(new_n511));
  XOR2_X1   g325(.A(new_n511), .B(KEYINPUT93), .Z(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n512), .A2(new_n498), .A3(new_n509), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n296), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT94), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT94), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n481), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n481), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n471), .A2(new_n478), .A3(new_n524), .ZN(new_n525));
  XOR2_X1   g339(.A(G110), .B(G122), .Z(new_n526));
  NAND3_X1  g340(.A1(new_n193), .A2(KEYINPUT5), .A3(new_n194), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n527), .B(G113), .C1(KEYINPUT5), .C2(new_n194), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n196), .A2(new_n193), .A3(new_n194), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT82), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n407), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n386), .A2(KEYINPUT82), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n397), .A2(new_n400), .A3(new_n197), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n526), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT85), .ZN(new_n537));
  INV_X1    g351(.A(new_n530), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n538), .B1(new_n382), .B2(new_n383), .ZN(new_n539));
  INV_X1    g353(.A(new_n526), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n397), .A2(new_n400), .A3(new_n197), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n541), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT85), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n544), .A3(new_n526), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n537), .A2(KEYINPUT6), .A3(new_n542), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n224), .A2(G125), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n547), .B1(new_n232), .B2(G125), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n246), .A2(G224), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n548), .B(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT6), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n552), .B(new_n526), .C1(new_n534), .C2(new_n535), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT86), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n543), .A2(KEYINPUT86), .A3(new_n552), .A4(new_n526), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n546), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT7), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n548), .B1(new_n559), .B2(new_n550), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT87), .ZN(new_n561));
  XOR2_X1   g375(.A(new_n526), .B(KEYINPUT8), .Z(new_n562));
  XNOR2_X1  g376(.A(new_n407), .B(new_n530), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n548), .A2(new_n550), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n564), .B(new_n542), .C1(new_n559), .C2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n558), .A2(new_n425), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(G210), .B1(G237), .B2(G902), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n558), .A2(new_n425), .A3(new_n568), .A4(new_n566), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(G214), .B1(G237), .B2(G902), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n433), .A2(new_n525), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n352), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g389(.A(KEYINPUT95), .B(G101), .Z(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(G3));
  INV_X1    g391(.A(KEYINPUT96), .ZN(new_n578));
  INV_X1    g392(.A(G472), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n295), .B1(new_n289), .B2(new_n278), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n351), .B(new_n282), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n428), .A2(new_n432), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n578), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n289), .A2(new_n278), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n296), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n290), .B1(new_n585), .B2(G472), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n586), .A2(KEYINPUT96), .A3(new_n351), .A4(new_n433), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n573), .ZN(new_n589));
  AND4_X1   g403(.A1(new_n425), .A2(new_n558), .A3(new_n568), .A4(new_n566), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n589), .B1(new_n590), .B2(KEYINPUT97), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n517), .A2(new_n479), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n514), .A2(new_n515), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT33), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n514), .A2(KEYINPUT33), .A3(new_n515), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n295), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n592), .B1(new_n597), .B2(new_n479), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT98), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT98), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n592), .B(new_n600), .C1(new_n597), .C2(new_n479), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n471), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT97), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n570), .A2(new_n604), .A3(new_n571), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n591), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n588), .A2(new_n478), .A3(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT34), .B(G104), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G6));
  NAND2_X1  g423(.A1(new_n470), .A2(G475), .ZN(new_n610));
  INV_X1    g424(.A(new_n462), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n610), .B1(new_n611), .B2(new_n463), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n524), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n591), .A2(new_n605), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n588), .A2(new_n478), .A3(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT35), .B(G107), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G9));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n335), .A2(new_n336), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n332), .A2(KEYINPUT36), .ZN(new_n621));
  OR2_X1    g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n619), .B1(new_n624), .B2(new_n349), .ZN(new_n625));
  INV_X1    g439(.A(new_n349), .ZN(new_n626));
  AOI211_X1 g440(.A(KEYINPUT99), .B(new_n626), .C1(new_n622), .C2(new_n623), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n348), .A2(new_n618), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n618), .B1(new_n348), .B2(new_n628), .ZN(new_n630));
  OR2_X1    g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n586), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n574), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT37), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G110), .ZN(G12));
  NOR2_X1   g449(.A1(new_n629), .A2(new_n630), .ZN(new_n636));
  AOI21_X1  g450(.A(KEYINPUT32), .B1(new_n584), .B2(new_n187), .ZN(new_n637));
  AOI211_X1 g451(.A(new_n283), .B(new_n285), .C1(new_n289), .C2(new_n278), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n636), .B1(new_n639), .B2(new_n301), .ZN(new_n640));
  INV_X1    g454(.A(new_n474), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT101), .B(G900), .Z(new_n642));
  AOI21_X1  g456(.A(new_n641), .B1(new_n475), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n582), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n614), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G128), .ZN(G30));
  XOR2_X1   g461(.A(new_n643), .B(KEYINPUT39), .Z(new_n648));
  NAND2_X1  g462(.A1(new_n433), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(KEYINPUT40), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n348), .A2(new_n628), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n650), .A2(new_n589), .A3(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT38), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n572), .B(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n471), .A2(new_n524), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n297), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n262), .B1(new_n658), .B2(new_n242), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT102), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n661), .A2(new_n251), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n579), .B1(new_n663), .B2(new_n425), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n639), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n649), .A2(KEYINPUT40), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n652), .A2(new_n657), .A3(new_n666), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G143), .ZN(G45));
  NAND2_X1  g483(.A1(new_n645), .A2(new_n606), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G146), .ZN(G48));
  INV_X1    g485(.A(KEYINPUT103), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n418), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n417), .A2(new_n674), .ZN(new_n675));
  AOI211_X1 g489(.A(new_n295), .B(new_n673), .C1(new_n406), .C2(new_n416), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n675), .A2(new_n676), .A3(new_n431), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n406), .A2(new_n416), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n296), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n673), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n417), .A2(new_n674), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n432), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT104), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n302), .A3(new_n351), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n591), .A2(new_n605), .A3(new_n478), .A4(new_n603), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT41), .B(G113), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  NAND2_X1  g505(.A1(new_n614), .A2(new_n478), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n687), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n191), .ZN(G18));
  AND3_X1   g508(.A1(new_n591), .A2(new_n605), .A3(new_n677), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n695), .A2(new_n302), .A3(new_n525), .A4(new_n631), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  AOI22_X1  g511(.A1(new_n298), .A2(new_n262), .B1(KEYINPUT31), .B2(new_n251), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n285), .B1(new_n698), .B2(new_n277), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n585), .B2(G472), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n677), .A2(new_n678), .ZN(new_n701));
  NOR4_X1   g515(.A1(new_n675), .A2(new_n676), .A3(KEYINPUT104), .A4(new_n431), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n700), .B(new_n351), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n591), .A2(new_n605), .A3(new_n478), .A4(new_n655), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n483), .ZN(G24));
  NAND2_X1  g520(.A1(new_n585), .A2(G472), .ZN(new_n707));
  INV_X1    g521(.A(new_n699), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n471), .A2(new_n602), .A3(new_n643), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n707), .A2(new_n651), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n591), .A2(new_n605), .A3(new_n677), .ZN(new_n711));
  OAI21_X1  g525(.A(KEYINPUT105), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n651), .B(new_n708), .C1(new_n580), .C2(new_n579), .ZN(new_n713));
  INV_X1    g527(.A(new_n709), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n695), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(new_n718), .B(KEYINPUT106), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  NAND2_X1  g534(.A1(new_n424), .A2(KEYINPUT107), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n421), .A2(new_n423), .A3(new_n722), .A4(G469), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n721), .A2(new_n419), .A3(new_n427), .A4(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n431), .A2(new_n589), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n724), .A2(new_n570), .A3(new_n571), .A4(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT108), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n570), .A2(new_n571), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT108), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(new_n729), .A3(new_n725), .A4(new_n724), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n351), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n732), .B1(new_n639), .B2(new_n301), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n731), .A2(new_n733), .A3(new_n709), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT42), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n731), .A2(KEYINPUT42), .A3(new_n733), .A4(new_n709), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT109), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n203), .ZN(G33));
  INV_X1    g554(.A(new_n643), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n731), .A2(new_n733), .A3(new_n613), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  NAND2_X1  g557(.A1(new_n421), .A2(new_n423), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n421), .A2(KEYINPUT45), .A3(new_n423), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(G469), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n427), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT46), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n748), .A2(KEYINPUT46), .A3(new_n427), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n419), .A3(new_n752), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n753), .A2(new_n432), .A3(new_n648), .ZN(new_n754));
  INV_X1    g568(.A(new_n586), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n464), .A2(new_n468), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(new_n610), .A3(new_n599), .A4(new_n601), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n758), .A3(KEYINPUT43), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n755), .A2(new_n651), .A3(new_n759), .A4(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n572), .A2(new_n589), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n767), .B1(new_n766), .B2(new_n768), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n754), .B(new_n765), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  INV_X1    g586(.A(new_n768), .ZN(new_n773));
  NOR4_X1   g587(.A1(new_n773), .A2(new_n302), .A3(new_n351), .A4(new_n714), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n753), .A2(new_n432), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT112), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n753), .A2(new_n779), .A3(new_n432), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n778), .A2(KEYINPUT47), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n753), .A2(new_n779), .A3(new_n432), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n779), .B1(new_n753), .B2(new_n432), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n776), .A2(new_n781), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT114), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  OAI21_X1  g602(.A(new_n696), .B1(new_n692), .B2(new_n687), .ZN(new_n789));
  OAI22_X1  g603(.A1(new_n687), .A2(new_n688), .B1(new_n703), .B2(new_n704), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n574), .B1(new_n352), .B2(new_n632), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n524), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT116), .B1(new_n521), .B2(new_n523), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n795), .A2(new_n756), .A3(new_n610), .A4(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n797), .B1(new_n471), .B2(new_n602), .ZN(new_n798));
  AND4_X1   g612(.A1(new_n478), .A2(new_n798), .A3(new_n572), .A4(new_n573), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n583), .A2(new_n587), .A3(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n612), .B1(new_n795), .B2(new_n796), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n645), .A2(new_n768), .A3(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n791), .A2(new_n793), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n731), .A2(new_n715), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n742), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n738), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n640), .B(new_n644), .C1(new_n606), .C2(new_n614), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n591), .A2(new_n605), .A3(new_n655), .ZN(new_n811));
  INV_X1    g625(.A(new_n724), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n812), .A2(new_n651), .A3(new_n643), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n666), .A2(new_n811), .A3(new_n813), .A4(new_n432), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n718), .A2(new_n810), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT52), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n718), .A2(new_n810), .A3(new_n814), .A4(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n817), .B1(new_n816), .B2(new_n819), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n808), .B(new_n809), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NOR4_X1   g636(.A1(new_n789), .A2(new_n790), .A3(new_n800), .A4(new_n792), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n742), .A2(new_n805), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n736), .B2(new_n737), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n823), .A2(new_n825), .A3(new_n803), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n816), .A2(new_n819), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT53), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n822), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT118), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n809), .B1(new_n826), .B2(new_n827), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n808), .B1(new_n820), .B2(new_n821), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n833), .B1(new_n834), .B2(new_n809), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT54), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT54), .B1(new_n822), .B2(new_n828), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n785), .A2(new_n781), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n675), .A2(new_n676), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n431), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT120), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n700), .A2(new_n351), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n762), .A2(new_n641), .A3(new_n759), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n768), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  AOI22_X1  g663(.A1(new_n785), .A2(new_n781), .B1(new_n431), .B2(new_n841), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n844), .A2(new_n849), .A3(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n654), .A2(new_n589), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(KEYINPUT50), .A3(new_n677), .A4(new_n847), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT50), .ZN(new_n856));
  INV_X1    g670(.A(new_n759), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT43), .B1(new_n757), .B2(new_n758), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n857), .A2(new_n858), .A3(new_n474), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n351), .A3(new_n677), .A4(new_n700), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n654), .A2(new_n589), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n856), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n855), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n846), .A2(new_n773), .A3(new_n684), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n651), .A3(new_n700), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n666), .A2(new_n474), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n773), .A2(new_n732), .A3(new_n684), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n866), .A2(new_n867), .A3(new_n471), .A4(new_n602), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n863), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n869), .A2(KEYINPUT119), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT51), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT119), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n853), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n866), .A2(new_n867), .A3(new_n603), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n847), .A2(new_n695), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n874), .A2(new_n473), .A3(new_n875), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n863), .A2(new_n865), .A3(new_n868), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n877), .B1(new_n848), .B2(new_n850), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n876), .B1(new_n878), .B2(new_n871), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n864), .A2(new_n733), .ZN(new_n880));
  XOR2_X1   g694(.A(KEYINPUT121), .B(KEYINPUT48), .Z(new_n881));
  XNOR2_X1  g695(.A(new_n880), .B(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n873), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n832), .A2(new_n836), .A3(new_n839), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT122), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n838), .B1(new_n829), .B2(new_n830), .ZN(new_n886));
  AOI211_X1 g700(.A(KEYINPUT118), .B(KEYINPUT54), .C1(new_n822), .C2(new_n828), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n888), .A2(new_n889), .A3(new_n836), .A4(new_n883), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n472), .A2(new_n246), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n885), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n351), .A2(new_n725), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT115), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n894), .A2(new_n757), .ZN(new_n895));
  INV_X1    g709(.A(new_n666), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n841), .B(KEYINPUT49), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n895), .A2(new_n654), .A3(new_n896), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n892), .A2(new_n898), .ZN(G75));
  NOR2_X1   g713(.A1(new_n829), .A2(new_n296), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT56), .B1(new_n900), .B2(new_n569), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n546), .A2(new_n557), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n551), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT55), .Z(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n901), .A2(new_n905), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n246), .A2(G952), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT123), .Z(new_n909));
  NOR3_X1   g723(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(G51));
  XNOR2_X1  g724(.A(new_n426), .B(KEYINPUT57), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n829), .A2(new_n830), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n911), .B1(new_n912), .B2(new_n837), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n680), .ZN(new_n914));
  OR3_X1    g728(.A1(new_n829), .A2(new_n296), .A3(new_n748), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n908), .B1(new_n914), .B2(new_n915), .ZN(G54));
  NAND3_X1  g730(.A1(new_n900), .A2(KEYINPUT58), .A3(G475), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n917), .A2(new_n459), .A3(new_n456), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n917), .B1(new_n459), .B2(new_n456), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n908), .ZN(G60));
  NAND2_X1  g734(.A1(new_n595), .A2(new_n596), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT124), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n832), .A2(new_n836), .A3(new_n839), .ZN(new_n923));
  NAND2_X1  g737(.A1(G478), .A2(G902), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT59), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n922), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n925), .B(new_n922), .C1(new_n912), .C2(new_n837), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n926), .A2(new_n909), .A3(new_n928), .ZN(G63));
  NAND2_X1  g743(.A1(G217), .A2(G902), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT60), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n930), .B(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n822), .A2(new_n828), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n909), .B1(new_n933), .B2(new_n340), .ZN(new_n934));
  INV_X1    g748(.A(new_n624), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n934), .B1(new_n935), .B2(new_n933), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g751(.A(new_n246), .B1(new_n477), .B2(G224), .ZN(new_n938));
  INV_X1    g752(.A(new_n823), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n938), .B1(new_n939), .B2(new_n246), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n902), .B1(G898), .B2(new_n246), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n940), .B(new_n941), .Z(G69));
  XNOR2_X1  g756(.A(new_n270), .B(new_n452), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n718), .A2(new_n810), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n771), .A2(new_n786), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n754), .A2(new_n733), .A3(new_n811), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n738), .A2(new_n742), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n246), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n246), .A2(G900), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n948), .A2(KEYINPUT126), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT126), .B1(new_n948), .B2(new_n950), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n943), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n944), .A2(new_n668), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT62), .Z(new_n955));
  AND2_X1   g769(.A1(new_n771), .A2(new_n786), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT125), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n649), .B1(new_n957), .B2(new_n798), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n798), .A2(new_n957), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n958), .A2(new_n733), .A3(new_n768), .A4(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n955), .A2(new_n956), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n943), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n961), .A2(new_n246), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n953), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(G227), .A2(G900), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(G953), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n964), .B(new_n966), .ZN(G72));
  XNOR2_X1  g781(.A(new_n271), .B(KEYINPUT127), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n945), .A2(new_n939), .A3(new_n947), .ZN(new_n969));
  NAND2_X1  g783(.A1(G472), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT63), .Z(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n262), .B(new_n968), .C1(new_n969), .C2(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n971), .B1(new_n961), .B2(new_n939), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n250), .ZN(new_n975));
  OAI221_X1 g789(.A(new_n973), .B1(G952), .B2(new_n246), .C1(new_n975), .C2(new_n968), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n271), .B(new_n250), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n835), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n976), .B1(new_n971), .B2(new_n978), .ZN(G57));
endmodule


