

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X2 U547 ( .A(n712), .ZN(n595) );
  XNOR2_X1 U548 ( .A(n644), .B(n643), .ZN(n646) );
  NAND2_X1 U549 ( .A1(G8), .A2(n653), .ZN(n693) );
  AND2_X1 U550 ( .A1(G137), .A2(n861), .ZN(n586) );
  XOR2_X1 U551 ( .A(KEYINPUT31), .B(n649), .Z(n513) );
  XOR2_X1 U552 ( .A(n738), .B(KEYINPUT97), .Z(n514) );
  AND2_X1 U553 ( .A1(n726), .A2(n732), .ZN(n515) );
  OR2_X1 U554 ( .A1(n695), .A2(n694), .ZN(n516) );
  AND2_X1 U555 ( .A1(n646), .A2(n645), .ZN(n517) );
  XNOR2_X1 U556 ( .A(KEYINPUT30), .B(KEYINPUT93), .ZN(n643) );
  INV_X1 U557 ( .A(G168), .ZN(n645) );
  NOR2_X1 U558 ( .A1(G1966), .A2(n693), .ZN(n667) );
  AND2_X1 U559 ( .A1(n660), .A2(n659), .ZN(n662) );
  XNOR2_X1 U560 ( .A(n662), .B(n661), .ZN(n683) );
  OR2_X1 U561 ( .A1(n742), .A2(n594), .ZN(n712) );
  NOR2_X1 U562 ( .A1(G2105), .A2(G2104), .ZN(n575) );
  NOR2_X1 U563 ( .A1(G651), .A2(n554), .ZN(n770) );
  NOR2_X1 U564 ( .A1(G2105), .A2(n578), .ZN(n862) );
  INV_X1 U565 ( .A(KEYINPUT23), .ZN(n587) );
  NOR2_X1 U566 ( .A1(G651), .A2(G543), .ZN(n775) );
  XNOR2_X1 U567 ( .A(n588), .B(n587), .ZN(n589) );
  NAND2_X1 U568 ( .A1(n590), .A2(n589), .ZN(n742) );
  INV_X1 U569 ( .A(G651), .ZN(n521) );
  NOR2_X1 U570 ( .A1(G543), .A2(n521), .ZN(n518) );
  XOR2_X1 U571 ( .A(KEYINPUT1), .B(n518), .Z(n769) );
  NAND2_X1 U572 ( .A1(G65), .A2(n769), .ZN(n520) );
  NAND2_X1 U573 ( .A1(G91), .A2(n775), .ZN(n519) );
  NAND2_X1 U574 ( .A1(n520), .A2(n519), .ZN(n525) );
  XOR2_X1 U575 ( .A(G543), .B(KEYINPUT0), .Z(n554) );
  NOR2_X1 U576 ( .A1(n554), .A2(n521), .ZN(n774) );
  NAND2_X1 U577 ( .A1(G78), .A2(n774), .ZN(n523) );
  NAND2_X1 U578 ( .A1(G53), .A2(n770), .ZN(n522) );
  NAND2_X1 U579 ( .A1(n523), .A2(n522), .ZN(n524) );
  OR2_X1 U580 ( .A1(n525), .A2(n524), .ZN(G299) );
  NAND2_X1 U581 ( .A1(G63), .A2(n769), .ZN(n527) );
  NAND2_X1 U582 ( .A1(G51), .A2(n770), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U584 ( .A(KEYINPUT6), .B(n528), .ZN(n537) );
  NAND2_X1 U585 ( .A1(G76), .A2(n774), .ZN(n533) );
  XOR2_X1 U586 ( .A(KEYINPUT4), .B(KEYINPUT68), .Z(n530) );
  NAND2_X1 U587 ( .A1(G89), .A2(n775), .ZN(n529) );
  XNOR2_X1 U588 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U589 ( .A(KEYINPUT67), .B(n531), .ZN(n532) );
  NAND2_X1 U590 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U591 ( .A(n534), .B(KEYINPUT5), .ZN(n535) );
  XNOR2_X1 U592 ( .A(n535), .B(KEYINPUT69), .ZN(n536) );
  NOR2_X1 U593 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U594 ( .A(KEYINPUT7), .B(n538), .Z(G168) );
  NAND2_X1 U595 ( .A1(G64), .A2(n769), .ZN(n540) );
  NAND2_X1 U596 ( .A1(G52), .A2(n770), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n546) );
  NAND2_X1 U598 ( .A1(n775), .A2(G90), .ZN(n541) );
  XOR2_X1 U599 ( .A(KEYINPUT65), .B(n541), .Z(n543) );
  NAND2_X1 U600 ( .A1(n774), .A2(G77), .ZN(n542) );
  NAND2_X1 U601 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U602 ( .A(KEYINPUT9), .B(n544), .Z(n545) );
  NOR2_X1 U603 ( .A1(n546), .A2(n545), .ZN(G171) );
  XOR2_X1 U604 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U605 ( .A1(G88), .A2(n775), .ZN(n547) );
  XNOR2_X1 U606 ( .A(n547), .B(KEYINPUT78), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n774), .A2(G75), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n549), .A2(n548), .ZN(n553) );
  NAND2_X1 U609 ( .A1(G62), .A2(n769), .ZN(n551) );
  NAND2_X1 U610 ( .A1(G50), .A2(n770), .ZN(n550) );
  NAND2_X1 U611 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U612 ( .A1(n553), .A2(n552), .ZN(G166) );
  INV_X1 U613 ( .A(G166), .ZN(G303) );
  NAND2_X1 U614 ( .A1(G74), .A2(G651), .ZN(n559) );
  NAND2_X1 U615 ( .A1(G49), .A2(n770), .ZN(n556) );
  NAND2_X1 U616 ( .A1(G87), .A2(n554), .ZN(n555) );
  NAND2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U618 ( .A1(n769), .A2(n557), .ZN(n558) );
  NAND2_X1 U619 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U620 ( .A(n560), .B(KEYINPUT76), .ZN(G288) );
  NAND2_X1 U621 ( .A1(G61), .A2(n769), .ZN(n562) );
  NAND2_X1 U622 ( .A1(G48), .A2(n770), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n566) );
  XOR2_X1 U624 ( .A(KEYINPUT2), .B(KEYINPUT77), .Z(n564) );
  NAND2_X1 U625 ( .A1(n774), .A2(G73), .ZN(n563) );
  XOR2_X1 U626 ( .A(n564), .B(n563), .Z(n565) );
  NOR2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U628 ( .A1(n775), .A2(G86), .ZN(n567) );
  NAND2_X1 U629 ( .A1(n568), .A2(n567), .ZN(G305) );
  NAND2_X1 U630 ( .A1(G60), .A2(n769), .ZN(n570) );
  NAND2_X1 U631 ( .A1(G85), .A2(n775), .ZN(n569) );
  NAND2_X1 U632 ( .A1(n570), .A2(n569), .ZN(n574) );
  NAND2_X1 U633 ( .A1(G72), .A2(n774), .ZN(n572) );
  NAND2_X1 U634 ( .A1(G47), .A2(n770), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n572), .A2(n571), .ZN(n573) );
  OR2_X1 U636 ( .A1(n574), .A2(n573), .ZN(G290) );
  XOR2_X2 U637 ( .A(KEYINPUT17), .B(n575), .Z(n861) );
  NAND2_X1 U638 ( .A1(G138), .A2(n861), .ZN(n577) );
  INV_X1 U639 ( .A(G2104), .ZN(n578) );
  NAND2_X1 U640 ( .A1(G102), .A2(n862), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n583) );
  AND2_X1 U642 ( .A1(n578), .A2(G2105), .ZN(n865) );
  NAND2_X1 U643 ( .A1(G126), .A2(n865), .ZN(n580) );
  AND2_X1 U644 ( .A1(G2105), .A2(G2104), .ZN(n866) );
  NAND2_X1 U645 ( .A1(G114), .A2(n866), .ZN(n579) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U647 ( .A(KEYINPUT83), .B(n581), .Z(n582) );
  NOR2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(KEYINPUT84), .B(n584), .ZN(n741) );
  NOR2_X1 U650 ( .A1(G1384), .A2(n741), .ZN(n713) );
  INV_X1 U651 ( .A(KEYINPUT64), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(n590) );
  NAND2_X1 U653 ( .A1(G101), .A2(n862), .ZN(n588) );
  INV_X1 U654 ( .A(G40), .ZN(n593) );
  NAND2_X1 U655 ( .A1(G125), .A2(n865), .ZN(n592) );
  NAND2_X1 U656 ( .A1(G113), .A2(n866), .ZN(n591) );
  NAND2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n743) );
  OR2_X1 U658 ( .A1(n593), .A2(n743), .ZN(n594) );
  NAND2_X2 U659 ( .A1(n713), .A2(n595), .ZN(n653) );
  NAND2_X1 U660 ( .A1(G56), .A2(n769), .ZN(n596) );
  XOR2_X1 U661 ( .A(KEYINPUT14), .B(n596), .Z(n602) );
  NAND2_X1 U662 ( .A1(n775), .A2(G81), .ZN(n597) );
  XNOR2_X1 U663 ( .A(n597), .B(KEYINPUT12), .ZN(n599) );
  NAND2_X1 U664 ( .A1(G68), .A2(n774), .ZN(n598) );
  NAND2_X1 U665 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U666 ( .A(KEYINPUT13), .B(n600), .Z(n601) );
  NOR2_X1 U667 ( .A1(n602), .A2(n601), .ZN(n604) );
  NAND2_X1 U668 ( .A1(n770), .A2(G43), .ZN(n603) );
  NAND2_X1 U669 ( .A1(n604), .A2(n603), .ZN(n942) );
  INV_X1 U670 ( .A(G1996), .ZN(n907) );
  NOR2_X1 U671 ( .A1(n653), .A2(n907), .ZN(n605) );
  XOR2_X1 U672 ( .A(n605), .B(KEYINPUT26), .Z(n607) );
  NAND2_X1 U673 ( .A1(n653), .A2(G1341), .ZN(n606) );
  NAND2_X1 U674 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U675 ( .A1(n942), .A2(n608), .ZN(n620) );
  NAND2_X1 U676 ( .A1(n770), .A2(G54), .ZN(n615) );
  NAND2_X1 U677 ( .A1(G79), .A2(n774), .ZN(n610) );
  NAND2_X1 U678 ( .A1(G66), .A2(n769), .ZN(n609) );
  NAND2_X1 U679 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U680 ( .A1(n775), .A2(G92), .ZN(n611) );
  XOR2_X1 U681 ( .A(KEYINPUT66), .B(n611), .Z(n612) );
  NOR2_X1 U682 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U683 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U684 ( .A(KEYINPUT15), .B(n616), .Z(n753) );
  NAND2_X1 U685 ( .A1(G1348), .A2(n653), .ZN(n618) );
  INV_X2 U686 ( .A(n653), .ZN(n636) );
  NAND2_X1 U687 ( .A1(G2067), .A2(n636), .ZN(n617) );
  NAND2_X1 U688 ( .A1(n618), .A2(n617), .ZN(n621) );
  NOR2_X1 U689 ( .A1(n753), .A2(n621), .ZN(n619) );
  NOR2_X1 U690 ( .A1(n620), .A2(n619), .ZN(n623) );
  AND2_X1 U691 ( .A1(n753), .A2(n621), .ZN(n622) );
  NOR2_X1 U692 ( .A1(n623), .A2(n622), .ZN(n630) );
  NAND2_X1 U693 ( .A1(n636), .A2(G2072), .ZN(n624) );
  XOR2_X1 U694 ( .A(n624), .B(KEYINPUT27), .Z(n627) );
  XOR2_X1 U695 ( .A(KEYINPUT90), .B(G1956), .Z(n966) );
  NOR2_X1 U696 ( .A1(n636), .A2(n966), .ZN(n625) );
  XNOR2_X1 U697 ( .A(KEYINPUT91), .B(n625), .ZN(n626) );
  NAND2_X1 U698 ( .A1(n627), .A2(n626), .ZN(n631) );
  NOR2_X1 U699 ( .A1(G299), .A2(n631), .ZN(n628) );
  XNOR2_X1 U700 ( .A(n628), .B(KEYINPUT92), .ZN(n629) );
  NOR2_X1 U701 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U702 ( .A1(n631), .A2(G299), .ZN(n632) );
  XOR2_X1 U703 ( .A(KEYINPUT28), .B(n632), .Z(n633) );
  NOR2_X2 U704 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U705 ( .A(KEYINPUT29), .B(n635), .ZN(n641) );
  INV_X1 U706 ( .A(G1961), .ZN(n962) );
  NAND2_X1 U707 ( .A1(n653), .A2(n962), .ZN(n638) );
  XNOR2_X1 U708 ( .A(KEYINPUT25), .B(G2078), .ZN(n914) );
  NAND2_X1 U709 ( .A1(n636), .A2(n914), .ZN(n637) );
  NAND2_X1 U710 ( .A1(n638), .A2(n637), .ZN(n647) );
  AND2_X1 U711 ( .A1(n647), .A2(G171), .ZN(n639) );
  XNOR2_X1 U712 ( .A(KEYINPUT89), .B(n639), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n641), .A2(n640), .ZN(n650) );
  NOR2_X1 U714 ( .A1(G2084), .A2(n653), .ZN(n663) );
  NOR2_X1 U715 ( .A1(n667), .A2(n663), .ZN(n642) );
  NAND2_X1 U716 ( .A1(G8), .A2(n642), .ZN(n644) );
  NOR2_X1 U717 ( .A1(G171), .A2(n647), .ZN(n648) );
  NOR2_X1 U718 ( .A1(n517), .A2(n648), .ZN(n649) );
  NAND2_X1 U719 ( .A1(n650), .A2(n513), .ZN(n665) );
  AND2_X1 U720 ( .A1(G286), .A2(G8), .ZN(n651) );
  NAND2_X1 U721 ( .A1(n665), .A2(n651), .ZN(n660) );
  INV_X1 U722 ( .A(G8), .ZN(n658) );
  NOR2_X1 U723 ( .A1(G1971), .A2(n693), .ZN(n652) );
  XNOR2_X1 U724 ( .A(n652), .B(KEYINPUT94), .ZN(n655) );
  NOR2_X1 U725 ( .A1(n653), .A2(G2090), .ZN(n654) );
  NOR2_X1 U726 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U727 ( .A1(n656), .A2(G303), .ZN(n657) );
  OR2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U729 ( .A(KEYINPUT95), .B(KEYINPUT32), .Z(n661) );
  NAND2_X1 U730 ( .A1(G8), .A2(n663), .ZN(n664) );
  XNOR2_X1 U731 ( .A(KEYINPUT88), .B(n664), .ZN(n669) );
  INV_X1 U732 ( .A(n665), .ZN(n666) );
  NOR2_X1 U733 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n682) );
  NAND2_X1 U735 ( .A1(G1976), .A2(G288), .ZN(n932) );
  AND2_X1 U736 ( .A1(n682), .A2(n932), .ZN(n670) );
  NAND2_X1 U737 ( .A1(n683), .A2(n670), .ZN(n675) );
  INV_X1 U738 ( .A(n932), .ZN(n673) );
  NOR2_X1 U739 ( .A1(G1976), .A2(G288), .ZN(n930) );
  NOR2_X1 U740 ( .A1(G1971), .A2(G303), .ZN(n671) );
  NOR2_X1 U741 ( .A1(n930), .A2(n671), .ZN(n672) );
  OR2_X1 U742 ( .A1(n673), .A2(n672), .ZN(n674) );
  AND2_X1 U743 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U744 ( .A1(n693), .A2(n676), .ZN(n677) );
  NOR2_X1 U745 ( .A1(KEYINPUT33), .A2(n677), .ZN(n680) );
  NAND2_X1 U746 ( .A1(n930), .A2(KEYINPUT33), .ZN(n678) );
  NOR2_X1 U747 ( .A1(n678), .A2(n693), .ZN(n679) );
  NOR2_X1 U748 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U749 ( .A(G1981), .B(G305), .Z(n947) );
  NAND2_X1 U750 ( .A1(n681), .A2(n947), .ZN(n689) );
  NAND2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n686) );
  NOR2_X1 U752 ( .A1(G2090), .A2(G303), .ZN(n684) );
  NAND2_X1 U753 ( .A1(G8), .A2(n684), .ZN(n685) );
  NAND2_X1 U754 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U755 ( .A1(n687), .A2(n693), .ZN(n688) );
  NAND2_X1 U756 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U757 ( .A(n690), .B(KEYINPUT96), .ZN(n695) );
  NOR2_X1 U758 ( .A1(G1981), .A2(G305), .ZN(n691) );
  XOR2_X1 U759 ( .A(n691), .B(KEYINPUT24), .Z(n692) );
  NOR2_X1 U760 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U761 ( .A1(G119), .A2(n865), .ZN(n697) );
  NAND2_X1 U762 ( .A1(G131), .A2(n861), .ZN(n696) );
  NAND2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n701) );
  NAND2_X1 U764 ( .A1(G107), .A2(n866), .ZN(n699) );
  NAND2_X1 U765 ( .A1(G95), .A2(n862), .ZN(n698) );
  NAND2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n700) );
  OR2_X1 U767 ( .A1(n701), .A2(n700), .ZN(n855) );
  NAND2_X1 U768 ( .A1(G1991), .A2(n855), .ZN(n702) );
  XOR2_X1 U769 ( .A(KEYINPUT87), .B(n702), .Z(n711) );
  NAND2_X1 U770 ( .A1(G129), .A2(n865), .ZN(n704) );
  NAND2_X1 U771 ( .A1(G141), .A2(n861), .ZN(n703) );
  NAND2_X1 U772 ( .A1(n704), .A2(n703), .ZN(n707) );
  NAND2_X1 U773 ( .A1(n862), .A2(G105), .ZN(n705) );
  XOR2_X1 U774 ( .A(KEYINPUT38), .B(n705), .Z(n706) );
  NOR2_X1 U775 ( .A1(n707), .A2(n706), .ZN(n709) );
  NAND2_X1 U776 ( .A1(n866), .A2(G117), .ZN(n708) );
  NAND2_X1 U777 ( .A1(n709), .A2(n708), .ZN(n873) );
  NAND2_X1 U778 ( .A1(G1996), .A2(n873), .ZN(n710) );
  NAND2_X1 U779 ( .A1(n711), .A2(n710), .ZN(n729) );
  INV_X1 U780 ( .A(n729), .ZN(n997) );
  XOR2_X1 U781 ( .A(G1986), .B(G290), .Z(n940) );
  NAND2_X1 U782 ( .A1(n997), .A2(n940), .ZN(n714) );
  NOR2_X1 U783 ( .A1(n713), .A2(n712), .ZN(n737) );
  NAND2_X1 U784 ( .A1(n714), .A2(n737), .ZN(n726) );
  NAND2_X1 U785 ( .A1(G140), .A2(n861), .ZN(n716) );
  NAND2_X1 U786 ( .A1(G104), .A2(n862), .ZN(n715) );
  NAND2_X1 U787 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U788 ( .A(KEYINPUT34), .B(n717), .ZN(n723) );
  NAND2_X1 U789 ( .A1(n865), .A2(G128), .ZN(n718) );
  XOR2_X1 U790 ( .A(KEYINPUT85), .B(n718), .Z(n720) );
  NAND2_X1 U791 ( .A1(n866), .A2(G116), .ZN(n719) );
  NAND2_X1 U792 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U793 ( .A(n721), .B(KEYINPUT35), .Z(n722) );
  NOR2_X1 U794 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U795 ( .A(KEYINPUT36), .B(n724), .Z(n725) );
  XOR2_X1 U796 ( .A(KEYINPUT86), .B(n725), .Z(n878) );
  XNOR2_X1 U797 ( .A(G2067), .B(KEYINPUT37), .ZN(n734) );
  NOR2_X1 U798 ( .A1(n878), .A2(n734), .ZN(n989) );
  NAND2_X1 U799 ( .A1(n989), .A2(n737), .ZN(n732) );
  NAND2_X1 U800 ( .A1(n516), .A2(n515), .ZN(n739) );
  NOR2_X1 U801 ( .A1(G1996), .A2(n873), .ZN(n994) );
  NOR2_X1 U802 ( .A1(G1986), .A2(G290), .ZN(n727) );
  NOR2_X1 U803 ( .A1(G1991), .A2(n855), .ZN(n988) );
  NOR2_X1 U804 ( .A1(n727), .A2(n988), .ZN(n728) );
  NOR2_X1 U805 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U806 ( .A1(n994), .A2(n730), .ZN(n731) );
  XNOR2_X1 U807 ( .A(KEYINPUT39), .B(n731), .ZN(n733) );
  NAND2_X1 U808 ( .A1(n733), .A2(n732), .ZN(n735) );
  NAND2_X1 U809 ( .A1(n878), .A2(n734), .ZN(n1006) );
  NAND2_X1 U810 ( .A1(n735), .A2(n1006), .ZN(n736) );
  NAND2_X1 U811 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U812 ( .A1(n739), .A2(n514), .ZN(n740) );
  XNOR2_X1 U813 ( .A(n740), .B(KEYINPUT40), .ZN(G329) );
  BUF_X1 U814 ( .A(n741), .Z(G164) );
  AND2_X1 U815 ( .A1(G452), .A2(G94), .ZN(G173) );
  NOR2_X1 U816 ( .A1(n743), .A2(n742), .ZN(G160) );
  INV_X1 U817 ( .A(G57), .ZN(G237) );
  INV_X1 U818 ( .A(G132), .ZN(G219) );
  INV_X1 U819 ( .A(G82), .ZN(G220) );
  NAND2_X1 U820 ( .A1(G7), .A2(G661), .ZN(n744) );
  XNOR2_X1 U821 ( .A(n744), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U822 ( .A(G223), .ZN(n812) );
  NAND2_X1 U823 ( .A1(n812), .A2(G567), .ZN(n745) );
  XOR2_X1 U824 ( .A(KEYINPUT11), .B(n745), .Z(G234) );
  INV_X1 U825 ( .A(G860), .ZN(n781) );
  OR2_X1 U826 ( .A1(n942), .A2(n781), .ZN(G153) );
  INV_X1 U827 ( .A(G171), .ZN(G301) );
  NAND2_X1 U828 ( .A1(G868), .A2(G301), .ZN(n747) );
  INV_X1 U829 ( .A(G868), .ZN(n792) );
  NAND2_X1 U830 ( .A1(n753), .A2(n792), .ZN(n746) );
  NAND2_X1 U831 ( .A1(n747), .A2(n746), .ZN(G284) );
  NOR2_X1 U832 ( .A1(G286), .A2(n792), .ZN(n748) );
  XNOR2_X1 U833 ( .A(n748), .B(KEYINPUT70), .ZN(n750) );
  NOR2_X1 U834 ( .A1(G299), .A2(G868), .ZN(n749) );
  NOR2_X1 U835 ( .A1(n750), .A2(n749), .ZN(G297) );
  NAND2_X1 U836 ( .A1(n781), .A2(G559), .ZN(n751) );
  INV_X1 U837 ( .A(n753), .ZN(n939) );
  NAND2_X1 U838 ( .A1(n751), .A2(n939), .ZN(n752) );
  XNOR2_X1 U839 ( .A(n752), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U840 ( .A1(n753), .A2(n792), .ZN(n754) );
  XNOR2_X1 U841 ( .A(n754), .B(KEYINPUT71), .ZN(n755) );
  NOR2_X1 U842 ( .A1(G559), .A2(n755), .ZN(n757) );
  NOR2_X1 U843 ( .A1(G868), .A2(n942), .ZN(n756) );
  NOR2_X1 U844 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U845 ( .A(KEYINPUT72), .B(n758), .ZN(G282) );
  NAND2_X1 U846 ( .A1(G123), .A2(n865), .ZN(n759) );
  XOR2_X1 U847 ( .A(KEYINPUT73), .B(n759), .Z(n760) );
  XNOR2_X1 U848 ( .A(n760), .B(KEYINPUT18), .ZN(n762) );
  NAND2_X1 U849 ( .A1(G111), .A2(n866), .ZN(n761) );
  NAND2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n766) );
  NAND2_X1 U851 ( .A1(G135), .A2(n861), .ZN(n764) );
  NAND2_X1 U852 ( .A1(G99), .A2(n862), .ZN(n763) );
  NAND2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n987) );
  XNOR2_X1 U855 ( .A(G2096), .B(n987), .ZN(n768) );
  INV_X1 U856 ( .A(G2100), .ZN(n767) );
  NAND2_X1 U857 ( .A1(n768), .A2(n767), .ZN(G156) );
  NAND2_X1 U858 ( .A1(G67), .A2(n769), .ZN(n772) );
  NAND2_X1 U859 ( .A1(G55), .A2(n770), .ZN(n771) );
  NAND2_X1 U860 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U861 ( .A(KEYINPUT74), .B(n773), .ZN(n779) );
  NAND2_X1 U862 ( .A1(G80), .A2(n774), .ZN(n777) );
  NAND2_X1 U863 ( .A1(G93), .A2(n775), .ZN(n776) );
  NAND2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n778) );
  OR2_X1 U865 ( .A1(n779), .A2(n778), .ZN(n793) );
  NAND2_X1 U866 ( .A1(G559), .A2(n939), .ZN(n780) );
  XOR2_X1 U867 ( .A(n942), .B(n780), .Z(n790) );
  NAND2_X1 U868 ( .A1(n781), .A2(n790), .ZN(n782) );
  XNOR2_X1 U869 ( .A(n782), .B(KEYINPUT75), .ZN(n783) );
  XOR2_X1 U870 ( .A(n793), .B(n783), .Z(G145) );
  XNOR2_X1 U871 ( .A(G166), .B(KEYINPUT79), .ZN(n784) );
  XNOR2_X1 U872 ( .A(n784), .B(KEYINPUT19), .ZN(n785) );
  XOR2_X1 U873 ( .A(n793), .B(n785), .Z(n787) );
  XNOR2_X1 U874 ( .A(G305), .B(G288), .ZN(n786) );
  XNOR2_X1 U875 ( .A(n787), .B(n786), .ZN(n788) );
  XNOR2_X1 U876 ( .A(n788), .B(G299), .ZN(n789) );
  XNOR2_X1 U877 ( .A(n789), .B(G290), .ZN(n881) );
  XOR2_X1 U878 ( .A(n881), .B(n790), .Z(n791) );
  NOR2_X1 U879 ( .A1(n792), .A2(n791), .ZN(n795) );
  NOR2_X1 U880 ( .A1(G868), .A2(n793), .ZN(n794) );
  NOR2_X1 U881 ( .A1(n795), .A2(n794), .ZN(G295) );
  NAND2_X1 U882 ( .A1(G2078), .A2(G2084), .ZN(n797) );
  XOR2_X1 U883 ( .A(KEYINPUT20), .B(KEYINPUT80), .Z(n796) );
  XNOR2_X1 U884 ( .A(n797), .B(n796), .ZN(n798) );
  NAND2_X1 U885 ( .A1(G2090), .A2(n798), .ZN(n799) );
  XNOR2_X1 U886 ( .A(KEYINPUT21), .B(n799), .ZN(n800) );
  NAND2_X1 U887 ( .A1(n800), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U888 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U889 ( .A1(G220), .A2(G219), .ZN(n801) );
  XOR2_X1 U890 ( .A(KEYINPUT22), .B(n801), .Z(n802) );
  NOR2_X1 U891 ( .A1(G218), .A2(n802), .ZN(n803) );
  NAND2_X1 U892 ( .A1(G96), .A2(n803), .ZN(n818) );
  NAND2_X1 U893 ( .A1(G2106), .A2(n818), .ZN(n808) );
  NAND2_X1 U894 ( .A1(G120), .A2(G108), .ZN(n804) );
  NOR2_X1 U895 ( .A1(G237), .A2(n804), .ZN(n805) );
  NAND2_X1 U896 ( .A1(G69), .A2(n805), .ZN(n817) );
  NAND2_X1 U897 ( .A1(G567), .A2(n817), .ZN(n806) );
  XOR2_X1 U898 ( .A(KEYINPUT81), .B(n806), .Z(n807) );
  NAND2_X1 U899 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U900 ( .A(KEYINPUT82), .B(n809), .Z(G319) );
  INV_X1 U901 ( .A(G319), .ZN(n811) );
  NAND2_X1 U902 ( .A1(G661), .A2(G483), .ZN(n810) );
  NOR2_X1 U903 ( .A1(n811), .A2(n810), .ZN(n814) );
  NAND2_X1 U904 ( .A1(n814), .A2(G36), .ZN(G176) );
  NAND2_X1 U905 ( .A1(G2106), .A2(n812), .ZN(G217) );
  AND2_X1 U906 ( .A1(G15), .A2(G2), .ZN(n813) );
  NAND2_X1 U907 ( .A1(G661), .A2(n813), .ZN(G259) );
  NAND2_X1 U908 ( .A1(G1), .A2(G3), .ZN(n815) );
  NAND2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U910 ( .A(n816), .B(KEYINPUT98), .ZN(G188) );
  XNOR2_X1 U911 ( .A(G96), .B(KEYINPUT99), .ZN(G221) );
  XOR2_X1 U912 ( .A(G108), .B(KEYINPUT108), .Z(G238) );
  INV_X1 U914 ( .A(G120), .ZN(G236) );
  NOR2_X1 U915 ( .A1(n818), .A2(n817), .ZN(G325) );
  INV_X1 U916 ( .A(G325), .ZN(G261) );
  XOR2_X1 U917 ( .A(KEYINPUT102), .B(G1986), .Z(n820) );
  XNOR2_X1 U918 ( .A(G1971), .B(G1976), .ZN(n819) );
  XNOR2_X1 U919 ( .A(n820), .B(n819), .ZN(n821) );
  XOR2_X1 U920 ( .A(n821), .B(KEYINPUT41), .Z(n823) );
  XNOR2_X1 U921 ( .A(G1996), .B(G1991), .ZN(n822) );
  XNOR2_X1 U922 ( .A(n823), .B(n822), .ZN(n827) );
  XOR2_X1 U923 ( .A(G1961), .B(G1956), .Z(n825) );
  XNOR2_X1 U924 ( .A(G1981), .B(G1966), .ZN(n824) );
  XNOR2_X1 U925 ( .A(n825), .B(n824), .ZN(n826) );
  XOR2_X1 U926 ( .A(n827), .B(n826), .Z(n829) );
  XNOR2_X1 U927 ( .A(KEYINPUT101), .B(G2474), .ZN(n828) );
  XNOR2_X1 U928 ( .A(n829), .B(n828), .ZN(G229) );
  XOR2_X1 U929 ( .A(G2096), .B(KEYINPUT43), .Z(n831) );
  XNOR2_X1 U930 ( .A(G2067), .B(KEYINPUT100), .ZN(n830) );
  XNOR2_X1 U931 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U932 ( .A(n832), .B(G2678), .Z(n834) );
  XNOR2_X1 U933 ( .A(G2090), .B(G2072), .ZN(n833) );
  XNOR2_X1 U934 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U935 ( .A(KEYINPUT42), .B(G2100), .Z(n836) );
  XNOR2_X1 U936 ( .A(G2078), .B(G2084), .ZN(n835) );
  XNOR2_X1 U937 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(G227) );
  NAND2_X1 U939 ( .A1(n865), .A2(G124), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n839), .B(KEYINPUT44), .ZN(n841) );
  NAND2_X1 U941 ( .A1(G112), .A2(n866), .ZN(n840) );
  NAND2_X1 U942 ( .A1(n841), .A2(n840), .ZN(n845) );
  NAND2_X1 U943 ( .A1(G136), .A2(n861), .ZN(n843) );
  NAND2_X1 U944 ( .A1(G100), .A2(n862), .ZN(n842) );
  NAND2_X1 U945 ( .A1(n843), .A2(n842), .ZN(n844) );
  NOR2_X1 U946 ( .A1(n845), .A2(n844), .ZN(G162) );
  NAND2_X1 U947 ( .A1(G130), .A2(n865), .ZN(n847) );
  NAND2_X1 U948 ( .A1(G118), .A2(n866), .ZN(n846) );
  NAND2_X1 U949 ( .A1(n847), .A2(n846), .ZN(n852) );
  NAND2_X1 U950 ( .A1(G142), .A2(n861), .ZN(n849) );
  NAND2_X1 U951 ( .A1(G106), .A2(n862), .ZN(n848) );
  NAND2_X1 U952 ( .A1(n849), .A2(n848), .ZN(n850) );
  XOR2_X1 U953 ( .A(n850), .B(KEYINPUT45), .Z(n851) );
  NOR2_X1 U954 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n853), .B(G164), .ZN(n860) );
  XOR2_X1 U956 ( .A(KEYINPUT103), .B(KEYINPUT46), .Z(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U958 ( .A(n856), .B(KEYINPUT105), .Z(n858) );
  XNOR2_X1 U959 ( .A(G160), .B(KEYINPUT48), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(n877) );
  NAND2_X1 U962 ( .A1(G139), .A2(n861), .ZN(n864) );
  NAND2_X1 U963 ( .A1(G103), .A2(n862), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n872) );
  NAND2_X1 U965 ( .A1(G127), .A2(n865), .ZN(n868) );
  NAND2_X1 U966 ( .A1(G115), .A2(n866), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U968 ( .A(KEYINPUT104), .B(n869), .Z(n870) );
  XNOR2_X1 U969 ( .A(KEYINPUT47), .B(n870), .ZN(n871) );
  NOR2_X1 U970 ( .A1(n872), .A2(n871), .ZN(n999) );
  XNOR2_X1 U971 ( .A(n999), .B(G162), .ZN(n875) );
  XNOR2_X1 U972 ( .A(n873), .B(n987), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n877), .B(n876), .ZN(n879) );
  XNOR2_X1 U975 ( .A(n879), .B(n878), .ZN(n880) );
  NOR2_X1 U976 ( .A1(G37), .A2(n880), .ZN(G395) );
  XNOR2_X1 U977 ( .A(G286), .B(n881), .ZN(n883) );
  XNOR2_X1 U978 ( .A(n942), .B(n939), .ZN(n882) );
  XNOR2_X1 U979 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U980 ( .A(n884), .B(G301), .ZN(n885) );
  NOR2_X1 U981 ( .A1(G37), .A2(n885), .ZN(n886) );
  XNOR2_X1 U982 ( .A(KEYINPUT106), .B(n886), .ZN(G397) );
  XOR2_X1 U983 ( .A(G2451), .B(G2430), .Z(n888) );
  XNOR2_X1 U984 ( .A(G2438), .B(G2443), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n888), .B(n887), .ZN(n894) );
  XOR2_X1 U986 ( .A(G2435), .B(G2454), .Z(n890) );
  XNOR2_X1 U987 ( .A(G1341), .B(G1348), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n892) );
  XOR2_X1 U989 ( .A(G2446), .B(G2427), .Z(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U991 ( .A(n894), .B(n893), .Z(n895) );
  NAND2_X1 U992 ( .A1(G14), .A2(n895), .ZN(n902) );
  NAND2_X1 U993 ( .A1(n902), .A2(G319), .ZN(n899) );
  NOR2_X1 U994 ( .A1(G229), .A2(G227), .ZN(n896) );
  XOR2_X1 U995 ( .A(KEYINPUT107), .B(n896), .Z(n897) );
  XNOR2_X1 U996 ( .A(n897), .B(KEYINPUT49), .ZN(n898) );
  NOR2_X1 U997 ( .A1(n899), .A2(n898), .ZN(n901) );
  NOR2_X1 U998 ( .A1(G395), .A2(G397), .ZN(n900) );
  NAND2_X1 U999 ( .A1(n901), .A2(n900), .ZN(G225) );
  INV_X1 U1000 ( .A(G225), .ZN(G308) );
  INV_X1 U1001 ( .A(G69), .ZN(G235) );
  INV_X1 U1002 ( .A(n902), .ZN(G401) );
  XOR2_X1 U1003 ( .A(G34), .B(KEYINPUT117), .Z(n904) );
  XNOR2_X1 U1004 ( .A(G2084), .B(KEYINPUT54), .ZN(n903) );
  XNOR2_X1 U1005 ( .A(n904), .B(n903), .ZN(n923) );
  XNOR2_X1 U1006 ( .A(G2072), .B(G33), .ZN(n906) );
  XNOR2_X1 U1007 ( .A(G1991), .B(G25), .ZN(n905) );
  NOR2_X1 U1008 ( .A1(n906), .A2(n905), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(G32), .B(n907), .ZN(n908) );
  NAND2_X1 U1010 ( .A1(n908), .A2(G28), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(KEYINPUT114), .B(G2067), .ZN(n909) );
  XNOR2_X1 U1012 ( .A(G26), .B(n909), .ZN(n910) );
  NOR2_X1 U1013 ( .A1(n911), .A2(n910), .ZN(n912) );
  NAND2_X1 U1014 ( .A1(n913), .A2(n912), .ZN(n916) );
  XOR2_X1 U1015 ( .A(G27), .B(n914), .Z(n915) );
  NOR2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n917) );
  XOR2_X1 U1017 ( .A(n917), .B(KEYINPUT115), .Z(n918) );
  XNOR2_X1 U1018 ( .A(KEYINPUT53), .B(n918), .ZN(n920) );
  XNOR2_X1 U1019 ( .A(G35), .B(G2090), .ZN(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1021 ( .A(KEYINPUT116), .B(n921), .Z(n922) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(KEYINPUT55), .B(KEYINPUT113), .ZN(n1011) );
  XNOR2_X1 U1024 ( .A(n924), .B(n1011), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(n925), .B(KEYINPUT118), .ZN(n926) );
  NOR2_X1 U1026 ( .A1(G29), .A2(n926), .ZN(n927) );
  XNOR2_X1 U1027 ( .A(KEYINPUT119), .B(n927), .ZN(n928) );
  NAND2_X1 U1028 ( .A1(n928), .A2(G11), .ZN(n929) );
  XNOR2_X1 U1029 ( .A(n929), .B(KEYINPUT120), .ZN(n1017) );
  XOR2_X1 U1030 ( .A(G16), .B(KEYINPUT56), .Z(n955) );
  XNOR2_X1 U1031 ( .A(G166), .B(G1971), .ZN(n937) );
  INV_X1 U1032 ( .A(n930), .ZN(n931) );
  NAND2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1034 ( .A(KEYINPUT121), .B(n933), .Z(n935) );
  XNOR2_X1 U1035 ( .A(G1956), .B(G299), .ZN(n934) );
  NOR2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(n938), .B(KEYINPUT122), .ZN(n953) );
  XNOR2_X1 U1039 ( .A(n939), .B(G1348), .ZN(n941) );
  NAND2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n946) );
  XOR2_X1 U1041 ( .A(n942), .B(G1341), .Z(n944) );
  XNOR2_X1 U1042 ( .A(G171), .B(G1961), .ZN(n943) );
  NAND2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(G1966), .B(G168), .ZN(n948) );
  NAND2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(n949), .B(KEYINPUT57), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n984) );
  XOR2_X1 U1051 ( .A(G1986), .B(G24), .Z(n958) );
  XNOR2_X1 U1052 ( .A(G1976), .B(KEYINPUT125), .ZN(n956) );
  XNOR2_X1 U1053 ( .A(n956), .B(G23), .ZN(n957) );
  NAND2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(G22), .B(G1971), .ZN(n959) );
  NOR2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1057 ( .A(KEYINPUT58), .B(n961), .Z(n979) );
  XOR2_X1 U1058 ( .A(G1966), .B(G21), .Z(n964) );
  XNOR2_X1 U1059 ( .A(n962), .B(G5), .ZN(n963) );
  NAND2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n976) );
  XNOR2_X1 U1061 ( .A(KEYINPUT59), .B(G1348), .ZN(n965) );
  XNOR2_X1 U1062 ( .A(n965), .B(G4), .ZN(n972) );
  XOR2_X1 U1063 ( .A(G1341), .B(G19), .Z(n968) );
  XNOR2_X1 U1064 ( .A(n966), .B(G20), .ZN(n967) );
  NAND2_X1 U1065 ( .A1(n968), .A2(n967), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(G6), .B(G1981), .ZN(n969) );
  NOR2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1069 ( .A(KEYINPUT123), .B(n973), .Z(n974) );
  XNOR2_X1 U1070 ( .A(KEYINPUT60), .B(n974), .ZN(n975) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1072 ( .A(KEYINPUT124), .B(n977), .Z(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1074 ( .A(KEYINPUT61), .B(n980), .Z(n981) );
  NOR2_X1 U1075 ( .A1(G16), .A2(n981), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(KEYINPUT126), .B(n982), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n1015) );
  XNOR2_X1 U1078 ( .A(G2084), .B(G160), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(KEYINPUT109), .B(n985), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n991) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(KEYINPUT110), .B(n992), .ZN(n1009) );
  XOR2_X1 U1084 ( .A(G2090), .B(G162), .Z(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1086 ( .A(n995), .B(KEYINPUT111), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(n996), .B(KEYINPUT51), .ZN(n998) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n1005) );
  XOR2_X1 U1089 ( .A(G164), .B(G2078), .Z(n1002) );
  XOR2_X1 U1090 ( .A(n999), .B(KEYINPUT112), .Z(n1000) );
  XNOR2_X1 U1091 ( .A(G2072), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1093 ( .A(KEYINPUT50), .B(n1003), .Z(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(KEYINPUT52), .B(n1010), .ZN(n1012) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(G29), .ZN(n1014) );
  NAND2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1101 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1102 ( .A(KEYINPUT127), .B(n1018), .Z(n1019) );
  XNOR2_X1 U1103 ( .A(KEYINPUT62), .B(n1019), .ZN(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

