

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742;

  AND2_X2 U369 ( .A1(n609), .A2(n608), .ZN(n705) );
  AND2_X1 U370 ( .A1(n536), .A2(n574), .ZN(n526) );
  AND2_X1 U371 ( .A1(n386), .A2(n668), .ZN(n382) );
  AND2_X1 U372 ( .A1(n522), .A2(n387), .ZN(n386) );
  XNOR2_X1 U373 ( .A(n446), .B(n445), .ZN(n563) );
  XNOR2_X1 U374 ( .A(n429), .B(n352), .ZN(n490) );
  XNOR2_X2 U375 ( .A(G125), .B(G146), .ZN(n482) );
  XNOR2_X2 U376 ( .A(n369), .B(n379), .ZN(n725) );
  XNOR2_X2 U377 ( .A(n485), .B(G134), .ZN(n379) );
  NOR2_X2 U378 ( .A1(n649), .A2(n537), .ZN(n416) );
  INV_X1 U379 ( .A(G953), .ZN(n732) );
  AND2_X2 U380 ( .A1(n731), .A2(n599), .ZN(n383) );
  XNOR2_X2 U381 ( .A(n368), .B(KEYINPUT77), .ZN(n397) );
  XNOR2_X2 U382 ( .A(n526), .B(n525), .ZN(n649) );
  OR2_X2 U383 ( .A1(n618), .A2(G902), .ZN(n474) );
  XNOR2_X2 U384 ( .A(n516), .B(KEYINPUT40), .ZN(n568) );
  XNOR2_X2 U385 ( .A(n473), .B(n461), .ZN(n701) );
  XNOR2_X1 U386 ( .A(KEYINPUT65), .B(KEYINPUT68), .ZN(n455) );
  NAND2_X1 U387 ( .A1(n606), .A2(n605), .ZN(n609) );
  BUF_X1 U388 ( .A(n527), .Z(n528) );
  XNOR2_X1 U389 ( .A(n515), .B(n514), .ZN(n635) );
  XNOR2_X1 U390 ( .A(n476), .B(n381), .ZN(n380) );
  XOR2_X1 U391 ( .A(n694), .B(n693), .Z(n695) );
  XNOR2_X1 U392 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U393 ( .A(n455), .B(KEYINPUT4), .ZN(n484) );
  XNOR2_X2 U394 ( .A(n367), .B(n489), .ZN(n585) );
  NOR2_X1 U395 ( .A1(n580), .A2(n346), .ZN(n363) );
  XNOR2_X1 U396 ( .A(n395), .B(KEYINPUT74), .ZN(n362) );
  INV_X1 U397 ( .A(n644), .ZN(n359) );
  XNOR2_X1 U398 ( .A(n484), .B(G137), .ZN(n369) );
  XOR2_X1 U399 ( .A(G122), .B(KEYINPUT9), .Z(n506) );
  NOR2_X1 U400 ( .A1(n361), .A2(n359), .ZN(n581) );
  XOR2_X1 U401 ( .A(G131), .B(G140), .Z(n491) );
  NAND2_X1 U402 ( .A1(G898), .A2(G953), .ZN(n521) );
  XNOR2_X1 U403 ( .A(n473), .B(n472), .ZN(n618) );
  XNOR2_X1 U404 ( .A(G143), .B(G122), .ZN(n492) );
  XOR2_X1 U405 ( .A(KEYINPUT12), .B(KEYINPUT104), .Z(n493) );
  XNOR2_X1 U406 ( .A(n495), .B(n494), .ZN(n496) );
  INV_X1 U407 ( .A(KEYINPUT11), .ZN(n494) );
  XNOR2_X1 U408 ( .A(G113), .B(G104), .ZN(n495) );
  NOR2_X1 U409 ( .A1(G953), .A2(G237), .ZN(n498) );
  NAND2_X1 U410 ( .A1(n397), .A2(n659), .ZN(n367) );
  AND2_X1 U411 ( .A1(n426), .A2(n635), .ZN(n425) );
  AND2_X1 U412 ( .A1(n574), .A2(n573), .ZN(n426) );
  XNOR2_X1 U413 ( .A(n519), .B(n518), .ZN(n576) );
  INV_X1 U414 ( .A(KEYINPUT91), .ZN(n518) );
  XNOR2_X1 U415 ( .A(n564), .B(n366), .ZN(n365) );
  INV_X1 U416 ( .A(KEYINPUT28), .ZN(n366) );
  XNOR2_X1 U417 ( .A(n576), .B(n520), .ZN(n572) );
  INV_X1 U418 ( .A(KEYINPUT19), .ZN(n520) );
  XNOR2_X1 U419 ( .A(n531), .B(n424), .ZN(n544) );
  INV_X1 U420 ( .A(KEYINPUT22), .ZN(n424) );
  NOR2_X1 U421 ( .A1(n537), .A2(n530), .ZN(n531) );
  NAND2_X1 U422 ( .A1(n705), .A2(n401), .ZN(n400) );
  AND2_X1 U423 ( .A1(n706), .A2(G478), .ZN(n401) );
  INV_X1 U424 ( .A(n714), .ZN(n403) );
  OR2_X1 U425 ( .A1(n706), .A2(G478), .ZN(n399) );
  XOR2_X1 U426 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n569) );
  NOR2_X1 U427 ( .A1(n631), .A2(n635), .ZN(n664) );
  XOR2_X1 U428 ( .A(KEYINPUT86), .B(KEYINPUT48), .Z(n583) );
  XNOR2_X1 U429 ( .A(G131), .B(G101), .ZN(n466) );
  NAND2_X1 U430 ( .A1(n372), .A2(KEYINPUT88), .ZN(n371) );
  NAND2_X1 U431 ( .A1(n737), .A2(KEYINPUT44), .ZN(n372) );
  AND2_X1 U432 ( .A1(n377), .A2(n375), .ZN(n374) );
  AND2_X1 U433 ( .A1(n378), .A2(KEYINPUT44), .ZN(n376) );
  XOR2_X1 U434 ( .A(KEYINPUT8), .B(n434), .Z(n504) );
  NAND2_X1 U435 ( .A1(n732), .A2(G234), .ZN(n434) );
  XNOR2_X1 U436 ( .A(n370), .B(n523), .ZN(n536) );
  INV_X1 U437 ( .A(KEYINPUT76), .ZN(n523) );
  INV_X1 U438 ( .A(G237), .ZN(n475) );
  INV_X1 U439 ( .A(n559), .ZN(n387) );
  INV_X1 U440 ( .A(KEYINPUT30), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n522), .B(KEYINPUT1), .ZN(n527) );
  XNOR2_X1 U442 ( .A(G113), .B(KEYINPUT71), .ZN(n463) );
  INV_X1 U443 ( .A(G122), .ZN(n478) );
  XOR2_X1 U444 ( .A(KEYINPUT98), .B(G140), .Z(n436) );
  XNOR2_X1 U445 ( .A(n490), .B(n431), .ZN(n432) );
  XNOR2_X1 U446 ( .A(G119), .B(G110), .ZN(n430) );
  XNOR2_X1 U447 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U448 ( .A(G116), .B(G107), .ZN(n508) );
  INV_X1 U449 ( .A(n608), .ZN(n654) );
  INV_X1 U450 ( .A(KEYINPUT0), .ZN(n408) );
  NOR2_X1 U451 ( .A1(n572), .A2(n422), .ZN(n407) );
  NAND2_X1 U452 ( .A1(n517), .A2(n521), .ZN(n422) );
  BUF_X1 U453 ( .A(n673), .Z(n388) );
  XNOR2_X1 U454 ( .A(n418), .B(n479), .ZN(n719) );
  XNOR2_X1 U455 ( .A(n477), .B(n419), .ZN(n418) );
  XNOR2_X1 U456 ( .A(n478), .B(n420), .ZN(n419) );
  INV_X1 U457 ( .A(KEYINPUT16), .ZN(n420) );
  XNOR2_X1 U458 ( .A(n497), .B(n496), .ZN(n500) );
  AND2_X1 U459 ( .A1(n614), .A2(G953), .ZN(n714) );
  NAND2_X1 U460 ( .A1(n585), .A2(n635), .ZN(n516) );
  NAND2_X1 U461 ( .A1(n360), .A2(n578), .ZN(n644) );
  XNOR2_X1 U462 ( .A(n577), .B(KEYINPUT36), .ZN(n360) );
  NOR2_X1 U463 ( .A1(n544), .A2(n351), .ZN(n390) );
  XNOR2_X1 U464 ( .A(n364), .B(KEYINPUT80), .ZN(n636) );
  NOR2_X1 U465 ( .A1(n411), .A2(n574), .ZN(n409) );
  NOR2_X1 U466 ( .A1(n402), .A2(n398), .ZN(n707) );
  NOR2_X1 U467 ( .A1(n708), .A2(n706), .ZN(n402) );
  INV_X1 U468 ( .A(KEYINPUT53), .ZN(n391) );
  INV_X1 U469 ( .A(n563), .ZN(n411) );
  AND2_X1 U470 ( .A1(n579), .A2(KEYINPUT47), .ZN(n346) );
  NOR2_X1 U471 ( .A1(n417), .A2(KEYINPUT2), .ZN(n347) );
  AND2_X1 U472 ( .A1(n487), .A2(G210), .ZN(n348) );
  OR2_X1 U473 ( .A1(G953), .A2(n651), .ZN(n349) );
  AND2_X1 U474 ( .A1(n563), .A2(n671), .ZN(n668) );
  AND2_X1 U475 ( .A1(n541), .A2(n396), .ZN(n350) );
  OR2_X1 U476 ( .A1(n423), .A2(n574), .ZN(n351) );
  XOR2_X1 U477 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n352) );
  AND2_X1 U478 ( .A1(n529), .A2(n539), .ZN(n353) );
  NAND2_X1 U479 ( .A1(n542), .A2(n541), .ZN(n354) );
  AND2_X1 U480 ( .A1(n353), .A2(n389), .ZN(n355) );
  AND2_X1 U481 ( .A1(n652), .A2(KEYINPUT2), .ZN(n356) );
  XOR2_X1 U482 ( .A(KEYINPUT75), .B(KEYINPUT38), .Z(n357) );
  XNOR2_X1 U483 ( .A(n510), .B(n384), .ZN(n706) );
  AND2_X1 U484 ( .A1(n399), .A2(n403), .ZN(n358) );
  NAND2_X1 U485 ( .A1(n363), .A2(n362), .ZN(n361) );
  NOR2_X1 U486 ( .A1(n572), .A2(n571), .ZN(n364) );
  NAND2_X1 U487 ( .A1(n365), .A2(n522), .ZN(n571) );
  NAND2_X1 U488 ( .A1(n382), .A2(n380), .ZN(n368) );
  XNOR2_X2 U489 ( .A(n725), .B(G146), .ZN(n473) );
  NAND2_X1 U490 ( .A1(n417), .A2(n356), .ZN(n608) );
  NAND2_X1 U491 ( .A1(n527), .A2(n668), .ZN(n370) );
  XNOR2_X2 U492 ( .A(n462), .B(G469), .ZN(n522) );
  OR2_X2 U493 ( .A1(n371), .A2(n543), .ZN(n373) );
  NAND2_X1 U494 ( .A1(n374), .A2(n373), .ZN(n554) );
  NAND2_X1 U495 ( .A1(n737), .A2(n376), .ZN(n375) );
  NAND2_X1 U496 ( .A1(n543), .A2(n378), .ZN(n377) );
  INV_X1 U497 ( .A(KEYINPUT88), .ZN(n378) );
  XNOR2_X1 U498 ( .A(n379), .B(n509), .ZN(n384) );
  NAND2_X1 U499 ( .A1(n383), .A2(n417), .ZN(n606) );
  BUF_X2 U500 ( .A(n705), .Z(n708) );
  XNOR2_X1 U501 ( .A(n390), .B(KEYINPUT32), .ZN(n740) );
  NAND2_X1 U502 ( .A1(n578), .A2(n411), .ZN(n423) );
  NAND2_X1 U503 ( .A1(n594), .A2(n593), .ZN(n607) );
  XNOR2_X1 U504 ( .A(n482), .B(n480), .ZN(n406) );
  NAND2_X1 U505 ( .A1(n385), .A2(n354), .ZN(n543) );
  INV_X1 U506 ( .A(n624), .ZN(n385) );
  NAND2_X1 U507 ( .A1(n410), .A2(n409), .ZN(n532) );
  INV_X1 U508 ( .A(n389), .ZN(n590) );
  NAND2_X1 U509 ( .A1(n389), .A2(n658), .ZN(n519) );
  XNOR2_X2 U510 ( .A(n488), .B(n348), .ZN(n389) );
  XNOR2_X1 U511 ( .A(n590), .B(n357), .ZN(n659) );
  XNOR2_X1 U512 ( .A(n392), .B(n391), .ZN(G75) );
  NAND2_X1 U513 ( .A1(n394), .A2(n393), .ZN(n392) );
  NOR2_X1 U514 ( .A1(n689), .A2(n349), .ZN(n393) );
  NAND2_X1 U515 ( .A1(n656), .A2(n655), .ZN(n394) );
  NAND2_X1 U516 ( .A1(n636), .A2(n541), .ZN(n579) );
  NAND2_X1 U517 ( .A1(n636), .A2(n350), .ZN(n395) );
  INV_X1 U518 ( .A(KEYINPUT47), .ZN(n396) );
  AND2_X1 U519 ( .A1(n397), .A2(n355), .ZN(n634) );
  NAND2_X1 U520 ( .A1(n400), .A2(n358), .ZN(n398) );
  XNOR2_X1 U521 ( .A(n404), .B(n483), .ZN(n405) );
  XNOR2_X1 U522 ( .A(n406), .B(n481), .ZN(n404) );
  XNOR2_X1 U523 ( .A(n405), .B(n486), .ZN(n421) );
  XNOR2_X2 U524 ( .A(n407), .B(n408), .ZN(n537) );
  INV_X1 U525 ( .A(n544), .ZN(n410) );
  XNOR2_X2 U526 ( .A(n413), .B(n412), .ZN(n485) );
  XNOR2_X2 U527 ( .A(KEYINPUT66), .B(KEYINPUT81), .ZN(n412) );
  XNOR2_X2 U528 ( .A(G143), .B(G128), .ZN(n413) );
  XNOR2_X2 U529 ( .A(n414), .B(KEYINPUT35), .ZN(n737) );
  NAND2_X1 U530 ( .A1(n415), .A2(n353), .ZN(n414) );
  XNOR2_X1 U531 ( .A(n416), .B(KEYINPUT34), .ZN(n415) );
  NAND2_X1 U532 ( .A1(n417), .A2(n732), .ZN(n717) );
  XNOR2_X2 U533 ( .A(n555), .B(KEYINPUT45), .ZN(n417) );
  XNOR2_X1 U534 ( .A(n421), .B(n719), .ZN(n692) );
  NAND2_X1 U535 ( .A1(n692), .A2(n595), .ZN(n488) );
  XNOR2_X1 U536 ( .A(n547), .B(KEYINPUT90), .ZN(n548) );
  INV_X1 U537 ( .A(KEYINPUT7), .ZN(n507) );
  XNOR2_X1 U538 ( .A(n430), .B(KEYINPUT24), .ZN(n431) );
  XNOR2_X1 U539 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U540 ( .A(n503), .B(n502), .ZN(n539) );
  XNOR2_X1 U541 ( .A(n712), .B(n711), .ZN(n713) );
  XOR2_X1 U542 ( .A(KEYINPUT97), .B(KEYINPUT99), .Z(n428) );
  XNOR2_X1 U543 ( .A(KEYINPUT72), .B(KEYINPUT23), .ZN(n427) );
  XNOR2_X1 U544 ( .A(n428), .B(n427), .ZN(n433) );
  INV_X1 U545 ( .A(n482), .ZN(n429) );
  XOR2_X1 U546 ( .A(n433), .B(n432), .Z(n440) );
  NAND2_X1 U547 ( .A1(G221), .A2(n504), .ZN(n438) );
  XNOR2_X1 U548 ( .A(G128), .B(G137), .ZN(n435) );
  XNOR2_X1 U549 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U550 ( .A(n440), .B(n439), .ZN(n710) );
  NOR2_X1 U551 ( .A1(G902), .A2(n710), .ZN(n446) );
  XOR2_X1 U552 ( .A(KEYINPUT101), .B(KEYINPUT25), .Z(n443) );
  XNOR2_X1 U553 ( .A(G902), .B(KEYINPUT15), .ZN(n595) );
  NAND2_X1 U554 ( .A1(n595), .A2(G234), .ZN(n441) );
  XNOR2_X1 U555 ( .A(n441), .B(KEYINPUT20), .ZN(n447) );
  NAND2_X1 U556 ( .A1(n447), .A2(G217), .ZN(n442) );
  XNOR2_X1 U557 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U558 ( .A(KEYINPUT100), .B(n444), .ZN(n445) );
  XOR2_X1 U559 ( .A(KEYINPUT102), .B(KEYINPUT21), .Z(n449) );
  NAND2_X1 U560 ( .A1(n447), .A2(G221), .ZN(n448) );
  XNOR2_X1 U561 ( .A(n449), .B(n448), .ZN(n671) );
  INV_X1 U562 ( .A(n668), .ZN(n533) );
  NAND2_X1 U563 ( .A1(G237), .A2(G234), .ZN(n450) );
  XNOR2_X1 U564 ( .A(n450), .B(KEYINPUT14), .ZN(n657) );
  OR2_X1 U565 ( .A1(n732), .A2(G902), .ZN(n451) );
  NAND2_X1 U566 ( .A1(n657), .A2(n451), .ZN(n453) );
  NOR2_X1 U567 ( .A1(G953), .A2(G952), .ZN(n452) );
  NOR2_X1 U568 ( .A1(n453), .A2(n452), .ZN(n517) );
  NAND2_X1 U569 ( .A1(G953), .A2(G900), .ZN(n454) );
  NAND2_X1 U570 ( .A1(n517), .A2(n454), .ZN(n559) );
  XOR2_X1 U571 ( .A(G101), .B(G104), .Z(n457) );
  XNOR2_X1 U572 ( .A(G107), .B(G110), .ZN(n456) );
  XNOR2_X1 U573 ( .A(n457), .B(n456), .ZN(n477) );
  XOR2_X1 U574 ( .A(n491), .B(KEYINPUT78), .Z(n459) );
  NAND2_X1 U575 ( .A1(G227), .A2(n732), .ZN(n458) );
  XNOR2_X1 U576 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U577 ( .A(n477), .B(n460), .ZN(n461) );
  OR2_X2 U578 ( .A1(n701), .A2(G902), .ZN(n462) );
  XNOR2_X1 U579 ( .A(n463), .B(G116), .ZN(n465) );
  XOR2_X1 U580 ( .A(KEYINPUT3), .B(G119), .Z(n464) );
  XNOR2_X1 U581 ( .A(n465), .B(n464), .ZN(n479) );
  NAND2_X1 U582 ( .A1(n498), .A2(G210), .ZN(n467) );
  XNOR2_X1 U583 ( .A(n467), .B(n466), .ZN(n470) );
  INV_X1 U584 ( .A(KEYINPUT103), .ZN(n468) );
  XNOR2_X1 U585 ( .A(n468), .B(KEYINPUT5), .ZN(n469) );
  XNOR2_X1 U586 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U587 ( .A(n479), .B(n471), .ZN(n472) );
  XNOR2_X2 U588 ( .A(n474), .B(G472), .ZN(n673) );
  INV_X1 U589 ( .A(G902), .ZN(n511) );
  NAND2_X1 U590 ( .A1(n511), .A2(n475), .ZN(n487) );
  NAND2_X1 U591 ( .A1(n487), .A2(G214), .ZN(n658) );
  NAND2_X1 U592 ( .A1(n673), .A2(n658), .ZN(n476) );
  XOR2_X1 U593 ( .A(KEYINPUT17), .B(KEYINPUT96), .Z(n481) );
  XNOR2_X1 U594 ( .A(KEYINPUT79), .B(KEYINPUT18), .ZN(n480) );
  NAND2_X1 U595 ( .A1(G224), .A2(n732), .ZN(n483) );
  XNOR2_X1 U596 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U597 ( .A(KEYINPUT87), .B(KEYINPUT39), .Z(n489) );
  XNOR2_X1 U598 ( .A(KEYINPUT13), .B(G475), .ZN(n503) );
  XNOR2_X1 U599 ( .A(n491), .B(n490), .ZN(n723) );
  XNOR2_X1 U600 ( .A(n493), .B(n492), .ZN(n497) );
  NAND2_X1 U601 ( .A1(n498), .A2(G214), .ZN(n499) );
  XNOR2_X1 U602 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U603 ( .A(n723), .B(n501), .Z(n611) );
  NOR2_X1 U604 ( .A1(G902), .A2(n611), .ZN(n502) );
  NAND2_X1 U605 ( .A1(G217), .A2(n504), .ZN(n505) );
  XNOR2_X1 U606 ( .A(n506), .B(n505), .ZN(n510) );
  NAND2_X1 U607 ( .A1(n706), .A2(n511), .ZN(n513) );
  INV_X1 U608 ( .A(G478), .ZN(n512) );
  XNOR2_X1 U609 ( .A(n513), .B(n512), .ZN(n540) );
  AND2_X1 U610 ( .A1(n539), .A2(n540), .ZN(n515) );
  INV_X1 U611 ( .A(KEYINPUT105), .ZN(n514) );
  XNOR2_X1 U612 ( .A(n568), .B(G131), .ZN(G33) );
  INV_X1 U613 ( .A(n540), .ZN(n529) );
  INV_X1 U614 ( .A(KEYINPUT6), .ZN(n524) );
  XNOR2_X1 U615 ( .A(n673), .B(n524), .ZN(n574) );
  XOR2_X1 U616 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n525) );
  NOR2_X1 U617 ( .A1(n529), .A2(n539), .ZN(n556) );
  NAND2_X1 U618 ( .A1(n671), .A2(n556), .ZN(n530) );
  NOR2_X1 U619 ( .A1(n528), .A2(n532), .ZN(n624) );
  NOR2_X1 U620 ( .A1(n533), .A2(n388), .ZN(n534) );
  NAND2_X1 U621 ( .A1(n534), .A2(n522), .ZN(n535) );
  OR2_X1 U622 ( .A1(n537), .A2(n535), .ZN(n626) );
  NAND2_X1 U623 ( .A1(n536), .A2(n388), .ZN(n677) );
  NOR2_X1 U624 ( .A1(n537), .A2(n677), .ZN(n538) );
  XNOR2_X1 U625 ( .A(n538), .B(KEYINPUT31), .ZN(n641) );
  NAND2_X1 U626 ( .A1(n626), .A2(n641), .ZN(n542) );
  NOR2_X1 U627 ( .A1(n540), .A2(n539), .ZN(n631) );
  INV_X1 U628 ( .A(n664), .ZN(n541) );
  NOR2_X1 U629 ( .A1(n544), .A2(n528), .ZN(n545) );
  NAND2_X1 U630 ( .A1(n411), .A2(n545), .ZN(n546) );
  NOR2_X1 U631 ( .A1(n546), .A2(n388), .ZN(n630) );
  XNOR2_X1 U632 ( .A(n528), .B(KEYINPUT94), .ZN(n578) );
  NOR2_X1 U633 ( .A1(n630), .A2(n740), .ZN(n549) );
  NOR2_X1 U634 ( .A1(KEYINPUT44), .A2(KEYINPUT89), .ZN(n547) );
  XNOR2_X1 U635 ( .A(n549), .B(n548), .ZN(n552) );
  INV_X1 U636 ( .A(KEYINPUT44), .ZN(n550) );
  NAND2_X1 U637 ( .A1(n550), .A2(n737), .ZN(n551) );
  NAND2_X1 U638 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U639 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U640 ( .A1(n659), .A2(n658), .ZN(n663) );
  INV_X1 U641 ( .A(n556), .ZN(n662) );
  NOR2_X1 U642 ( .A1(n663), .A2(n662), .ZN(n558) );
  XNOR2_X1 U643 ( .A(KEYINPUT106), .B(KEYINPUT41), .ZN(n557) );
  XNOR2_X1 U644 ( .A(n558), .B(n557), .ZN(n682) );
  INV_X1 U645 ( .A(n671), .ZN(n560) );
  NOR2_X1 U646 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U647 ( .A(KEYINPUT70), .B(n561), .Z(n562) );
  NOR2_X1 U648 ( .A1(n563), .A2(n562), .ZN(n573) );
  NAND2_X1 U649 ( .A1(n573), .A2(n673), .ZN(n564) );
  NOR2_X1 U650 ( .A1(n682), .A2(n571), .ZN(n567) );
  XNOR2_X1 U651 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n566) );
  XNOR2_X1 U652 ( .A(n567), .B(n566), .ZN(n741) );
  NAND2_X1 U653 ( .A1(n568), .A2(n741), .ZN(n570) );
  XNOR2_X1 U654 ( .A(n570), .B(n569), .ZN(n582) );
  XOR2_X1 U655 ( .A(KEYINPUT108), .B(n425), .Z(n575) );
  NOR2_X1 U656 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U657 ( .A(KEYINPUT83), .B(n634), .Z(n580) );
  NAND2_X1 U658 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U659 ( .A(n584), .B(n583), .ZN(n594) );
  NAND2_X1 U660 ( .A1(n585), .A2(n631), .ZN(n586) );
  XOR2_X1 U661 ( .A(KEYINPUT109), .B(n586), .Z(n736) );
  INV_X1 U662 ( .A(n736), .ZN(n592) );
  NAND2_X1 U663 ( .A1(n425), .A2(n658), .ZN(n587) );
  NOR2_X1 U664 ( .A1(n528), .A2(n587), .ZN(n589) );
  INV_X1 U665 ( .A(KEYINPUT43), .ZN(n588) );
  XNOR2_X1 U666 ( .A(n589), .B(n588), .ZN(n591) );
  AND2_X1 U667 ( .A1(n591), .A2(n590), .ZN(n647) );
  NOR2_X1 U668 ( .A1(n592), .A2(n647), .ZN(n593) );
  XNOR2_X2 U669 ( .A(n607), .B(KEYINPUT85), .ZN(n731) );
  INV_X1 U670 ( .A(n595), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n597), .A2(KEYINPUT2), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n596), .A2(KEYINPUT67), .ZN(n601) );
  INV_X1 U673 ( .A(n601), .ZN(n598) );
  OR2_X1 U674 ( .A1(n598), .A2(n597), .ZN(n599) );
  INV_X1 U675 ( .A(n599), .ZN(n604) );
  INV_X1 U676 ( .A(KEYINPUT67), .ZN(n600) );
  NAND2_X1 U677 ( .A1(n600), .A2(KEYINPUT2), .ZN(n602) );
  AND2_X1 U678 ( .A1(n602), .A2(n601), .ZN(n603) );
  OR2_X1 U679 ( .A1(n604), .A2(n603), .ZN(n605) );
  INV_X1 U680 ( .A(n607), .ZN(n652) );
  NAND2_X1 U681 ( .A1(n705), .A2(G475), .ZN(n613) );
  XNOR2_X1 U682 ( .A(KEYINPUT119), .B(KEYINPUT59), .ZN(n610) );
  XNOR2_X1 U683 ( .A(n613), .B(n612), .ZN(n615) );
  INV_X1 U684 ( .A(G952), .ZN(n614) );
  NOR2_X2 U685 ( .A1(n615), .A2(n714), .ZN(n616) );
  XNOR2_X1 U686 ( .A(n616), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U687 ( .A1(n705), .A2(G472), .ZN(n620) );
  XOR2_X1 U688 ( .A(KEYINPUT62), .B(KEYINPUT93), .Z(n617) );
  XNOR2_X1 U689 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U690 ( .A(n620), .B(n619), .ZN(n621) );
  NOR2_X2 U691 ( .A1(n621), .A2(n714), .ZN(n623) );
  XNOR2_X1 U692 ( .A(KEYINPUT95), .B(KEYINPUT63), .ZN(n622) );
  XNOR2_X1 U693 ( .A(n623), .B(n622), .ZN(G57) );
  XOR2_X1 U694 ( .A(G101), .B(n624), .Z(G3) );
  INV_X1 U695 ( .A(n635), .ZN(n638) );
  NOR2_X1 U696 ( .A1(n638), .A2(n626), .ZN(n625) );
  XOR2_X1 U697 ( .A(G104), .B(n625), .Z(G6) );
  INV_X1 U698 ( .A(n631), .ZN(n642) );
  NOR2_X1 U699 ( .A1(n642), .A2(n626), .ZN(n628) );
  XNOR2_X1 U700 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U702 ( .A(G107), .B(n629), .ZN(G9) );
  XOR2_X1 U703 ( .A(G110), .B(n630), .Z(G12) );
  XOR2_X1 U704 ( .A(G128), .B(KEYINPUT29), .Z(n633) );
  NAND2_X1 U705 ( .A1(n631), .A2(n636), .ZN(n632) );
  XNOR2_X1 U706 ( .A(n633), .B(n632), .ZN(G30) );
  XOR2_X1 U707 ( .A(G143), .B(n634), .Z(G45) );
  NAND2_X1 U708 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U709 ( .A(n637), .B(G146), .ZN(G48) );
  NOR2_X1 U710 ( .A1(n638), .A2(n641), .ZN(n639) );
  XOR2_X1 U711 ( .A(KEYINPUT110), .B(n639), .Z(n640) );
  XNOR2_X1 U712 ( .A(G113), .B(n640), .ZN(G15) );
  NOR2_X1 U713 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U714 ( .A(G116), .B(n643), .Z(G18) );
  XNOR2_X1 U715 ( .A(KEYINPUT37), .B(KEYINPUT111), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U717 ( .A(G125), .B(n646), .ZN(G27) );
  XOR2_X1 U718 ( .A(G140), .B(n647), .Z(n648) );
  XNOR2_X1 U719 ( .A(KEYINPUT112), .B(n648), .ZN(G42) );
  NOR2_X1 U720 ( .A1(n649), .A2(n682), .ZN(n650) );
  XOR2_X1 U721 ( .A(KEYINPUT117), .B(n650), .Z(n651) );
  XOR2_X1 U722 ( .A(KEYINPUT84), .B(n347), .Z(n656) );
  NOR2_X1 U723 ( .A1(n731), .A2(KEYINPUT2), .ZN(n653) );
  NOR2_X1 U724 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U725 ( .A1(G952), .A2(n657), .ZN(n687) );
  NOR2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U727 ( .A(KEYINPUT115), .B(n660), .Z(n661) );
  NOR2_X1 U728 ( .A1(n662), .A2(n661), .ZN(n666) );
  NOR2_X1 U729 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U730 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U731 ( .A1(n649), .A2(n667), .ZN(n684) );
  NOR2_X1 U732 ( .A1(n528), .A2(n668), .ZN(n669) );
  XNOR2_X1 U733 ( .A(n669), .B(KEYINPUT113), .ZN(n670) );
  XNOR2_X1 U734 ( .A(n670), .B(KEYINPUT50), .ZN(n676) );
  NOR2_X1 U735 ( .A1(n563), .A2(n671), .ZN(n672) );
  XOR2_X1 U736 ( .A(KEYINPUT49), .B(n672), .Z(n674) );
  NOR2_X1 U737 ( .A1(n674), .A2(n388), .ZN(n675) );
  NAND2_X1 U738 ( .A1(n676), .A2(n675), .ZN(n678) );
  NAND2_X1 U739 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U740 ( .A(n679), .B(KEYINPUT114), .ZN(n680) );
  XNOR2_X1 U741 ( .A(KEYINPUT51), .B(n680), .ZN(n681) );
  NOR2_X1 U742 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U743 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U744 ( .A(n685), .B(KEYINPUT52), .ZN(n686) );
  NOR2_X1 U745 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U746 ( .A(n688), .B(KEYINPUT116), .ZN(n689) );
  NAND2_X1 U747 ( .A1(n705), .A2(G210), .ZN(n696) );
  XOR2_X1 U748 ( .A(KEYINPUT92), .B(KEYINPUT82), .Z(n691) );
  XNOR2_X1 U749 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n690) );
  XNOR2_X1 U750 ( .A(n691), .B(n690), .ZN(n694) );
  BUF_X1 U751 ( .A(n692), .Z(n693) );
  XNOR2_X1 U752 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X2 U753 ( .A1(n697), .A2(n714), .ZN(n698) );
  XNOR2_X1 U754 ( .A(n698), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U755 ( .A1(n708), .A2(G469), .ZN(n703) );
  XNOR2_X1 U756 ( .A(KEYINPUT58), .B(KEYINPUT118), .ZN(n699) );
  XOR2_X1 U757 ( .A(n699), .B(KEYINPUT57), .Z(n700) );
  XNOR2_X1 U758 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U759 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U760 ( .A1(n714), .A2(n704), .ZN(G54) );
  XNOR2_X1 U761 ( .A(KEYINPUT120), .B(n707), .ZN(G63) );
  NAND2_X1 U762 ( .A1(n708), .A2(G217), .ZN(n712) );
  INV_X1 U763 ( .A(KEYINPUT121), .ZN(n709) );
  XNOR2_X1 U764 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U765 ( .A1(n714), .A2(n713), .ZN(G66) );
  NAND2_X1 U766 ( .A1(G953), .A2(G224), .ZN(n715) );
  XNOR2_X1 U767 ( .A(KEYINPUT61), .B(n715), .ZN(n716) );
  NAND2_X1 U768 ( .A1(n716), .A2(G898), .ZN(n718) );
  NAND2_X1 U769 ( .A1(n718), .A2(n717), .ZN(n722) );
  OR2_X1 U770 ( .A1(n732), .A2(G898), .ZN(n720) );
  NAND2_X1 U771 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U772 ( .A(n722), .B(n721), .Z(G69) );
  XNOR2_X1 U773 ( .A(G227), .B(KEYINPUT124), .ZN(n726) );
  XNOR2_X1 U774 ( .A(n723), .B(KEYINPUT122), .ZN(n724) );
  XOR2_X1 U775 ( .A(n725), .B(n724), .Z(n729) );
  XNOR2_X1 U776 ( .A(n726), .B(n729), .ZN(n727) );
  NAND2_X1 U777 ( .A1(n727), .A2(G900), .ZN(n728) );
  NAND2_X1 U778 ( .A1(n728), .A2(G953), .ZN(n735) );
  XNOR2_X1 U779 ( .A(n729), .B(KEYINPUT123), .ZN(n730) );
  XNOR2_X1 U780 ( .A(n731), .B(n730), .ZN(n733) );
  NAND2_X1 U781 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U782 ( .A1(n735), .A2(n734), .ZN(G72) );
  XNOR2_X1 U783 ( .A(G134), .B(n736), .ZN(G36) );
  XNOR2_X1 U784 ( .A(n737), .B(G122), .ZN(n738) );
  XNOR2_X1 U785 ( .A(n738), .B(KEYINPUT125), .ZN(G24) );
  XOR2_X1 U786 ( .A(G119), .B(KEYINPUT126), .Z(n739) );
  XNOR2_X1 U787 ( .A(n740), .B(n739), .ZN(G21) );
  XOR2_X1 U788 ( .A(G137), .B(n741), .Z(n742) );
  XNOR2_X1 U789 ( .A(KEYINPUT127), .B(n742), .ZN(G39) );
endmodule

