//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT96), .B(G952), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(G234), .A2(G237), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT21), .B(G898), .ZN(new_n192));
  NAND4_X1  g006(.A1(new_n192), .A2(G902), .A3(G953), .A4(new_n190), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT4), .ZN(new_n196));
  INV_X1    g010(.A(G104), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G107), .ZN(new_n198));
  INV_X1    g012(.A(G101), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G107), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT80), .A3(G104), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n201), .A2(KEYINPUT80), .A3(KEYINPUT3), .A4(G104), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n200), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n198), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n207), .B1(new_n204), .B2(new_n205), .ZN(new_n208));
  OAI22_X1  g022(.A1(new_n196), .A2(new_n206), .B1(new_n208), .B2(new_n199), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n204), .A2(new_n205), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(new_n198), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(KEYINPUT4), .A3(G101), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G113), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT2), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT2), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G113), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G116), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT67), .B1(new_n220), .B2(G119), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n222));
  INV_X1    g036(.A(G119), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n223), .A3(G116), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n220), .A2(G119), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n219), .A2(new_n226), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n218), .A2(new_n221), .A3(new_n224), .A4(new_n225), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n213), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n201), .A2(G104), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n199), .B1(new_n231), .B2(new_n198), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n206), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n220), .A2(G119), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT5), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n214), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n226), .B2(new_n235), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n233), .A2(new_n228), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(G110), .B(G122), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT83), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n240), .B(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n230), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT84), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n227), .A2(new_n228), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n246), .B1(new_n209), .B2(new_n212), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n245), .B1(new_n247), .B2(new_n238), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n243), .A2(new_n248), .A3(KEYINPUT6), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT6), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n250), .B(new_n245), .C1(new_n247), .C2(new_n238), .ZN(new_n251));
  INV_X1    g065(.A(G146), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G143), .ZN(new_n253));
  INV_X1    g067(.A(G143), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G146), .ZN(new_n255));
  AND2_X1   g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(G143), .B(G146), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT0), .B(G128), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n260), .A2(KEYINPUT85), .A3(G125), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT85), .B1(new_n260), .B2(G125), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT1), .B1(new_n254), .B2(G146), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n254), .A2(G146), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n252), .A2(G143), .ZN(new_n265));
  OAI211_X1 g079(.A(G128), .B(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G128), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n253), .B(new_n255), .C1(KEYINPUT1), .C2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(G125), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NOR3_X1   g083(.A1(new_n261), .A2(new_n262), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G224), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(G953), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n270), .B(new_n273), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n249), .A2(new_n251), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(KEYINPUT7), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n272), .A2(KEYINPUT86), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n277), .B1(new_n270), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n262), .A2(new_n269), .ZN(new_n280));
  INV_X1    g094(.A(new_n261), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n278), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(new_n276), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n242), .B(KEYINPUT8), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n233), .B1(new_n228), .B2(new_n237), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n285), .B1(new_n286), .B2(new_n238), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n243), .A2(new_n279), .A3(new_n284), .A4(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G210), .B1(G237), .B2(G902), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n275), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n288), .A2(new_n289), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n249), .A2(new_n274), .A3(new_n251), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n291), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n187), .B(new_n195), .C1(new_n293), .C2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(G237), .A2(G953), .ZN(new_n298));
  AND2_X1   g112(.A1(KEYINPUT88), .A2(G143), .ZN(new_n299));
  NOR2_X1   g113(.A1(KEYINPUT88), .A2(G143), .ZN(new_n300));
  OAI211_X1 g114(.A(G214), .B(new_n298), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G237), .ZN(new_n302));
  INV_X1    g116(.A(G953), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n303), .A3(G214), .ZN(new_n304));
  NAND2_X1  g118(.A1(KEYINPUT88), .A2(G143), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT18), .ZN(new_n307));
  INV_X1    g121(.A(G131), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n301), .B(new_n306), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(G125), .B(G140), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n310), .A2(new_n252), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n252), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n301), .A2(new_n306), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G131), .ZN(new_n314));
  OAI221_X1 g128(.A(new_n309), .B1(new_n311), .B2(new_n312), .C1(new_n314), .C2(new_n307), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT17), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n301), .A2(new_n308), .A3(new_n306), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n314), .A2(KEYINPUT92), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G125), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G140), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT16), .ZN(new_n323));
  OR3_X1    g137(.A1(new_n321), .A2(KEYINPUT16), .A3(G140), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n323), .A2(G146), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(G146), .B1(new_n323), .B2(new_n324), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n318), .B(new_n327), .C1(new_n316), .C2(new_n314), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n301), .A2(new_n308), .A3(new_n306), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n308), .B1(new_n301), .B2(new_n306), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT92), .B1(new_n331), .B2(new_n316), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n315), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G113), .B(G122), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(new_n197), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n335), .B(new_n315), .C1(new_n328), .C2(new_n332), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n289), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G475), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT20), .ZN(new_n342));
  NOR2_X1   g156(.A1(G475), .A2(G902), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(KEYINPUT93), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT89), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n329), .B2(new_n330), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT90), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT19), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n310), .A2(KEYINPUT90), .A3(KEYINPUT19), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n325), .B1(new_n351), .B2(new_n252), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n314), .A2(KEYINPUT89), .A3(new_n317), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n346), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n315), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(KEYINPUT91), .A3(new_n336), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n338), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT91), .B1(new_n355), .B2(new_n336), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n342), .B(new_n344), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  XOR2_X1   g174(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n361));
  NAND2_X1  g175(.A1(new_n355), .A2(new_n336), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT91), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(new_n338), .A3(new_n356), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n361), .B1(new_n365), .B2(new_n344), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n341), .B1(new_n360), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT15), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G478), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n254), .A2(G128), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n267), .A2(G143), .ZN(new_n371));
  INV_X1    g185(.A(G134), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G122), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G116), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n220), .A2(G122), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G107), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n376), .A3(new_n201), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n373), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT13), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n370), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n254), .A2(KEYINPUT13), .A3(G128), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n382), .A2(new_n383), .A3(new_n371), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n380), .B1(new_n372), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT9), .B(G234), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(KEYINPUT78), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n303), .A2(G217), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n220), .A2(KEYINPUT14), .A3(G122), .ZN(new_n390));
  OAI211_X1 g204(.A(G107), .B(new_n390), .C1(new_n377), .C2(KEYINPUT14), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n372), .B1(new_n370), .B2(new_n371), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n391), .B(new_n379), .C1(new_n373), .C2(new_n392), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n385), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n389), .B1(new_n385), .B2(new_n393), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n289), .B(new_n369), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(KEYINPUT95), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n394), .A2(new_n395), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT94), .B1(new_n398), .B2(G902), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n385), .A2(new_n393), .ZN(new_n400));
  INV_X1    g214(.A(new_n389), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n385), .A2(new_n389), .A3(new_n393), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT94), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n405), .A3(new_n289), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n399), .A2(new_n406), .A3(new_n368), .A4(G478), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n397), .A2(new_n407), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n297), .A2(new_n367), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT72), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n266), .A2(new_n268), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT65), .B1(new_n372), .B2(G137), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT11), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n372), .A2(G137), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT11), .ZN(new_n417));
  OAI211_X1 g231(.A(KEYINPUT65), .B(new_n417), .C1(new_n372), .C2(G137), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n415), .A2(new_n308), .A3(new_n416), .A4(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G137), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G134), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n416), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G131), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n413), .A2(KEYINPUT66), .A3(new_n419), .A4(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT66), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n266), .A2(new_n423), .A3(new_n268), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n418), .A2(new_n416), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n417), .B1(new_n421), .B2(KEYINPUT65), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n427), .A2(new_n428), .A3(G131), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n425), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT64), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n257), .B(new_n432), .C1(new_n258), .C2(new_n259), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(KEYINPUT0), .A2(G128), .ZN(new_n435));
  OR2_X1    g249(.A1(KEYINPUT0), .A2(G128), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n435), .B(new_n436), .C1(new_n264), .C2(new_n265), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n432), .B1(new_n437), .B2(new_n257), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(G131), .B1(new_n427), .B2(new_n428), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n419), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n246), .B1(new_n431), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n260), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n413), .A2(new_n419), .A3(new_n423), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n227), .A2(KEYINPUT68), .A3(new_n228), .ZN(new_n448));
  AOI21_X1  g262(.A(KEYINPUT68), .B1(new_n227), .B2(new_n228), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n412), .B1(new_n443), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n426), .A2(new_n429), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n260), .B1(new_n440), .B2(new_n419), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT68), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n229), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n227), .A2(new_n228), .A3(KEYINPUT68), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(KEYINPUT28), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT26), .B(G101), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n298), .A2(G210), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n461), .B(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n463), .A2(new_n464), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n460), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n452), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT29), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n467), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n455), .A2(KEYINPUT30), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n430), .A2(new_n424), .B1(new_n439), .B2(new_n441), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n229), .B(new_n473), .C1(new_n474), .C2(KEYINPUT30), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n445), .B(new_n446), .C1(new_n448), .C2(new_n449), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n410), .B1(new_n471), .B2(new_n477), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n458), .B(new_n457), .C1(new_n453), .C2(new_n454), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT28), .ZN(new_n481));
  INV_X1    g295(.A(new_n460), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT29), .B1(new_n465), .B2(new_n466), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT73), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n460), .B1(new_n480), .B2(KEYINPUT28), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(KEYINPUT73), .A3(new_n484), .ZN(new_n489));
  AOI21_X1  g303(.A(G902), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n477), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT29), .B1(new_n452), .B2(new_n468), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT72), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n478), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(G472), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n451), .A2(new_n467), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n475), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT31), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n475), .A2(KEYINPUT31), .A3(new_n496), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n452), .A2(new_n482), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n499), .A2(new_n500), .B1(new_n501), .B2(new_n467), .ZN(new_n502));
  NOR2_X1   g316(.A1(G472), .A2(G902), .ZN(new_n503));
  XOR2_X1   g317(.A(new_n503), .B(KEYINPUT71), .Z(new_n504));
  OAI21_X1  g318(.A(KEYINPUT32), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n475), .A2(KEYINPUT31), .A3(new_n496), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT31), .B1(new_n475), .B2(new_n496), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n476), .B1(new_n474), .B2(new_n246), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n460), .B1(new_n508), .B2(new_n412), .ZN(new_n509));
  OAI22_X1  g323(.A1(new_n506), .A2(new_n507), .B1(new_n509), .B2(new_n472), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT32), .ZN(new_n511));
  INV_X1    g325(.A(new_n504), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n505), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n495), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G217), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n516), .B1(G234), .B2(new_n289), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT22), .B(G137), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n303), .A2(G221), .A3(G234), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G110), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT75), .ZN(new_n523));
  OAI211_X1 g337(.A(G119), .B(new_n267), .C1(new_n523), .C2(KEYINPUT23), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT23), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n525), .B1(new_n223), .B2(G128), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT75), .B1(new_n223), .B2(G128), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n522), .B(new_n524), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT76), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n267), .A2(G119), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n267), .A2(G119), .ZN(new_n531));
  OAI211_X1 g345(.A(KEYINPUT75), .B(new_n530), .C1(new_n531), .C2(new_n525), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT76), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n532), .A2(new_n533), .A3(new_n522), .A4(new_n524), .ZN(new_n534));
  INV_X1    g348(.A(new_n531), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n530), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n522), .A2(KEYINPUT24), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT24), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(G110), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT74), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n540), .B1(new_n537), .B2(new_n539), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n536), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n529), .A2(new_n534), .A3(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n325), .A2(new_n311), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT77), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n532), .A2(new_n524), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G110), .ZN(new_n549));
  INV_X1    g363(.A(new_n542), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n550), .A2(new_n530), .A3(new_n535), .A4(new_n551), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n549), .B(new_n552), .C1(new_n326), .C2(new_n325), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n546), .A2(new_n547), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n547), .B1(new_n546), .B2(new_n553), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n521), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n546), .A2(new_n553), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n520), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT25), .B1(new_n559), .B2(new_n289), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT25), .ZN(new_n561));
  AOI211_X1 g375(.A(new_n561), .B(G902), .C1(new_n556), .C2(new_n558), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n517), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n517), .A2(G902), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  OR2_X1    g381(.A1(new_n387), .A2(G902), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G221), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(KEYINPUT79), .ZN(new_n570));
  XNOR2_X1  g384(.A(G110), .B(G140), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n303), .A2(G227), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT81), .ZN(new_n575));
  INV_X1    g389(.A(new_n200), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n210), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n232), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n266), .A2(new_n268), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n575), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n233), .A2(new_n413), .A3(KEYINPUT81), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n579), .A2(new_n580), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n441), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT12), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n584), .A2(KEYINPUT12), .A3(new_n441), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT10), .ZN(new_n590));
  NOR4_X1   g404(.A1(new_n580), .A2(new_n206), .A3(new_n590), .A4(new_n232), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(new_n213), .B2(new_n444), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n581), .A2(new_n590), .A3(new_n582), .ZN(new_n593));
  INV_X1    g407(.A(new_n441), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n574), .B1(new_n589), .B2(new_n595), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n594), .B1(new_n592), .B2(new_n593), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n597), .A2(new_n598), .A3(new_n573), .ZN(new_n599));
  OAI21_X1  g413(.A(KEYINPUT82), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n584), .A2(KEYINPUT12), .A3(new_n441), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT12), .B1(new_n584), .B2(new_n441), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n595), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n573), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT82), .ZN(new_n605));
  INV_X1    g419(.A(new_n598), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(new_n595), .A3(new_n574), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n600), .A2(G469), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(G469), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n610), .A2(new_n289), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n595), .B(new_n574), .C1(new_n601), .C2(new_n602), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n573), .B1(new_n597), .B2(new_n598), .ZN(new_n613));
  AOI21_X1  g427(.A(G902), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n611), .B1(new_n614), .B2(new_n610), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n570), .B1(new_n609), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n409), .A2(new_n515), .A3(new_n567), .A4(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G101), .ZN(G3));
  INV_X1    g432(.A(G478), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n399), .A2(new_n406), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT97), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n400), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n398), .A2(KEYINPUT33), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(KEYINPUT33), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n404), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n623), .A2(new_n625), .A3(G478), .A4(new_n289), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n367), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n628), .A2(new_n297), .ZN(new_n629));
  INV_X1    g443(.A(G472), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n510), .B2(new_n289), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n502), .A2(new_n504), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n566), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n629), .A2(new_n633), .A3(new_n616), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT34), .B(G104), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  OAI21_X1  g450(.A(new_n344), .B1(new_n357), .B2(new_n358), .ZN(new_n637));
  INV_X1    g451(.A(new_n361), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n365), .A2(new_n361), .A3(new_n344), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AOI22_X1  g456(.A1(G475), .A2(new_n340), .B1(new_n397), .B2(new_n407), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n365), .A2(KEYINPUT98), .A3(new_n361), .A4(new_n344), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n297), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n646), .A2(new_n633), .A3(new_n616), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n647), .B(KEYINPUT99), .Z(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT35), .B(G107), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  INV_X1    g464(.A(KEYINPUT100), .ZN(new_n651));
  INV_X1    g465(.A(new_n517), .ZN(new_n652));
  INV_X1    g466(.A(new_n558), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n557), .A2(KEYINPUT77), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n546), .A2(new_n547), .A3(new_n553), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n653), .B1(new_n656), .B2(new_n521), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n561), .B1(new_n657), .B2(G902), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n559), .A2(KEYINPUT25), .A3(new_n289), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n652), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n656), .B1(KEYINPUT36), .B2(new_n521), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n521), .A2(KEYINPUT36), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n654), .A2(new_n655), .A3(new_n662), .ZN(new_n663));
  AOI211_X1 g477(.A(G902), .B(new_n517), .C1(new_n661), .C2(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n651), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n664), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n563), .A3(KEYINPUT100), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n631), .A2(new_n632), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n668), .A2(new_n409), .A3(new_n616), .A4(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  INV_X1    g486(.A(new_n187), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n292), .B1(new_n275), .B2(new_n290), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n294), .A2(new_n291), .A3(new_n295), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n495), .B2(new_n514), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n191), .B(KEYINPUT102), .ZN(new_n679));
  INV_X1    g493(.A(G900), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n190), .A2(new_n680), .A3(G902), .A4(G953), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n681), .B(KEYINPUT101), .Z(new_n682));
  NAND2_X1  g496(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n645), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n678), .A2(new_n668), .A3(new_n616), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n505), .A2(new_n513), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n475), .A2(new_n476), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n472), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n289), .B1(new_n480), .B2(new_n472), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n630), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n688), .B1(new_n689), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n694), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n514), .A2(KEYINPUT104), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n683), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n616), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT40), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n674), .A2(new_n675), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n658), .A2(new_n659), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n664), .B1(new_n707), .B2(new_n517), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n673), .B1(new_n397), .B2(new_n407), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(new_n367), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n711), .B1(KEYINPUT40), .B2(new_n701), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n713));
  OR3_X1    g527(.A1(new_n703), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n713), .B1(new_n703), .B2(new_n712), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n254), .ZN(G45));
  INV_X1    g531(.A(G475), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n339), .B2(new_n289), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n639), .B2(new_n359), .ZN(new_n720));
  INV_X1    g534(.A(new_n627), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n720), .A2(new_n721), .A3(new_n684), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n678), .A2(new_n668), .A3(new_n616), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G146), .ZN(G48));
  NAND2_X1  g538(.A1(new_n612), .A2(new_n613), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n289), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(G469), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n614), .A2(new_n610), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n569), .A3(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n515), .A2(new_n629), .A3(new_n567), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT41), .B(G113), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G15));
  NAND4_X1  g547(.A1(new_n515), .A2(new_n646), .A3(new_n730), .A4(new_n567), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G116), .ZN(G18));
  NAND2_X1  g549(.A1(new_n639), .A2(new_n359), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n397), .A2(new_n407), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n736), .A2(new_n195), .A3(new_n341), .A4(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n729), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n668), .A2(new_n515), .A3(new_n739), .A4(new_n676), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G119), .ZN(G21));
  OAI22_X1  g555(.A1(new_n506), .A2(new_n507), .B1(new_n472), .B2(new_n488), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n742), .A2(new_n512), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n566), .A2(new_n743), .A3(new_n631), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n367), .A2(new_n704), .A3(new_n709), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n744), .A2(new_n730), .A3(new_n745), .A4(new_n195), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT107), .B(G122), .Z(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G24));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n510), .A2(new_n289), .ZN(new_n750));
  AOI22_X1  g564(.A1(new_n750), .A2(G472), .B1(new_n512), .B2(new_n742), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n721), .B1(new_n736), .B2(new_n341), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n666), .A2(new_n563), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n751), .A2(new_n752), .A3(new_n753), .A4(new_n683), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n676), .A2(new_n569), .A3(new_n728), .A4(new_n727), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n749), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n755), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n708), .A2(new_n743), .A3(new_n631), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n757), .A2(new_n758), .A3(KEYINPUT108), .A4(new_n722), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G125), .ZN(G27));
  XOR2_X1   g575(.A(new_n611), .B(KEYINPUT109), .Z(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n614), .B2(new_n610), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n597), .B1(new_n588), .B2(new_n587), .ZN(new_n765));
  OAI211_X1 g579(.A(G469), .B(new_n607), .C1(new_n765), .C2(new_n574), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n604), .A2(KEYINPUT110), .A3(G469), .A4(new_n607), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n764), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n764), .A2(new_n768), .A3(KEYINPUT111), .A4(new_n769), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n566), .B1(new_n495), .B2(new_n514), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n674), .A2(new_n675), .A3(new_n187), .ZN(new_n776));
  INV_X1    g590(.A(new_n569), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n774), .A2(new_n775), .A3(new_n722), .A4(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT42), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n782));
  INV_X1    g596(.A(new_n778), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n783), .B1(new_n772), .B2(new_n773), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(KEYINPUT42), .A3(new_n775), .A4(new_n722), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n781), .A2(new_n782), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n782), .B1(new_n781), .B2(new_n785), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G131), .ZN(G33));
  NAND3_X1  g603(.A1(new_n784), .A2(new_n775), .A3(new_n685), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G134), .ZN(G36));
  NAND2_X1  g605(.A1(new_n720), .A2(new_n627), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT43), .Z(new_n793));
  INV_X1    g607(.A(new_n669), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(new_n794), .A3(new_n753), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT44), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n797), .A2(new_n798), .A3(new_n776), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT45), .B1(new_n600), .B2(new_n608), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n604), .A2(KEYINPUT45), .A3(new_n607), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(G469), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n762), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT46), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AOI22_X1  g619(.A1(new_n803), .A2(new_n804), .B1(new_n610), .B2(new_n614), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n777), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT113), .B1(new_n807), .B2(new_n700), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n807), .A2(KEYINPUT113), .A3(new_n700), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n799), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G137), .ZN(G39));
  XNOR2_X1  g625(.A(new_n807), .B(KEYINPUT47), .ZN(new_n812));
  INV_X1    g626(.A(new_n776), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n722), .A2(new_n566), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n515), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  NAND2_X1  g631(.A1(new_n727), .A2(new_n728), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n792), .B1(KEYINPUT49), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(KEYINPUT49), .B2(new_n818), .ZN(new_n820));
  INV_X1    g634(.A(new_n570), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n706), .A2(new_n567), .A3(new_n821), .A4(new_n187), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n698), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT114), .ZN(new_n824));
  INV_X1    g638(.A(new_n679), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n793), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n744), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n189), .B1(new_n827), .B2(new_n755), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n775), .A2(new_n826), .A3(new_n730), .A4(new_n813), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT48), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n730), .A2(new_n813), .ZN(new_n831));
  NOR4_X1   g645(.A1(new_n698), .A2(new_n566), .A3(new_n191), .A4(new_n831), .ZN(new_n832));
  AOI211_X1 g646(.A(new_n828), .B(new_n830), .C1(new_n752), .C2(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n827), .A2(new_n776), .ZN(new_n834));
  XOR2_X1   g648(.A(new_n834), .B(KEYINPUT117), .Z(new_n835));
  NOR2_X1   g649(.A1(new_n818), .A2(new_n821), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n835), .B1(new_n812), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT50), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n187), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n706), .A2(new_n730), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n827), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n838), .B2(new_n839), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n826), .A2(new_n730), .A3(new_n758), .A4(new_n813), .ZN(new_n844));
  OAI211_X1 g658(.A(KEYINPUT119), .B(KEYINPUT50), .C1(new_n827), .C2(new_n841), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n832), .A2(new_n720), .A3(new_n721), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n843), .A2(new_n844), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n837), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n836), .B(KEYINPUT118), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n812), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n847), .B1(new_n835), .B2(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n833), .B(new_n850), .C1(KEYINPUT51), .C2(new_n853), .ZN(new_n854));
  AND4_X1   g668(.A1(new_n617), .A2(new_n731), .A3(new_n734), .A4(new_n746), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n628), .B1(new_n367), .B2(new_n737), .ZN(new_n856));
  INV_X1    g670(.A(new_n297), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n633), .A3(new_n616), .A4(new_n857), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n670), .A2(new_n740), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n784), .A2(new_n722), .A3(new_n758), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n408), .A2(new_n719), .A3(new_n684), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n644), .A2(new_n813), .A3(new_n642), .A4(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(new_n668), .A3(new_n515), .A4(new_n616), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n790), .A2(new_n861), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT115), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT115), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n790), .A2(new_n861), .A3(new_n864), .A4(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n860), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT52), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n760), .A2(new_n686), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n708), .B2(new_n683), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n367), .A2(new_n569), .A3(new_n704), .A4(new_n709), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n708), .A2(new_n872), .A3(new_n683), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n875), .A2(new_n774), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT104), .B1(new_n514), .B2(new_n696), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n688), .B(new_n694), .C1(new_n505), .C2(new_n513), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n723), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n870), .B1(new_n871), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT72), .B1(new_n491), .B2(new_n492), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT73), .B1(new_n488), .B2(new_n484), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT28), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n885), .B1(new_n476), .B2(new_n479), .ZN(new_n886));
  NOR4_X1   g700(.A1(new_n886), .A2(new_n460), .A3(new_n486), .A4(new_n483), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n289), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n630), .B1(new_n889), .B2(new_n493), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n676), .B1(new_n689), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n609), .A2(new_n615), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n892), .A2(new_n821), .A3(new_n665), .A4(new_n667), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  AOI22_X1  g708(.A1(new_n894), .A2(new_n685), .B1(new_n756), .B2(new_n759), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n698), .A2(new_n774), .A3(new_n876), .A4(new_n875), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n895), .A2(KEYINPUT52), .A3(new_n723), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n882), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n869), .A2(new_n898), .A3(new_n788), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT53), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n869), .A2(new_n898), .A3(new_n788), .A4(KEYINPUT53), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT54), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n781), .A2(new_n785), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT53), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n882), .B2(new_n897), .ZN(new_n907));
  AOI22_X1  g721(.A1(new_n899), .A2(new_n900), .B1(new_n869), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT54), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n904), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n854), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(G952), .A2(G953), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n824), .B1(new_n912), .B2(new_n913), .ZN(G75));
  NOR2_X1   g728(.A1(new_n303), .A2(G952), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n908), .A2(new_n289), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT56), .B1(new_n917), .B2(G210), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n249), .A2(new_n251), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(new_n274), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT55), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n916), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n907), .A2(new_n869), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n901), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n924), .A2(KEYINPUT120), .A3(G902), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n908), .B2(new_n289), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n925), .A2(new_n927), .A3(new_n292), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT56), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n921), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT121), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT121), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n928), .A2(new_n933), .A3(new_n930), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n922), .B1(new_n932), .B2(new_n934), .ZN(G51));
  AOI221_X4 g749(.A(KEYINPUT54), .B1(new_n907), .B2(new_n869), .C1(new_n899), .C2(new_n900), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n909), .B1(new_n901), .B2(new_n923), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n762), .B(KEYINPUT57), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n725), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n800), .A2(new_n802), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n925), .A2(new_n927), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n915), .B1(new_n940), .B2(new_n942), .ZN(G54));
  AND2_X1   g757(.A1(KEYINPUT58), .A2(G475), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n925), .A2(new_n927), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n365), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n947), .A2(new_n948), .A3(new_n915), .ZN(G60));
  INV_X1    g763(.A(KEYINPUT122), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n623), .A2(new_n625), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(G478), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT59), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n952), .B1(new_n911), .B2(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n952), .A2(new_n954), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n936), .B2(new_n937), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n916), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n950), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n909), .B1(new_n901), .B2(new_n902), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n954), .B1(new_n936), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n951), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n962), .A2(KEYINPUT122), .A3(new_n916), .A4(new_n957), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n959), .A2(new_n963), .ZN(G63));
  NAND2_X1  g778(.A1(new_n661), .A2(new_n663), .ZN(new_n965));
  NAND2_X1  g779(.A1(G217), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT60), .Z(new_n967));
  NAND3_X1  g781(.A1(new_n924), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n924), .A2(new_n967), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n916), .B(new_n968), .C1(new_n969), .C2(new_n559), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(G66));
  OAI21_X1  g786(.A(G953), .B1(new_n192), .B2(new_n271), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(KEYINPUT123), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n860), .A2(new_n303), .ZN(new_n975));
  MUX2_X1   g789(.A(KEYINPUT123), .B(new_n974), .S(new_n975), .Z(new_n976));
  OAI21_X1  g790(.A(new_n919), .B1(G898), .B2(new_n303), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT124), .Z(new_n978));
  XOR2_X1   g792(.A(new_n976), .B(new_n978), .Z(G69));
  OAI211_X1 g793(.A(new_n775), .B(new_n745), .C1(new_n809), .C2(new_n808), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n810), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n895), .A2(new_n723), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n816), .A2(new_n788), .A3(new_n790), .A4(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n303), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(G900), .B2(new_n303), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n473), .B1(new_n474), .B2(KEYINPUT30), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n351), .B(KEYINPUT125), .Z(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT126), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT62), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n716), .B2(new_n982), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n983), .A2(KEYINPUT62), .A3(new_n715), .A4(new_n714), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n701), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n996), .A2(new_n775), .A3(new_n813), .A4(new_n856), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n810), .A2(new_n816), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n991), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n993), .A2(new_n994), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n816), .A2(new_n997), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n1000), .A2(KEYINPUT126), .A3(new_n810), .A4(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(G953), .B1(new_n999), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n990), .B1(new_n1003), .B2(new_n989), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n303), .B1(G227), .B2(G900), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1005), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n990), .B(new_n1007), .C1(new_n1003), .C2(new_n989), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1006), .A2(new_n1008), .ZN(G72));
  NAND4_X1  g823(.A1(new_n999), .A2(new_n859), .A3(new_n855), .A4(new_n1002), .ZN(new_n1010));
  XNOR2_X1  g824(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n630), .A2(new_n289), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1011), .B(new_n1012), .Z(new_n1013));
  AOI21_X1  g827(.A(new_n691), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  NOR3_X1   g828(.A1(new_n981), .A2(new_n984), .A3(new_n860), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1013), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR3_X1   g831(.A1(new_n1017), .A2(new_n472), .A3(new_n690), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1016), .B1(new_n491), .B2(new_n497), .ZN(new_n1019));
  AND2_X1   g833(.A1(new_n903), .A2(new_n1019), .ZN(new_n1020));
  NOR4_X1   g834(.A1(new_n1014), .A2(new_n1018), .A3(new_n915), .A4(new_n1020), .ZN(G57));
endmodule


