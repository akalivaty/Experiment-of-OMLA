//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 1 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n602, new_n603, new_n605,
    new_n606, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1220,
    new_n1221, new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT67), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  AOI21_X1  g042(.A(KEYINPUT68), .B1(new_n467), .B2(G101), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n465), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n462), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n472), .A2(new_n475), .ZN(G160));
  INV_X1    g051(.A(new_n464), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  XNOR2_X1  g058(.A(KEYINPUT3), .B(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n480), .B(new_n482), .C1(new_n483), .C2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n488), .A2(new_n490), .A3(G2104), .ZN(new_n491));
  AND2_X1   g066(.A1(G126), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n463), .B2(new_n464), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n463), .B2(new_n464), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n496), .B(new_n499), .C1(new_n464), .C2(new_n463), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n494), .B1(new_n498), .B2(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n504), .A2(new_n506), .B1(new_n503), .B2(G543), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n505), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(new_n512), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n507), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n510), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n513), .A2(G51), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n520), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n507), .A2(G89), .A3(new_n515), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(G168));
  NAND2_X1  g101(.A1(new_n507), .A2(G64), .ZN(new_n527));
  NAND2_X1  g102(.A1(G77), .A2(G543), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n509), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n507), .A2(G90), .A3(new_n515), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n513), .A2(G52), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT70), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  NOR3_X1   g109(.A1(new_n529), .A2(new_n532), .A3(KEYINPUT70), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  AOI22_X1  g112(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n509), .ZN(new_n539));
  INV_X1    g114(.A(G81), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n515), .A2(G543), .ZN(new_n541));
  XNOR2_X1  g116(.A(KEYINPUT71), .B(G43), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n516), .A2(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  INV_X1    g124(.A(new_n516), .ZN(new_n550));
  INV_X1    g125(.A(G53), .ZN(new_n551));
  OAI21_X1  g126(.A(KEYINPUT9), .B1(new_n541), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n513), .A2(new_n553), .A3(G53), .ZN(new_n554));
  AOI22_X1  g129(.A1(G91), .A2(new_n550), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n504), .A2(new_n506), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n503), .A2(G543), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n556), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(KEYINPUT72), .B1(new_n561), .B2(G651), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT72), .ZN(new_n564));
  NOR3_X1   g139(.A1(new_n563), .A2(new_n564), .A3(new_n509), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n555), .B1(new_n562), .B2(new_n565), .ZN(G299));
  INV_X1    g141(.A(G168), .ZN(G286));
  OAI221_X1 g142(.A(new_n514), .B1(new_n516), .B2(new_n517), .C1(new_n508), .C2(new_n509), .ZN(G303));
  OAI21_X1  g143(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n557), .A2(G87), .A3(new_n515), .A4(new_n558), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n513), .A2(G49), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  NAND2_X1  g147(.A1(new_n507), .A2(G61), .ZN(new_n573));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G651), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n507), .A2(G86), .A3(new_n515), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n513), .A2(G48), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n576), .A2(new_n579), .ZN(G305));
  AOI22_X1  g155(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n509), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n513), .A2(G47), .ZN(new_n583));
  INV_X1    g158(.A(G85), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n516), .B2(new_n584), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n582), .A2(new_n585), .ZN(G290));
  NAND3_X1  g161(.A1(new_n507), .A2(G92), .A3(new_n515), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G66), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n559), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(G54), .B2(new_n513), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(G868), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(G171), .B2(G868), .ZN(G321));
  XOR2_X1   g171(.A(G321), .B(KEYINPUT73), .Z(G284));
  NAND2_X1  g172(.A1(G286), .A2(G868), .ZN(new_n598));
  INV_X1    g173(.A(G299), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(G868), .ZN(G297));
  OAI21_X1  g175(.A(new_n598), .B1(new_n599), .B2(G868), .ZN(G280));
  AND2_X1   g176(.A1(new_n589), .A2(new_n593), .ZN(new_n602));
  XOR2_X1   g177(.A(KEYINPUT74), .B(G559), .Z(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(G860), .B2(new_n603), .ZN(G148));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G868), .B2(new_n544), .ZN(G323));
  XNOR2_X1  g182(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g183(.A1(new_n484), .A2(new_n467), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT12), .Z(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT13), .Z(new_n611));
  XOR2_X1   g186(.A(KEYINPUT75), .B(G2100), .Z(new_n612));
  OR2_X1    g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n463), .A2(new_n464), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n615), .A2(new_n462), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n616), .A2(G123), .B1(new_n479), .B2(G135), .ZN(new_n617));
  NOR3_X1   g192(.A1(new_n462), .A2(KEYINPUT76), .A3(G111), .ZN(new_n618));
  OAI21_X1  g193(.A(KEYINPUT76), .B1(new_n462), .B2(G111), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n619), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n617), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND3_X1  g197(.A1(new_n613), .A2(new_n614), .A3(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(G2427), .B(G2438), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2430), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n627), .A2(KEYINPUT14), .A3(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT77), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G1341), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G1348), .ZN(new_n633));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n635), .B(new_n636), .Z(new_n637));
  OR2_X1    g212(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(G14), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n639), .B1(new_n633), .B2(new_n637), .ZN(new_n640));
  AND2_X1   g215(.A1(new_n638), .A2(new_n640), .ZN(G401));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT78), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2072), .B(G2078), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2067), .B(G2678), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT18), .Z(new_n647));
  OR2_X1    g222(.A1(new_n643), .A2(new_n645), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n643), .A2(new_n645), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n644), .B(KEYINPUT17), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n644), .B(KEYINPUT79), .Z(new_n652));
  OAI211_X1 g227(.A(new_n647), .B(new_n651), .C1(new_n648), .C2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2096), .B(G2100), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT80), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n653), .B(new_n655), .ZN(G227));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT81), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1956), .B(G2474), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n659), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT20), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n659), .B1(new_n661), .B2(new_n663), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n661), .A2(new_n663), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n665), .B(new_n668), .C1(new_n658), .C2(new_n667), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT82), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(new_n675), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(G229));
  AOI22_X1  g253(.A1(new_n479), .A2(G141), .B1(G105), .B2(new_n467), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n616), .A2(G129), .ZN(new_n680));
  NAND3_X1  g255(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT26), .Z(new_n682));
  NAND3_X1  g257(.A1(new_n679), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(G29), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT90), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g262(.A(KEYINPUT90), .B1(G29), .B2(G32), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT27), .B(G1996), .Z(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g266(.A1(KEYINPUT24), .A2(G34), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n684), .B1(KEYINPUT24), .B2(G34), .ZN(new_n693));
  OAI22_X1  g268(.A1(G160), .A2(new_n684), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G5), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G171), .B2(new_n695), .ZN(new_n697));
  OAI221_X1 g272(.A(new_n691), .B1(G2084), .B2(new_n694), .C1(new_n697), .C2(G1961), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT91), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n695), .A2(G21), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G168), .B2(new_n695), .ZN(new_n701));
  INV_X1    g276(.A(G1966), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT30), .B(G28), .ZN(new_n704));
  OR2_X1    g279(.A1(KEYINPUT31), .A2(G11), .ZN(new_n705));
  NAND2_X1  g280(.A1(KEYINPUT31), .A2(G11), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n704), .A2(new_n684), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(new_n621), .B2(new_n684), .ZN(new_n708));
  OAI21_X1  g283(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n484), .A2(new_n492), .B1(new_n710), .B2(new_n490), .ZN(new_n711));
  INV_X1    g286(.A(new_n500), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n499), .B1(new_n484), .B2(new_n496), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n684), .A2(G27), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G2078), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n708), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n717), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n720), .A2(G2078), .B1(G2084), .B2(new_n694), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n703), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n684), .A2(G35), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G162), .B2(new_n684), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT29), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G2090), .ZN(new_n726));
  AOI211_X1 g301(.A(new_n722), .B(new_n726), .C1(G1961), .C2(new_n697), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n695), .A2(G20), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT92), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT23), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n599), .B2(new_n695), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT93), .B(G1956), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n695), .A2(G4), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n602), .B2(new_n695), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1348), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n695), .A2(G19), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n544), .B2(new_n695), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1341), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n684), .A2(G26), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT28), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n616), .A2(G128), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n479), .A2(G140), .ZN(new_n743));
  OR2_X1    g318(.A1(G104), .A2(G2105), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n744), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n741), .B1(new_n747), .B2(new_n684), .ZN(new_n748));
  INV_X1    g323(.A(G2067), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n689), .B2(new_n690), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n684), .A2(G33), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT25), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n479), .A2(G139), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n484), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n757), .A2(new_n462), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n752), .B1(new_n759), .B2(new_n684), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G2072), .ZN(new_n761));
  NOR4_X1   g336(.A1(new_n736), .A2(new_n739), .A3(new_n751), .A4(new_n761), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n699), .A2(new_n727), .A3(new_n733), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n695), .A2(G22), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G166), .B2(new_n695), .ZN(new_n765));
  INV_X1    g340(.A(G1971), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT88), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n695), .A2(G6), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n509), .B1(new_n573), .B2(new_n574), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n577), .A2(new_n578), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n771), .B1(new_n774), .B2(new_n695), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT32), .B(G1981), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT85), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n775), .B(new_n777), .Z(new_n778));
  NOR3_X1   g353(.A1(new_n769), .A2(new_n770), .A3(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(G74), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n509), .B1(new_n559), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n570), .A2(new_n571), .ZN(new_n782));
  OAI21_X1  g357(.A(KEYINPUT86), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT86), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n569), .A2(new_n784), .A3(new_n570), .A4(new_n571), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  MUX2_X1   g361(.A(G23), .B(new_n786), .S(G16), .Z(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT33), .B(G1976), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT87), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n779), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(KEYINPUT34), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n695), .A2(G24), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n582), .A2(new_n585), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n796), .B2(new_n695), .ZN(new_n797));
  INV_X1    g372(.A(G1986), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n799), .A2(KEYINPUT84), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(KEYINPUT84), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n616), .A2(G119), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n479), .A2(G131), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n462), .A2(G107), .ZN(new_n804));
  OAI21_X1  g379(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n802), .B(new_n803), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G25), .B(new_n806), .S(G29), .Z(new_n807));
  XOR2_X1   g382(.A(KEYINPUT35), .B(G1991), .Z(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT83), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n807), .B(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n800), .A2(KEYINPUT89), .A3(new_n801), .A4(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n793), .B2(KEYINPUT34), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n794), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(KEYINPUT36), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT36), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n794), .A2(new_n815), .A3(new_n812), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n763), .B1(new_n814), .B2(new_n816), .ZN(G311));
  NAND2_X1  g392(.A1(new_n814), .A2(new_n816), .ZN(new_n818));
  INV_X1    g393(.A(new_n763), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(G150));
  NAND2_X1  g395(.A1(new_n602), .A2(G559), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT94), .B(KEYINPUT38), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(G80), .A2(G543), .ZN(new_n824));
  INV_X1    g399(.A(G67), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n559), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(KEYINPUT95), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT95), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n828), .B(new_n824), .C1(new_n559), .C2(new_n825), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n827), .A2(G651), .A3(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT96), .B(G55), .Z(new_n831));
  AOI22_X1  g406(.A1(new_n550), .A2(G93), .B1(new_n513), .B2(new_n831), .ZN(new_n832));
  AND3_X1   g407(.A1(new_n830), .A2(new_n544), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n544), .B1(new_n830), .B2(new_n832), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n823), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT39), .ZN(new_n838));
  AOI21_X1  g413(.A(G860), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n838), .B2(new_n837), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT97), .Z(new_n841));
  NAND2_X1  g416(.A1(new_n830), .A2(new_n832), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G860), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT98), .B(KEYINPUT37), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n841), .A2(new_n845), .ZN(G145));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n806), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(new_n610), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n806), .B(KEYINPUT100), .ZN(new_n850));
  INV_X1    g425(.A(new_n610), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n616), .A2(G130), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n479), .A2(G142), .ZN(new_n855));
  OR2_X1    g430(.A1(G106), .A2(G2105), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n856), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n853), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n858), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n849), .A2(new_n852), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n498), .A2(new_n500), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n494), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n491), .A2(new_n493), .A3(KEYINPUT99), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n863), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n746), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n683), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n759), .ZN(new_n870));
  INV_X1    g445(.A(new_n683), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n868), .B(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n759), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n862), .A2(new_n870), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n621), .B(G160), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(G162), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n870), .A2(new_n874), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n882), .A2(new_n861), .A3(new_n859), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n883), .A2(new_n876), .A3(new_n875), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(new_n880), .A3(new_n875), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n887), .A2(KEYINPUT102), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(KEYINPUT102), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n885), .B(new_n886), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g466(.A(new_n835), .B(new_n605), .ZN(new_n892));
  NAND2_X1  g467(.A1(G299), .A2(new_n594), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n564), .B1(new_n563), .B2(new_n509), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n561), .A2(KEYINPUT72), .A3(G651), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n896), .A2(new_n555), .A3(new_n589), .A4(new_n593), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n893), .A2(KEYINPUT41), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT41), .B1(new_n893), .B2(new_n897), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n892), .A2(new_n901), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n893), .A2(new_n897), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n902), .B1(new_n903), .B2(new_n892), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n786), .A2(new_n774), .ZN(new_n906));
  AOI21_X1  g481(.A(G305), .B1(new_n783), .B2(new_n785), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(G290), .A2(G166), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n796), .A2(G303), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n910), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n906), .B2(new_n907), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n905), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n916), .B1(new_n905), .B2(new_n917), .ZN(new_n919));
  OAI21_X1  g494(.A(G868), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G868), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n842), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(G295));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n922), .ZN(G331));
  AND3_X1   g499(.A1(new_n912), .A2(new_n914), .A3(KEYINPUT104), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT104), .B1(new_n912), .B2(new_n914), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(G286), .B1(new_n534), .B2(new_n535), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n527), .A2(new_n528), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(G651), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n530), .A2(new_n531), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT70), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n934), .A2(new_n533), .A3(G168), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n929), .B(new_n935), .C1(new_n833), .C2(new_n834), .ZN(new_n936));
  INV_X1    g511(.A(new_n544), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n842), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n830), .A2(new_n544), .A3(new_n832), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n934), .A2(new_n533), .A3(G168), .ZN(new_n940));
  AOI21_X1  g515(.A(G168), .B1(new_n934), .B2(new_n533), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n938), .B(new_n939), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n936), .A2(new_n942), .A3(new_n903), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(KEYINPUT103), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n929), .A2(new_n935), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT103), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n835), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n947), .A3(new_n936), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n900), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n943), .B1(new_n949), .B2(KEYINPUT106), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT106), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n951), .A3(new_n900), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n928), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n944), .A2(new_n947), .A3(new_n903), .A4(new_n936), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n936), .A2(new_n942), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n900), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(new_n956), .A3(new_n915), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT105), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n954), .A2(new_n956), .A3(new_n959), .A4(new_n915), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n958), .A2(new_n886), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n953), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n954), .A2(new_n956), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n927), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n958), .A2(new_n965), .A3(new_n886), .A4(new_n960), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n966), .A2(new_n962), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT44), .B1(new_n963), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n953), .A2(new_n961), .A3(KEYINPUT43), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n968), .A2(new_n972), .ZN(G397));
  INV_X1    g548(.A(G1384), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n867), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n473), .A2(new_n474), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(G2105), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n467), .A2(KEYINPUT68), .A3(G101), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n469), .A2(new_n470), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n979), .A2(G40), .A3(new_n465), .A4(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n977), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1996), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(new_n683), .ZN(new_n987));
  XOR2_X1   g562(.A(new_n987), .B(KEYINPUT107), .Z(new_n988));
  XNOR2_X1  g563(.A(new_n746), .B(new_n749), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT108), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n871), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n985), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n991), .A2(new_n992), .A3(new_n984), .ZN(new_n993));
  INV_X1    g568(.A(new_n808), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n806), .A2(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n806), .A2(new_n994), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n984), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(G290), .A2(G1986), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n796), .A2(new_n798), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n984), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n988), .A2(new_n993), .A3(new_n997), .A4(new_n1000), .ZN(new_n1001));
  XOR2_X1   g576(.A(new_n1001), .B(KEYINPUT109), .Z(new_n1002));
  INV_X1    g577(.A(KEYINPUT49), .ZN(new_n1003));
  INV_X1    g578(.A(G1981), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n576), .B2(new_n579), .ZN(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT115), .B(G1981), .Z(new_n1006));
  NOR3_X1   g581(.A1(new_n772), .A2(new_n773), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1003), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G8), .ZN(new_n1009));
  AOI22_X1  g584(.A1(KEYINPUT99), .A2(new_n711), .B1(new_n498), .B2(new_n500), .ZN(new_n1010));
  AOI21_X1  g585(.A(G1384), .B1(new_n1010), .B2(new_n865), .ZN(new_n1011));
  INV_X1    g586(.A(G40), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n472), .A2(new_n475), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1009), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1006), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n576), .A2(new_n579), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(G1981), .B1(new_n772), .B2(new_n773), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(KEYINPUT49), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1008), .A2(new_n1014), .A3(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n783), .A2(G1976), .A3(new_n785), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n783), .A2(KEYINPUT112), .A3(G1976), .A4(new_n785), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n1014), .A3(new_n1023), .ZN(new_n1024));
  XOR2_X1   g599(.A(KEYINPUT113), .B(G1976), .Z(new_n1025));
  NAND2_X1  g600(.A1(G288), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(KEYINPUT114), .A3(new_n1027), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1019), .B1(new_n1024), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n867), .A2(new_n1013), .A3(new_n974), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n1023), .A2(G8), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1027), .B1(new_n1035), .B2(new_n1022), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT118), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1035), .A2(new_n1022), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1024), .A2(KEYINPUT52), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .A4(new_n1019), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1037), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1043));
  OAI211_X1 g618(.A(KEYINPUT55), .B(G8), .C1(new_n510), .C2(new_n518), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT110), .ZN(new_n1047));
  AOI21_X1  g622(.A(G1384), .B1(new_n863), .B2(new_n711), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1013), .B1(new_n1048), .B2(KEYINPUT45), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n976), .A2(G1384), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1051), .B1(new_n1010), .B2(new_n865), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1047), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n976), .B1(G164), .B2(G1384), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n866), .B1(new_n712), .B2(new_n713), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n711), .A2(KEYINPUT99), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1050), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1054), .A2(new_n1057), .A3(KEYINPUT110), .A4(new_n1013), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1053), .A2(new_n766), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n867), .A2(new_n1060), .A3(new_n974), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT111), .B(G2090), .Z(new_n1063));
  NAND4_X1  g638(.A1(new_n1061), .A2(new_n1013), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  AOI211_X1 g639(.A(new_n1009), .B(new_n1046), .C1(new_n1059), .C2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1046), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n714), .A2(new_n1060), .A3(new_n974), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n1013), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1060), .B1(new_n867), .B2(new_n974), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n1063), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1059), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1066), .B1(new_n1072), .B2(G8), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1065), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1042), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT126), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1042), .A2(new_n1074), .A3(KEYINPUT126), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT45), .B1(new_n867), .B2(new_n974), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1013), .B1(G164), .B2(new_n1051), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n718), .A2(KEYINPUT53), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1061), .A2(new_n1013), .A3(new_n1062), .ZN(new_n1085));
  INV_X1    g660(.A(G1961), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1082), .A2(new_n1084), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(G2078), .B1(new_n1053), .B2(new_n1058), .ZN(new_n1088));
  OAI211_X1 g663(.A(G301), .B(new_n1087), .C1(new_n1088), .C2(KEYINPUT53), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n472), .A2(KEYINPUT125), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n979), .A2(G40), .A3(new_n1084), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n472), .A2(KEYINPUT125), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n977), .A2(new_n1094), .A3(new_n1057), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1090), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n714), .A2(new_n974), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n983), .B1(new_n1097), .B2(new_n976), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT110), .B1(new_n1098), .B2(new_n1057), .ZN(new_n1099));
  AND4_X1   g674(.A1(KEYINPUT110), .A2(new_n1054), .A3(new_n1057), .A4(new_n1013), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n718), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1096), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(KEYINPUT54), .B(new_n1089), .C1(new_n1103), .C2(G301), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT127), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1088), .A2(KEYINPUT53), .ZN(new_n1107));
  OAI21_X1  g682(.A(G171), .B1(new_n1107), .B2(new_n1096), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1108), .A2(KEYINPUT127), .A3(KEYINPUT54), .A4(new_n1089), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1087), .ZN(new_n1111));
  OAI21_X1  g686(.A(G171), .B1(new_n1107), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1096), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1113), .B(G301), .C1(KEYINPUT53), .C2(new_n1088), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n702), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(G2084), .B2(new_n1085), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1118), .A2(G286), .ZN(new_n1119));
  OAI21_X1  g694(.A(G8), .B1(new_n1118), .B2(G286), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT51), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1120), .A2(KEYINPUT51), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1115), .A2(new_n1116), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n1124));
  NAND2_X1  g699(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1125));
  INV_X1    g700(.A(G1956), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n896), .A2(new_n1128), .A3(new_n555), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT56), .B(G2072), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1098), .A2(new_n1057), .A3(new_n1130), .ZN(new_n1131));
  AND4_X1   g706(.A1(new_n1125), .A2(new_n1127), .A3(new_n1129), .A4(new_n1131), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1127), .A2(new_n1131), .B1(new_n1125), .B2(new_n1129), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1124), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1137));
  XOR2_X1   g712(.A(new_n1137), .B(KEYINPUT123), .Z(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT121), .B(G1996), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1054), .A2(new_n1057), .A3(new_n1013), .A4(new_n1140), .ZN(new_n1141));
  XOR2_X1   g716(.A(KEYINPUT58), .B(G1341), .Z(new_n1142));
  NAND2_X1  g717(.A1(new_n1034), .A2(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1136), .B(new_n1139), .C1(new_n1144), .C2(new_n937), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n937), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1138), .B1(new_n1146), .B2(new_n1135), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1125), .A2(new_n1129), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1127), .A2(new_n1125), .A3(new_n1131), .A4(new_n1129), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1151), .A2(KEYINPUT61), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1134), .A2(new_n1148), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(G1348), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1085), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(KEYINPUT120), .B1(new_n1034), .B2(G2067), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT120), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1011), .A2(new_n1158), .A3(new_n749), .A4(new_n1013), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1156), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT60), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1156), .A2(KEYINPUT60), .A3(new_n1157), .A4(new_n1159), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1163), .A2(KEYINPUT124), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1163), .A2(KEYINPUT124), .A3(new_n594), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n594), .B1(new_n1163), .B2(KEYINPUT124), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1154), .B1(new_n1162), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1152), .A2(new_n1160), .A3(new_n602), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1151), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1110), .B(new_n1123), .C1(new_n1168), .C2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1122), .A2(new_n1121), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1112), .B1(new_n1172), .B2(KEYINPUT62), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1173), .B1(KEYINPUT62), .B2(new_n1172), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1079), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n1118), .A2(G8), .A3(G168), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1042), .A2(new_n1074), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT63), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT116), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT116), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1038), .A2(new_n1039), .A3(new_n1181), .A4(new_n1019), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1009), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1184));
  OR2_X1    g759(.A1(new_n1184), .A2(new_n1066), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1118), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1186), .B1(new_n1066), .B2(new_n1184), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1183), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(KEYINPUT119), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT119), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1183), .A2(new_n1190), .A3(new_n1185), .A4(new_n1187), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1179), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1014), .ZN(new_n1193));
  NOR2_X1   g768(.A1(G288), .A2(G1976), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1019), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1193), .B1(new_n1195), .B2(new_n1016), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1196), .B1(new_n1183), .B2(new_n1065), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT117), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1184), .A2(new_n1066), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1200), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1201));
  OAI21_X1  g776(.A(KEYINPUT117), .B1(new_n1201), .B2(new_n1196), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1192), .A2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1002), .B1(new_n1175), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n991), .A2(new_n984), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n986), .B(KEYINPUT46), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(KEYINPUT47), .ZN(new_n1209));
  AND2_X1   g784(.A1(new_n988), .A2(new_n993), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1210), .A2(new_n997), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n984), .A2(new_n998), .ZN(new_n1212));
  XOR2_X1   g787(.A(new_n1212), .B(KEYINPUT48), .Z(new_n1213));
  OAI21_X1  g788(.A(new_n1209), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1210), .A2(new_n995), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1215), .B1(G2067), .B2(new_n746), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1214), .B1(new_n984), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1205), .A2(new_n1217), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g793(.A1(G227), .A2(new_n460), .ZN(new_n1220));
  NAND3_X1  g794(.A1(new_n676), .A2(new_n1220), .A3(new_n677), .ZN(new_n1221));
  AOI21_X1  g795(.A(new_n1221), .B1(new_n638), .B2(new_n640), .ZN(new_n1222));
  OAI211_X1 g796(.A(new_n890), .B(new_n1222), .C1(new_n970), .C2(new_n971), .ZN(G225));
  INV_X1    g797(.A(G225), .ZN(G308));
endmodule


