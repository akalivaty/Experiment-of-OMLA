//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n571, new_n572,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n583, new_n584, new_n585, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1214, new_n1215,
    new_n1216;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT65), .Z(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  OR2_X1    g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(G137), .A3(new_n463), .ZN(new_n464));
  AND3_X1   g039(.A1(new_n463), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT68), .B1(new_n463), .B2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(G101), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n469), .B1(new_n460), .B2(new_n461), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  AND3_X1   g046(.A1(KEYINPUT67), .A2(G113), .A3(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(KEYINPUT67), .B1(G113), .B2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n468), .B1(G2105), .B2(new_n476), .ZN(G160));
  AOI21_X1  g052(.A(new_n463), .B1(new_n460), .B2(new_n461), .ZN(new_n478));
  OR2_X1    g053(.A1(new_n478), .A2(KEYINPUT69), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(KEYINPUT69), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G112), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  AND2_X1   g061(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n487));
  NOR2_X1   g062(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n486), .B1(new_n490), .B2(G136), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n483), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  OAI211_X1 g068(.A(G126), .B(G2105), .C1(new_n487), .C2(new_n488), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n495), .A2(new_n497), .A3(G2104), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT70), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n494), .A2(new_n501), .A3(new_n498), .ZN(new_n502));
  XOR2_X1   g077(.A(KEYINPUT71), .B(KEYINPUT4), .Z(new_n503));
  NAND2_X1  g078(.A1(new_n463), .A2(G138), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n489), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G138), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(G2105), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT4), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n507), .B(new_n509), .C1(new_n488), .C2(new_n487), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n500), .A2(new_n502), .B1(new_n505), .B2(new_n510), .ZN(G164));
  OR2_X1    g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(new_n516), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  INV_X1    g098(.A(new_n520), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  OAI21_X1  g100(.A(G543), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G50), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n522), .A2(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n517), .A2(new_n528), .ZN(G166));
  NAND3_X1  g104(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G543), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n533), .B1(new_n519), .B2(new_n520), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT72), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G51), .ZN(new_n537));
  OAI211_X1 g112(.A(KEYINPUT73), .B(new_n530), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT73), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n537), .B1(new_n532), .B2(new_n535), .ZN(new_n540));
  INV_X1    g115(.A(new_n530), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n514), .A2(new_n521), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(KEYINPUT7), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n544), .A2(KEYINPUT7), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n543), .A2(G89), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n538), .A2(new_n542), .A3(new_n547), .ZN(G286));
  INV_X1    g123(.A(G286), .ZN(G168));
  XOR2_X1   g124(.A(KEYINPUT74), .B(G52), .Z(new_n550));
  NOR2_X1   g125(.A1(new_n536), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G90), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n552), .A2(new_n516), .B1(new_n522), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(G171));
  AND2_X1   g130(.A1(new_n512), .A2(new_n513), .ZN(new_n556));
  INV_X1    g131(.A(G56), .ZN(new_n557));
  INV_X1    g132(.A(G68), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n556), .A2(new_n557), .B1(new_n558), .B2(new_n533), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT75), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n561));
  OAI221_X1 g136(.A(new_n561), .B1(new_n558), .B2(new_n533), .C1(new_n556), .C2(new_n557), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n560), .A2(G651), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n532), .A2(new_n535), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n564), .A2(G43), .B1(G81), .B2(new_n543), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(G860), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  XOR2_X1   g143(.A(new_n568), .B(KEYINPUT76), .Z(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND4_X1  g147(.A1(G319), .A2(G483), .A3(G661), .A4(new_n572), .ZN(G188));
  NAND2_X1  g148(.A1(new_n534), .A2(G53), .ZN(new_n574));
  NAND2_X1  g149(.A1(KEYINPUT77), .A2(KEYINPUT9), .ZN(new_n575));
  XOR2_X1   g150(.A(new_n574), .B(new_n575), .Z(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n556), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(G651), .B1(new_n543), .B2(G91), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(G299));
  INV_X1    g156(.A(G171), .ZN(G301));
  NAND2_X1  g157(.A1(G166), .A2(KEYINPUT78), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n584), .B1(new_n517), .B2(new_n528), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n583), .A2(new_n585), .ZN(G303));
  NAND2_X1  g161(.A1(new_n543), .A2(G87), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n534), .A2(G49), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G288));
  NAND2_X1  g165(.A1(new_n543), .A2(G86), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT79), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(new_n512), .B2(new_n513), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n534), .A2(G48), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n591), .A2(new_n596), .A3(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n556), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(new_n543), .B2(G85), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n564), .A2(G47), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  AND3_X1   g180(.A1(new_n514), .A2(new_n521), .A3(G92), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT10), .Z(new_n607));
  AOI22_X1  g182(.A1(new_n514), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n516), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n564), .A2(G54), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n605), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n605), .B1(new_n613), .B2(G868), .ZN(G321));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(G299), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G168), .B2(new_n616), .ZN(G297));
  OAI21_X1  g193(.A(new_n617), .B1(G168), .B2(new_n616), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n613), .A2(new_n620), .ZN(new_n622));
  MUX2_X1   g197(.A(new_n566), .B(new_n622), .S(G868), .Z(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n482), .A2(G123), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT80), .Z(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT81), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(G111), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n627), .A2(new_n628), .B1(new_n630), .B2(G2105), .ZN(new_n631));
  AOI22_X1  g206(.A1(new_n490), .A2(G135), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(G2096), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(G2096), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n465), .A2(new_n466), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(new_n462), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT13), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2100), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n634), .A2(new_n635), .A3(new_n640), .ZN(G156));
  INV_X1    g216(.A(G14), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(KEYINPUT14), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n648), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n642), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT82), .ZN(new_n656));
  INV_X1    g231(.A(new_n653), .ZN(new_n657));
  INV_X1    g232(.A(new_n654), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NOR3_X1   g234(.A1(new_n653), .A2(KEYINPUT82), .A3(new_n654), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT83), .Z(G401));
  XNOR2_X1  g237(.A(KEYINPUT86), .B(G2100), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT84), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(G2072), .A2(G2078), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n442), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n669), .B(KEYINPUT17), .Z(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(new_n666), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2084), .B(G2090), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT85), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n667), .A2(new_n669), .A3(new_n673), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT18), .ZN(new_n677));
  OR3_X1    g252(.A1(new_n671), .A2(new_n666), .A3(new_n673), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n675), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n679), .A2(G2096), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(G2096), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n664), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n679), .A2(G2096), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n679), .A2(G2096), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n683), .A2(new_n684), .A3(new_n663), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(G227));
  XOR2_X1   g261(.A(G1991), .B(G1996), .Z(new_n687));
  XOR2_X1   g262(.A(G1971), .B(G1976), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n690), .A2(new_n691), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  MUX2_X1   g272(.A(new_n697), .B(new_n696), .S(new_n689), .Z(new_n698));
  OR3_X1    g273(.A1(new_n695), .A2(new_n698), .A3(KEYINPUT87), .ZN(new_n699));
  OAI21_X1  g274(.A(KEYINPUT87), .B1(new_n695), .B2(new_n698), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n701), .B1(new_n699), .B2(new_n700), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n687), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n704), .ZN(new_n706));
  INV_X1    g281(.A(new_n687), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n706), .A2(new_n707), .A3(new_n702), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1981), .B(G1986), .ZN(new_n709));
  AND3_X1   g284(.A1(new_n705), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n705), .B2(new_n708), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(G229));
  NOR2_X1   g287(.A1(G6), .A2(G16), .ZN(new_n713));
  AND3_X1   g288(.A1(new_n591), .A2(new_n596), .A3(new_n597), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(G16), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT32), .ZN(new_n716));
  INV_X1    g291(.A(G1981), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G23), .ZN(new_n720));
  INV_X1    g295(.A(G288), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n719), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT33), .B(G1976), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n719), .A2(G22), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G166), .B2(new_n719), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT89), .Z(new_n727));
  AOI21_X1  g302(.A(new_n724), .B1(new_n727), .B2(G1971), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n718), .B(new_n728), .C1(G1971), .C2(new_n727), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT88), .B(KEYINPUT34), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G25), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n482), .A2(G119), .ZN(new_n735));
  OAI21_X1  g310(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n736));
  INV_X1    g311(.A(G107), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(G2105), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n490), .B2(G131), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n734), .B1(new_n740), .B2(new_n733), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT35), .B(G1991), .Z(new_n742));
  XOR2_X1   g317(.A(new_n741), .B(new_n742), .Z(new_n743));
  MUX2_X1   g318(.A(G24), .B(G290), .S(G16), .Z(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G1986), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT90), .B(KEYINPUT36), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n731), .A2(new_n732), .A3(new_n746), .A4(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT91), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n731), .A2(new_n732), .A3(new_n746), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n749), .A2(new_n750), .B1(KEYINPUT36), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n748), .A2(KEYINPUT91), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n733), .A2(G35), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G162), .B2(new_n733), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT29), .B(G2090), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT24), .ZN(new_n759));
  INV_X1    g334(.A(G34), .ZN(new_n760));
  AOI21_X1  g335(.A(G29), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n759), .B2(new_n760), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G160), .B2(new_n733), .ZN(new_n763));
  INV_X1    g338(.A(G2084), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(G29), .A2(G33), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n462), .A2(G127), .ZN(new_n767));
  AND2_X1   g342(.A1(G115), .A2(G2104), .ZN(new_n768));
  OAI21_X1  g343(.A(G2105), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT25), .ZN(new_n770));
  NAND2_X1  g345(.A1(G103), .A2(G2104), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(G2105), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n463), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n490), .A2(G139), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n766), .B1(new_n776), .B2(G29), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT93), .B(G2072), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n758), .A2(new_n765), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n733), .A2(G32), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n482), .A2(G129), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT94), .B(KEYINPUT26), .Z(new_n783));
  NAND3_X1  g358(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n636), .A2(G105), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n490), .A2(G141), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n782), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n781), .B1(new_n789), .B2(new_n733), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT27), .B(G1996), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n790), .B(new_n791), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n719), .A2(G20), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT23), .Z(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G299), .B2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1956), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n733), .A2(G27), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G164), .B2(new_n733), .ZN(new_n798));
  INV_X1    g373(.A(G2078), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n719), .A2(G5), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G171), .B2(new_n719), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1961), .ZN(new_n804));
  NOR4_X1   g379(.A1(new_n780), .A2(new_n792), .A3(new_n801), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n719), .A2(G4), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n613), .B2(new_n719), .ZN(new_n807));
  INV_X1    g382(.A(G1348), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  MUX2_X1   g384(.A(G19), .B(new_n566), .S(G16), .Z(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(G1341), .Z(new_n811));
  NAND2_X1  g386(.A1(new_n490), .A2(G140), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT92), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n479), .A2(G128), .A3(new_n480), .ZN(new_n815));
  OR2_X1    g390(.A1(G104), .A2(G2105), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n816), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n814), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(G29), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n733), .A2(G26), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT28), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(G2067), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n805), .A2(new_n809), .A3(new_n811), .A4(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT31), .B(G11), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT30), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G28), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT95), .Z(new_n829));
  OAI211_X1 g404(.A(new_n829), .B(new_n733), .C1(new_n827), .C2(G28), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n826), .B(new_n830), .C1(new_n633), .C2(new_n733), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT96), .ZN(new_n832));
  NOR2_X1   g407(.A1(G168), .A2(new_n719), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(new_n719), .B2(G21), .ZN(new_n834));
  INV_X1    g409(.A(G1966), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n832), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  OR3_X1    g413(.A1(new_n825), .A2(KEYINPUT97), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(KEYINPUT97), .B1(new_n825), .B2(new_n838), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n754), .A2(new_n841), .ZN(G311));
  NAND2_X1  g417(.A1(new_n754), .A2(new_n841), .ZN(G150));
  NAND2_X1  g418(.A1(new_n564), .A2(G55), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT98), .B(G93), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n543), .A2(new_n845), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n844), .B(new_n846), .C1(new_n516), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G860), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT100), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT37), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n613), .A2(G559), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT38), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n566), .A2(new_n848), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n566), .A2(new_n848), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n853), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT99), .Z(new_n860));
  OAI21_X1  g435(.A(new_n567), .B1(new_n857), .B2(new_n858), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n851), .B1(new_n860), .B2(new_n861), .ZN(G145));
  XOR2_X1   g437(.A(new_n492), .B(G160), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n633), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT101), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  INV_X1    g441(.A(G118), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n866), .B1(new_n867), .B2(G2105), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(new_n490), .B2(G142), .ZN(new_n869));
  INV_X1    g444(.A(G130), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n638), .B(new_n869), .C1(new_n870), .C2(new_n481), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n637), .B(KEYINPUT12), .Z(new_n872));
  OAI21_X1  g447(.A(new_n869), .B1(new_n481), .B2(new_n870), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n871), .A2(new_n740), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n740), .B1(new_n871), .B2(new_n874), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n865), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n871), .A2(new_n874), .ZN(new_n878));
  INV_X1    g453(.A(new_n740), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n871), .A2(new_n740), .A3(new_n874), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n880), .A2(KEYINPUT101), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n818), .A2(new_n775), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n504), .B1(new_n460), .B2(new_n461), .ZN(new_n885));
  XNOR2_X1  g460(.A(KEYINPUT71), .B(KEYINPUT4), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n510), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n463), .A2(G114), .ZN(new_n888));
  OAI21_X1  g463(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(new_n478), .B2(G126), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n776), .A2(new_n814), .A3(new_n815), .A4(new_n817), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n884), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n892), .B1(new_n884), .B2(new_n893), .ZN(new_n896));
  INV_X1    g471(.A(new_n789), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n884), .A2(new_n893), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n499), .B1(new_n505), .B2(new_n510), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n789), .B1(new_n901), .B2(new_n894), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n883), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT102), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n897), .B1(new_n895), .B2(new_n896), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(new_n789), .A3(new_n894), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n908), .A3(new_n883), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n864), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  OR3_X1    g485(.A1(new_n898), .A2(new_n902), .A3(KEYINPUT103), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n907), .A2(KEYINPUT103), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n911), .A2(new_n881), .A3(new_n880), .A4(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(G37), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n909), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n908), .B1(new_n907), .B2(new_n883), .ZN(new_n916));
  OAI22_X1  g491(.A1(new_n915), .A2(new_n916), .B1(new_n907), .B2(new_n883), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n864), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g495(.A1(new_n848), .A2(new_n616), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n714), .B(G166), .ZN(new_n922));
  XNOR2_X1  g497(.A(G290), .B(G288), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(new_n924), .B2(new_n923), .ZN(new_n926));
  INV_X1    g501(.A(new_n923), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n927), .A2(KEYINPUT105), .A3(new_n922), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(KEYINPUT106), .B2(KEYINPUT42), .ZN(new_n931));
  NAND2_X1  g506(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n931), .B(new_n932), .Z(new_n933));
  XOR2_X1   g508(.A(new_n856), .B(KEYINPUT104), .Z(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(new_n622), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n612), .A2(G299), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n610), .A2(new_n576), .A3(new_n580), .A4(new_n611), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n936), .A2(KEYINPUT41), .A3(new_n937), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT41), .B1(new_n936), .B2(new_n937), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n939), .B1(new_n935), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n933), .B(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n921), .B1(new_n944), .B2(new_n616), .ZN(G295));
  OAI21_X1  g520(.A(new_n921), .B1(new_n944), .B2(new_n616), .ZN(G331));
  NOR2_X1   g521(.A1(G286), .A2(KEYINPUT107), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n856), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(G171), .B1(G286), .B2(KEYINPUT107), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n854), .B(new_n855), .C1(KEYINPUT107), .C2(G286), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n949), .B1(new_n948), .B2(new_n950), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n942), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n948), .A2(new_n950), .ZN(new_n955));
  INV_X1    g530(.A(new_n949), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n938), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(new_n958), .A3(new_n951), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n954), .A2(new_n959), .A3(KEYINPUT108), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n957), .A2(new_n961), .A3(new_n958), .A4(new_n951), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n929), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n964));
  INV_X1    g539(.A(G37), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n954), .A2(new_n959), .A3(new_n930), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n963), .A2(new_n964), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n965), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n930), .B1(new_n954), .B2(new_n959), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT43), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n964), .B1(new_n968), .B2(new_n969), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n972), .B1(new_n973), .B2(new_n964), .ZN(new_n974));
  MUX2_X1   g549(.A(new_n971), .B(new_n974), .S(KEYINPUT44), .Z(G397));
  INV_X1    g550(.A(KEYINPUT124), .ZN(new_n976));
  AOI21_X1  g551(.A(G1384), .B1(new_n887), .B2(new_n891), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT45), .ZN(new_n978));
  OAI21_X1  g553(.A(G2105), .B1(new_n470), .B2(new_n474), .ZN(new_n979));
  XOR2_X1   g554(.A(KEYINPUT109), .B(G40), .Z(new_n980));
  AND4_X1   g555(.A1(new_n979), .A2(new_n467), .A3(new_n464), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n494), .A2(new_n501), .A3(new_n498), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n501), .B1(new_n494), .B2(new_n498), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n887), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1384), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT45), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n982), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n799), .ZN(new_n989));
  XNOR2_X1  g564(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n985), .A2(KEYINPUT45), .A3(new_n986), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(new_n900), .B2(G1384), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n992), .A2(new_n799), .A3(new_n994), .A4(new_n981), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT119), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n979), .A2(new_n467), .A3(new_n464), .A4(new_n980), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n892), .A2(new_n986), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n998), .B1(new_n999), .B2(new_n993), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n1000), .A2(KEYINPUT119), .A3(new_n799), .A4(new_n992), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(KEYINPUT53), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT120), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n998), .B1(new_n977), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1961), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n1002), .A2(new_n1003), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1003), .B1(new_n1002), .B2(new_n1009), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n991), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n981), .B1(new_n999), .B2(KEYINPUT50), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1005), .B1(new_n985), .B2(new_n986), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1014), .A2(new_n1015), .A3(G2090), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n993), .B1(G164), .B2(G1384), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n998), .B1(new_n977), .B2(KEYINPUT45), .ZN(new_n1018));
  AOI21_X1  g593(.A(G1971), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1013), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n583), .A2(G8), .A3(new_n585), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(KEYINPUT111), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n583), .A2(G8), .A3(new_n585), .A4(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1971), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n982), .B2(new_n987), .ZN(new_n1031));
  INV_X1    g606(.A(G2090), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1004), .A2(new_n1032), .A3(new_n1006), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n1033), .A3(KEYINPUT110), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1020), .A2(G8), .A3(new_n1029), .A4(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(G305), .A2(G1981), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n543), .A2(G86), .B1(G48), .B2(new_n534), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(new_n717), .A3(new_n596), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1036), .A2(KEYINPUT49), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G8), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1040), .B1(new_n981), .B2(new_n977), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT49), .ZN(new_n1043));
  NOR2_X1   g618(.A1(G305), .A2(G1981), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n717), .B1(new_n1037), .B2(new_n596), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT112), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1048), .B(new_n1043), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1042), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1041), .ZN(new_n1051));
  INV_X1    g626(.A(G1976), .ZN(new_n1052));
  NOR2_X1   g627(.A1(G288), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT52), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT52), .B1(G288), .B2(new_n1052), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1041), .B(new_n1055), .C1(new_n1052), .C2(G288), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1050), .A2(new_n1057), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1035), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1005), .B1(new_n892), .B2(new_n986), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(new_n1061), .B2(new_n998), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n985), .A2(new_n1005), .A3(new_n986), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n981), .B(KEYINPUT114), .C1(new_n977), .C2(new_n1005), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1062), .A2(new_n1032), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n1031), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT115), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(new_n1068), .A3(new_n1031), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(G8), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1029), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1012), .A2(new_n1059), .A3(new_n1072), .A4(G171), .ZN(new_n1073));
  NAND2_X1  g648(.A1(G286), .A2(G8), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n992), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n981), .B1(new_n977), .B2(KEYINPUT45), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n835), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1004), .A2(new_n764), .A3(new_n1006), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1076), .B1(new_n1081), .B2(G8), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1014), .A2(new_n1015), .A3(G2084), .ZN(new_n1083));
  AOI21_X1  g658(.A(G1966), .B1(new_n1000), .B2(new_n992), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT118), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1079), .A2(new_n1080), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(G168), .A3(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1075), .A2(new_n1040), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1082), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1074), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1090), .A2(KEYINPUT62), .A3(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n976), .B1(new_n1073), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1091), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1094), .B(new_n1095), .C1(new_n1096), .C2(new_n1082), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1002), .A2(new_n1009), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT120), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1002), .A2(new_n1003), .A3(new_n1009), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(G301), .B1(new_n1101), .B2(new_n991), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1035), .A2(new_n1058), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1103), .B1(new_n1071), .B2(new_n1070), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1097), .A2(new_n1102), .A3(new_n1104), .A4(KEYINPUT124), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT62), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1093), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1093), .A2(new_n1105), .A3(KEYINPUT125), .A4(new_n1106), .ZN(new_n1110));
  XOR2_X1   g685(.A(G299), .B(KEYINPUT57), .Z(new_n1111));
  NAND3_X1  g686(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1112));
  INV_X1    g687(.A(G1956), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT56), .B(G2072), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n988), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1111), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1007), .A2(new_n808), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n999), .A2(new_n998), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n823), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1122), .A2(new_n612), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1111), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1117), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT60), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1121), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n613), .B1(new_n1127), .B2(KEYINPUT117), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1129), .B(new_n612), .C1(new_n1121), .C2(new_n1126), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1127), .A2(KEYINPUT117), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1131), .A2(new_n1132), .B1(new_n1126), .B2(new_n1121), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n1117), .A2(KEYINPUT61), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1117), .A2(KEYINPUT61), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT58), .B(G1341), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1119), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(G1996), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1137), .B1(new_n988), .B2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1139), .A2(new_n566), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1140), .A2(KEYINPUT59), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(KEYINPUT59), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1134), .A2(new_n1135), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1125), .B1(new_n1133), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT54), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n463), .B1(new_n476), .B2(KEYINPUT122), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(KEYINPUT122), .B2(new_n476), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n799), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n468), .A2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1147), .A2(new_n994), .A3(new_n978), .A4(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n991), .A2(new_n1009), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1151), .A2(G171), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1145), .B1(new_n1102), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT123), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(G171), .ZN(new_n1157));
  OAI221_X1 g732(.A(KEYINPUT54), .B1(new_n1012), .B2(G171), .C1(new_n1155), .C2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1059), .A2(new_n1072), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1144), .A2(new_n1153), .A3(new_n1158), .A4(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1050), .ZN(new_n1163));
  NOR2_X1   g738(.A1(G288), .A2(G1976), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT113), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1044), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1058), .ZN(new_n1167));
  OAI22_X1  g742(.A1(new_n1166), .A2(new_n1051), .B1(new_n1167), .B2(new_n1035), .ZN(new_n1168));
  AOI211_X1 g743(.A(new_n1040), .B(G286), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT63), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1020), .A2(G8), .A3(new_n1034), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n1071), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT116), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n1174), .A2(new_n1175), .A3(new_n1058), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1175), .B1(new_n1174), .B2(new_n1058), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1035), .B(new_n1172), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1171), .B1(new_n1159), .B2(new_n1170), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1168), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1109), .A2(new_n1110), .A3(new_n1162), .A4(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n994), .A2(new_n998), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n789), .B(G1996), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n818), .B(new_n823), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n740), .A2(new_n742), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n740), .A2(new_n742), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(G290), .B(G1986), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1182), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1181), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1182), .ZN(new_n1191));
  NOR3_X1   g766(.A1(new_n1191), .A2(G1986), .A3(G290), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1192), .B(KEYINPUT48), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1193), .B1(new_n1187), .B2(new_n1182), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1138), .A2(KEYINPUT46), .ZN(new_n1195));
  AND3_X1   g770(.A1(new_n1184), .A2(new_n789), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(KEYINPUT46), .B1(new_n1182), .B2(new_n1138), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1197), .A2(KEYINPUT126), .ZN(new_n1198));
  AND2_X1   g773(.A1(new_n1197), .A2(KEYINPUT126), .ZN(new_n1199));
  OAI22_X1  g774(.A1(new_n1196), .A2(new_n1191), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  XOR2_X1   g775(.A(new_n1200), .B(KEYINPUT47), .Z(new_n1201));
  NAND2_X1  g776(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1202));
  OAI22_X1  g777(.A1(new_n1202), .A2(new_n1185), .B1(G2067), .B2(new_n818), .ZN(new_n1203));
  AOI211_X1 g778(.A(new_n1194), .B(new_n1201), .C1(new_n1182), .C2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1190), .A2(new_n1204), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g780(.A1(new_n682), .A2(new_n685), .A3(G319), .ZN(new_n1207));
  OAI211_X1 g781(.A(new_n661), .B(new_n1207), .C1(new_n710), .C2(new_n711), .ZN(new_n1208));
  AOI21_X1  g782(.A(new_n1208), .B1(new_n914), .B2(new_n918), .ZN(new_n1209));
  INV_X1    g783(.A(KEYINPUT127), .ZN(new_n1210));
  AND3_X1   g784(.A1(new_n1209), .A2(new_n971), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g785(.A(new_n1210), .B1(new_n1209), .B2(new_n971), .ZN(new_n1212));
  NOR2_X1   g786(.A1(new_n1211), .A2(new_n1212), .ZN(G308));
  NAND2_X1  g787(.A1(new_n1209), .A2(new_n971), .ZN(new_n1214));
  NAND2_X1  g788(.A1(new_n1214), .A2(KEYINPUT127), .ZN(new_n1215));
  NAND3_X1  g789(.A1(new_n1209), .A2(new_n971), .A3(new_n1210), .ZN(new_n1216));
  NAND2_X1  g790(.A1(new_n1215), .A2(new_n1216), .ZN(G225));
endmodule


