

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581;

  XNOR2_X1 U323 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U324 ( .A(n412), .B(n411), .ZN(n413) );
  NOR2_X1 U325 ( .A1(n458), .A2(n543), .ZN(n429) );
  XOR2_X1 U326 ( .A(n418), .B(n417), .Z(n528) );
  INV_X1 U327 ( .A(G190GAT), .ZN(n453) );
  XNOR2_X1 U328 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U329 ( .A(n456), .B(n455), .ZN(G1351GAT) );
  XOR2_X1 U330 ( .A(G29GAT), .B(G43GAT), .Z(n292) );
  XNOR2_X1 U331 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n291) );
  XNOR2_X1 U332 ( .A(n292), .B(n291), .ZN(n414) );
  XNOR2_X1 U333 ( .A(G50GAT), .B(KEYINPUT76), .ZN(n293) );
  XNOR2_X1 U334 ( .A(n293), .B(G162GAT), .ZN(n317) );
  XOR2_X1 U335 ( .A(n414), .B(n317), .Z(n306) );
  XOR2_X1 U336 ( .A(G99GAT), .B(G85GAT), .Z(n385) );
  XOR2_X1 U337 ( .A(G36GAT), .B(G190GAT), .Z(n356) );
  XOR2_X1 U338 ( .A(n385), .B(n356), .Z(n295) );
  NAND2_X1 U339 ( .A1(G232GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U341 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n297) );
  XNOR2_X1 U342 ( .A(G106GAT), .B(G92GAT), .ZN(n296) );
  XNOR2_X1 U343 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U344 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U345 ( .A(G134GAT), .B(KEYINPUT77), .Z(n340) );
  XOR2_X1 U346 ( .A(KEYINPUT78), .B(KEYINPUT9), .Z(n301) );
  XNOR2_X1 U347 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n340), .B(n302), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n306), .B(n305), .ZN(n553) );
  XOR2_X1 U352 ( .A(G211GAT), .B(G218GAT), .Z(n308) );
  XNOR2_X1 U353 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U355 ( .A(G197GAT), .B(n309), .Z(n357) );
  XOR2_X1 U356 ( .A(KEYINPUT91), .B(KEYINPUT22), .Z(n311) );
  XNOR2_X1 U357 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U359 ( .A(KEYINPUT88), .B(n312), .Z(n314) );
  NAND2_X1 U360 ( .A1(G228GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U362 ( .A(G22GAT), .B(G155GAT), .Z(n367) );
  XOR2_X1 U363 ( .A(n315), .B(n367), .Z(n319) );
  XNOR2_X1 U364 ( .A(G106GAT), .B(G78GAT), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n316), .B(G148GAT), .ZN(n380) );
  XNOR2_X1 U366 ( .A(n317), .B(n380), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U368 ( .A(n357), .B(n320), .ZN(n324) );
  XOR2_X1 U369 ( .A(KEYINPUT90), .B(KEYINPUT2), .Z(n322) );
  XNOR2_X1 U370 ( .A(KEYINPUT3), .B(KEYINPUT89), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U372 ( .A(G141GAT), .B(n323), .ZN(n337) );
  XNOR2_X1 U373 ( .A(n324), .B(n337), .ZN(n463) );
  XOR2_X1 U374 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n326) );
  XNOR2_X1 U375 ( .A(G148GAT), .B(G155GAT), .ZN(n325) );
  XNOR2_X1 U376 ( .A(n326), .B(n325), .ZN(n330) );
  XOR2_X1 U377 ( .A(G85GAT), .B(G162GAT), .Z(n328) );
  XNOR2_X1 U378 ( .A(G29GAT), .B(G127GAT), .ZN(n327) );
  XNOR2_X1 U379 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U380 ( .A(n330), .B(n329), .ZN(n347) );
  XOR2_X1 U381 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n332) );
  XNOR2_X1 U382 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n331) );
  XNOR2_X1 U383 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U384 ( .A(G57GAT), .B(n333), .Z(n335) );
  NAND2_X1 U385 ( .A1(G225GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U386 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U387 ( .A(n336), .B(KEYINPUT92), .Z(n339) );
  XOR2_X1 U388 ( .A(n337), .B(KEYINPUT93), .Z(n338) );
  XNOR2_X1 U389 ( .A(n339), .B(n338), .ZN(n341) );
  XOR2_X1 U390 ( .A(n341), .B(n340), .Z(n345) );
  XOR2_X1 U391 ( .A(G113GAT), .B(G1GAT), .Z(n404) );
  XOR2_X1 U392 ( .A(G120GAT), .B(KEYINPUT82), .Z(n343) );
  XNOR2_X1 U393 ( .A(KEYINPUT0), .B(KEYINPUT81), .ZN(n342) );
  XNOR2_X1 U394 ( .A(n343), .B(n342), .ZN(n433) );
  XNOR2_X1 U395 ( .A(n404), .B(n433), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U397 ( .A(n347), .B(n346), .Z(n469) );
  XNOR2_X1 U398 ( .A(KEYINPUT84), .B(KEYINPUT85), .ZN(n348) );
  XNOR2_X1 U399 ( .A(n348), .B(G183GAT), .ZN(n349) );
  XOR2_X1 U400 ( .A(n349), .B(KEYINPUT18), .Z(n351) );
  XNOR2_X1 U401 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n350) );
  XOR2_X1 U402 ( .A(n351), .B(n350), .Z(n437) );
  XOR2_X1 U403 ( .A(KEYINPUT98), .B(KEYINPUT96), .Z(n353) );
  NAND2_X1 U404 ( .A1(G226GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U406 ( .A(KEYINPUT97), .B(n354), .ZN(n361) );
  XNOR2_X1 U407 ( .A(G176GAT), .B(G92GAT), .ZN(n355) );
  XNOR2_X1 U408 ( .A(n355), .B(G64GAT), .ZN(n394) );
  XOR2_X1 U409 ( .A(n394), .B(n356), .Z(n359) );
  XOR2_X1 U410 ( .A(G169GAT), .B(G8GAT), .Z(n403) );
  XNOR2_X1 U411 ( .A(n403), .B(n357), .ZN(n358) );
  XNOR2_X1 U412 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U413 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U414 ( .A(n437), .B(n362), .Z(n458) );
  INV_X1 U415 ( .A(n553), .ZN(n539) );
  XOR2_X1 U416 ( .A(KEYINPUT36), .B(n539), .Z(n579) );
  XOR2_X1 U417 ( .A(KEYINPUT79), .B(KEYINPUT15), .Z(n364) );
  XNOR2_X1 U418 ( .A(G8GAT), .B(G64GAT), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n366) );
  XNOR2_X1 U420 ( .A(G71GAT), .B(G57GAT), .ZN(n365) );
  XNOR2_X1 U421 ( .A(n365), .B(KEYINPUT13), .ZN(n393) );
  XOR2_X1 U422 ( .A(n366), .B(n393), .Z(n369) );
  XOR2_X1 U423 ( .A(G15GAT), .B(G127GAT), .Z(n434) );
  XNOR2_X1 U424 ( .A(n434), .B(n367), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U426 ( .A(KEYINPUT80), .B(KEYINPUT12), .Z(n371) );
  NAND2_X1 U427 ( .A1(G231GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U429 ( .A(n373), .B(n372), .Z(n378) );
  XOR2_X1 U430 ( .A(G78GAT), .B(G211GAT), .Z(n375) );
  XNOR2_X1 U431 ( .A(G1GAT), .B(G183GAT), .ZN(n374) );
  XNOR2_X1 U432 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n376), .B(KEYINPUT14), .ZN(n377) );
  XOR2_X1 U434 ( .A(n378), .B(n377), .Z(n535) );
  INV_X1 U435 ( .A(n535), .ZN(n576) );
  NOR2_X1 U436 ( .A1(n579), .A2(n576), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n379), .B(KEYINPUT45), .ZN(n399) );
  XOR2_X1 U438 ( .A(n380), .B(KEYINPUT72), .Z(n382) );
  NAND2_X1 U439 ( .A1(G230GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U440 ( .A(n382), .B(n381), .ZN(n398) );
  XOR2_X1 U441 ( .A(KEYINPUT75), .B(KEYINPUT70), .Z(n384) );
  XNOR2_X1 U442 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n383) );
  XOR2_X1 U443 ( .A(n384), .B(n383), .Z(n386) );
  XNOR2_X1 U444 ( .A(n386), .B(n385), .ZN(n388) );
  XNOR2_X1 U445 ( .A(G120GAT), .B(G204GAT), .ZN(n387) );
  XNOR2_X1 U446 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U447 ( .A(KEYINPUT71), .B(KEYINPUT33), .Z(n390) );
  XNOR2_X1 U448 ( .A(KEYINPUT74), .B(KEYINPUT73), .ZN(n389) );
  XOR2_X1 U449 ( .A(n390), .B(n389), .Z(n391) );
  XNOR2_X1 U450 ( .A(n392), .B(n391), .ZN(n396) );
  XNOR2_X1 U451 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U453 ( .A(n398), .B(n397), .ZN(n572) );
  NAND2_X1 U454 ( .A1(n399), .A2(n572), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n400), .B(KEYINPUT115), .ZN(n419) );
  XOR2_X1 U456 ( .A(G141GAT), .B(G197GAT), .Z(n402) );
  XNOR2_X1 U457 ( .A(G15GAT), .B(G22GAT), .ZN(n401) );
  XNOR2_X1 U458 ( .A(n402), .B(n401), .ZN(n418) );
  XOR2_X1 U459 ( .A(G50GAT), .B(G36GAT), .Z(n406) );
  XNOR2_X1 U460 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n412) );
  XOR2_X1 U462 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n408) );
  XNOR2_X1 U463 ( .A(KEYINPUT30), .B(KEYINPUT66), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n410) );
  AND2_X1 U465 ( .A1(G229GAT), .A2(G233GAT), .ZN(n409) );
  XOR2_X1 U466 ( .A(KEYINPUT67), .B(n413), .Z(n416) );
  XNOR2_X1 U467 ( .A(n414), .B(KEYINPUT29), .ZN(n415) );
  XNOR2_X1 U468 ( .A(n416), .B(n415), .ZN(n417) );
  INV_X1 U469 ( .A(n528), .ZN(n568) );
  NAND2_X1 U470 ( .A1(n419), .A2(n568), .ZN(n427) );
  XOR2_X1 U471 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n421) );
  XNOR2_X1 U472 ( .A(KEYINPUT41), .B(n572), .ZN(n548) );
  NAND2_X1 U473 ( .A1(n548), .A2(n528), .ZN(n420) );
  XNOR2_X1 U474 ( .A(n421), .B(n420), .ZN(n422) );
  NAND2_X1 U475 ( .A1(n576), .A2(n422), .ZN(n423) );
  NOR2_X1 U476 ( .A1(n539), .A2(n423), .ZN(n425) );
  XNOR2_X1 U477 ( .A(KEYINPUT47), .B(KEYINPUT114), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n425), .B(n424), .ZN(n426) );
  NAND2_X1 U479 ( .A1(n427), .A2(n426), .ZN(n428) );
  XOR2_X1 U480 ( .A(KEYINPUT48), .B(n428), .Z(n543) );
  XNOR2_X1 U481 ( .A(n429), .B(KEYINPUT54), .ZN(n430) );
  AND2_X1 U482 ( .A1(n469), .A2(n430), .ZN(n567) );
  NAND2_X1 U483 ( .A1(n463), .A2(n567), .ZN(n431) );
  XNOR2_X1 U484 ( .A(n431), .B(KEYINPUT122), .ZN(n432) );
  XNOR2_X1 U485 ( .A(n432), .B(KEYINPUT55), .ZN(n452) );
  XOR2_X1 U486 ( .A(n434), .B(n433), .Z(n436) );
  XNOR2_X1 U487 ( .A(G43GAT), .B(G99GAT), .ZN(n435) );
  XNOR2_X1 U488 ( .A(n436), .B(n435), .ZN(n438) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n451) );
  XOR2_X1 U490 ( .A(KEYINPUT83), .B(KEYINPUT86), .Z(n440) );
  XNOR2_X1 U491 ( .A(G190GAT), .B(G134GAT), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U493 ( .A(G71GAT), .B(G176GAT), .Z(n442) );
  XNOR2_X1 U494 ( .A(G169GAT), .B(KEYINPUT20), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U496 ( .A(n444), .B(n443), .Z(n449) );
  XOR2_X1 U497 ( .A(KEYINPUT64), .B(KEYINPUT87), .Z(n446) );
  NAND2_X1 U498 ( .A1(G227GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U500 ( .A(G113GAT), .B(n447), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U502 ( .A(n451), .B(n450), .Z(n459) );
  INV_X1 U503 ( .A(n459), .ZN(n524) );
  NAND2_X1 U504 ( .A1(n452), .A2(n524), .ZN(n563) );
  NOR2_X1 U505 ( .A1(n553), .A2(n563), .ZN(n456) );
  XNOR2_X1 U506 ( .A(KEYINPUT126), .B(KEYINPUT58), .ZN(n454) );
  XNOR2_X1 U507 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n476) );
  INV_X1 U508 ( .A(n469), .ZN(n513) );
  NAND2_X1 U509 ( .A1(n528), .A2(n572), .ZN(n485) );
  NOR2_X1 U510 ( .A1(n539), .A2(n576), .ZN(n457) );
  XNOR2_X1 U511 ( .A(n457), .B(KEYINPUT16), .ZN(n473) );
  INV_X1 U512 ( .A(n458), .ZN(n517) );
  XNOR2_X1 U513 ( .A(KEYINPUT27), .B(n517), .ZN(n462) );
  NAND2_X1 U514 ( .A1(n513), .A2(n462), .ZN(n542) );
  XOR2_X1 U515 ( .A(KEYINPUT28), .B(n463), .Z(n521) );
  NOR2_X1 U516 ( .A1(n542), .A2(n521), .ZN(n525) );
  NAND2_X1 U517 ( .A1(n459), .A2(n525), .ZN(n460) );
  XOR2_X1 U518 ( .A(KEYINPUT99), .B(n460), .Z(n472) );
  NOR2_X1 U519 ( .A1(n463), .A2(n524), .ZN(n461) );
  XNOR2_X1 U520 ( .A(n461), .B(KEYINPUT26), .ZN(n566) );
  NAND2_X1 U521 ( .A1(n462), .A2(n566), .ZN(n468) );
  NAND2_X1 U522 ( .A1(n524), .A2(n517), .ZN(n464) );
  NAND2_X1 U523 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n465), .B(KEYINPUT25), .ZN(n466) );
  XOR2_X1 U525 ( .A(KEYINPUT100), .B(n466), .Z(n467) );
  NAND2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n470) );
  NAND2_X1 U527 ( .A1(n470), .A2(n469), .ZN(n471) );
  NAND2_X1 U528 ( .A1(n472), .A2(n471), .ZN(n482) );
  NAND2_X1 U529 ( .A1(n473), .A2(n482), .ZN(n474) );
  XOR2_X1 U530 ( .A(KEYINPUT101), .B(n474), .Z(n503) );
  NOR2_X1 U531 ( .A1(n485), .A2(n503), .ZN(n480) );
  NAND2_X1 U532 ( .A1(n513), .A2(n480), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n476), .B(n475), .ZN(G1324GAT) );
  NAND2_X1 U534 ( .A1(n480), .A2(n517), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n477), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(G15GAT), .B(KEYINPUT35), .Z(n479) );
  NAND2_X1 U537 ( .A1(n480), .A2(n524), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(G1326GAT) );
  NAND2_X1 U539 ( .A1(n521), .A2(n480), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n481), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U541 ( .A1(n576), .A2(n482), .ZN(n483) );
  NOR2_X1 U542 ( .A1(n483), .A2(n579), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n484), .B(KEYINPUT37), .ZN(n511) );
  NOR2_X1 U544 ( .A1(n511), .A2(n485), .ZN(n487) );
  XNOR2_X1 U545 ( .A(KEYINPUT104), .B(KEYINPUT38), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U547 ( .A(KEYINPUT103), .B(n488), .Z(n499) );
  NAND2_X1 U548 ( .A1(n513), .A2(n499), .ZN(n490) );
  XOR2_X1 U549 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U551 ( .A(G29GAT), .B(n491), .ZN(G1328GAT) );
  XOR2_X1 U552 ( .A(G36GAT), .B(KEYINPUT105), .Z(n493) );
  NAND2_X1 U553 ( .A1(n499), .A2(n517), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(G1329GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT40), .B(KEYINPUT108), .Z(n495) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(KEYINPUT107), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(n498) );
  NAND2_X1 U558 ( .A1(n524), .A2(n499), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n496), .B(KEYINPUT106), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(G1330GAT) );
  XOR2_X1 U561 ( .A(G50GAT), .B(KEYINPUT109), .Z(n501) );
  NAND2_X1 U562 ( .A1(n499), .A2(n521), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(G1331GAT) );
  NAND2_X1 U564 ( .A1(n568), .A2(n548), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n502), .B(KEYINPUT110), .ZN(n512) );
  NOR2_X1 U566 ( .A1(n512), .A2(n503), .ZN(n508) );
  NAND2_X1 U567 ( .A1(n513), .A2(n508), .ZN(n504) );
  XNOR2_X1 U568 ( .A(KEYINPUT42), .B(n504), .ZN(n505) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(n505), .ZN(G1332GAT) );
  NAND2_X1 U570 ( .A1(n508), .A2(n517), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n506), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U572 ( .A1(n524), .A2(n508), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n507), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U575 ( .A1(n508), .A2(n521), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n515) );
  NOR2_X1 U578 ( .A1(n512), .A2(n511), .ZN(n520) );
  NAND2_X1 U579 ( .A1(n520), .A2(n513), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  NAND2_X1 U582 ( .A1(n520), .A2(n517), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n518), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U584 ( .A1(n524), .A2(n520), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(KEYINPUT44), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n530) );
  NAND2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U591 ( .A1(n526), .A2(n543), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n527), .B(KEYINPUT116), .ZN(n538) );
  NAND2_X1 U593 ( .A1(n528), .A2(n538), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G113GAT), .B(n531), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U597 ( .A1(n548), .A2(n538), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U599 ( .A(G120GAT), .B(n534), .Z(G1341GAT) );
  NAND2_X1 U600 ( .A1(n538), .A2(n535), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n536), .B(KEYINPUT50), .ZN(n537) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U604 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  NOR2_X1 U606 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U607 ( .A1(n544), .A2(n566), .ZN(n552) );
  NOR2_X1 U608 ( .A1(n568), .A2(n552), .ZN(n545) );
  XOR2_X1 U609 ( .A(G141GAT), .B(n545), .Z(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n547) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(n550) );
  INV_X1 U613 ( .A(n548), .ZN(n559) );
  NOR2_X1 U614 ( .A1(n559), .A2(n552), .ZN(n549) );
  XOR2_X1 U615 ( .A(n550), .B(n549), .Z(G1345GAT) );
  NOR2_X1 U616 ( .A1(n576), .A2(n552), .ZN(n551) );
  XOR2_X1 U617 ( .A(G155GAT), .B(n551), .Z(G1346GAT) );
  NOR2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n555) );
  XNOR2_X1 U619 ( .A(G162GAT), .B(KEYINPUT121), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(G1347GAT) );
  XNOR2_X1 U621 ( .A(G169GAT), .B(KEYINPUT123), .ZN(n558) );
  NOR2_X1 U622 ( .A1(n563), .A2(n568), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(KEYINPUT124), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1348GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n563), .ZN(n561) );
  XNOR2_X1 U626 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(n562), .ZN(G1349GAT) );
  NOR2_X1 U629 ( .A1(n576), .A2(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(G183GAT), .B(KEYINPUT125), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1350GAT) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n578) );
  NOR2_X1 U633 ( .A1(n568), .A2(n578), .ZN(n570) );
  XNOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(n571), .ZN(G1352GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n578), .ZN(n574) );
  XNOR2_X1 U638 ( .A(KEYINPUT61), .B(KEYINPUT127), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U640 ( .A(G204GAT), .B(n575), .Z(G1353GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n578), .ZN(n577) );
  XOR2_X1 U642 ( .A(G211GAT), .B(n577), .Z(G1354GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT62), .B(n580), .Z(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

