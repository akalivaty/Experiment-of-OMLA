

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n718, n719, n720, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751;

  XNOR2_X1 U372 ( .A(n715), .B(n716), .ZN(n352) );
  XNOR2_X1 U373 ( .A(n720), .B(n718), .ZN(n350) );
  NOR2_X1 U374 ( .A1(n641), .A2(n657), .ZN(n563) );
  NOR2_X1 U375 ( .A1(n550), .A2(n617), .ZN(n570) );
  XNOR2_X1 U376 ( .A(n543), .B(KEYINPUT22), .ZN(n550) );
  XNOR2_X1 U377 ( .A(n535), .B(KEYINPUT33), .ZN(n696) );
  INV_X1 U378 ( .A(n559), .ZN(n354) );
  NAND2_X1 U379 ( .A1(n558), .A2(n608), .ZN(n535) );
  XNOR2_X1 U380 ( .A(n390), .B(n587), .ZN(n664) );
  NOR2_X1 U381 ( .A1(n565), .A2(n566), .ZN(n654) );
  XNOR2_X1 U382 ( .A(n541), .B(n351), .ZN(n608) );
  INV_X1 U383 ( .A(KEYINPUT6), .ZN(n351) );
  XNOR2_X1 U384 ( .A(n732), .B(n389), .ZN(n513) );
  XNOR2_X1 U385 ( .A(n485), .B(n484), .ZN(n732) );
  XNOR2_X1 U386 ( .A(n489), .B(G134), .ZN(n507) );
  XNOR2_X1 U387 ( .A(G113), .B(G143), .ZN(n466) );
  XNOR2_X1 U388 ( .A(n373), .B(G128), .ZN(n489) );
  INV_X2 U389 ( .A(G953), .ZN(n487) );
  NOR2_X1 U390 ( .A1(G953), .A2(G237), .ZN(n525) );
  INV_X1 U391 ( .A(G143), .ZN(n373) );
  XNOR2_X1 U392 ( .A(n481), .B(KEYINPUT3), .ZN(n482) );
  XNOR2_X1 U393 ( .A(n480), .B(n479), .ZN(n483) );
  NOR2_X1 U394 ( .A1(n350), .A2(n722), .ZN(G66) );
  XNOR2_X2 U395 ( .A(n385), .B(n534), .ZN(n541) );
  NOR2_X1 U396 ( .A1(n352), .A2(n722), .ZN(G63) );
  NAND2_X2 U397 ( .A1(n391), .A2(n422), .ZN(n731) );
  XNOR2_X2 U398 ( .A(n353), .B(n538), .ZN(n748) );
  NOR2_X2 U399 ( .A1(n537), .A2(n599), .ZN(n353) );
  AND2_X2 U400 ( .A1(n432), .A2(n573), .ZN(n360) );
  XNOR2_X2 U401 ( .A(n505), .B(n504), .ZN(n559) );
  NOR2_X2 U402 ( .A1(n405), .A2(n404), .ZN(n615) );
  NOR2_X2 U403 ( .A1(n597), .A2(n586), .ZN(n585) );
  XNOR2_X2 U404 ( .A(n557), .B(KEYINPUT99), .ZN(n641) );
  OR2_X2 U405 ( .A1(n748), .A2(KEYINPUT44), .ZN(n540) );
  AND2_X2 U406 ( .A1(n393), .A2(n360), .ZN(n431) );
  XNOR2_X2 U407 ( .A(KEYINPUT32), .B(n551), .ZN(n751) );
  NOR2_X2 U408 ( .A1(n646), .A2(n751), .ZN(n553) );
  BUF_X1 U409 ( .A(n541), .Z(n679) );
  INV_X1 U410 ( .A(KEYINPUT4), .ZN(n371) );
  INV_X1 U411 ( .A(G125), .ZN(n384) );
  NOR2_X1 U412 ( .A1(n654), .A2(n658), .ZN(n691) );
  XNOR2_X1 U413 ( .A(n419), .B(KEYINPUT106), .ZN(n689) );
  XNOR2_X1 U414 ( .A(n591), .B(KEYINPUT1), .ZN(n674) );
  XNOR2_X1 U415 ( .A(n518), .B(n517), .ZN(n676) );
  XNOR2_X1 U416 ( .A(n371), .B(KEYINPUT68), .ZN(n506) );
  XNOR2_X1 U417 ( .A(n384), .B(G146), .ZN(n486) );
  XOR2_X1 U418 ( .A(G131), .B(G140), .Z(n509) );
  BUF_X1 U419 ( .A(n611), .Z(n355) );
  OR2_X1 U420 ( .A1(n628), .A2(n624), .ZN(n356) );
  NAND2_X1 U421 ( .A1(n664), .A2(n593), .ZN(n421) );
  OR2_X2 U422 ( .A1(n628), .A2(n624), .ZN(n742) );
  AND2_X1 U423 ( .A1(n750), .A2(KEYINPUT46), .ZN(n404) );
  AND2_X1 U424 ( .A1(n411), .A2(n407), .ZN(n406) );
  XNOR2_X1 U425 ( .A(n412), .B(n516), .ZN(n523) );
  XNOR2_X1 U426 ( .A(n742), .B(n450), .ZN(n449) );
  INV_X1 U427 ( .A(KEYINPUT76), .ZN(n450) );
  OR2_X1 U428 ( .A1(n566), .A2(n564), .ZN(n419) );
  XNOR2_X1 U429 ( .A(n398), .B(n366), .ZN(n628) );
  XNOR2_X1 U430 ( .A(KEYINPUT90), .B(n662), .ZN(n614) );
  INV_X1 U431 ( .A(n676), .ZN(n379) );
  NOR2_X1 U432 ( .A1(n633), .A2(G902), .ZN(n385) );
  XNOR2_X1 U433 ( .A(n524), .B(n453), .ZN(n452) );
  OR2_X1 U434 ( .A1(n718), .A2(G902), .ZN(n454) );
  INV_X1 U435 ( .A(KEYINPUT25), .ZN(n453) );
  XOR2_X1 U436 ( .A(G110), .B(G107), .Z(n485) );
  XNOR2_X1 U437 ( .A(n447), .B(n446), .ZN(n445) );
  XNOR2_X1 U438 ( .A(G119), .B(G128), .ZN(n446) );
  XNOR2_X1 U439 ( .A(n448), .B(G140), .ZN(n447) );
  INV_X1 U440 ( .A(G110), .ZN(n448) );
  XNOR2_X1 U441 ( .A(n444), .B(n443), .ZN(n442) );
  XNOR2_X1 U442 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n444) );
  XNOR2_X1 U443 ( .A(G137), .B(KEYINPUT80), .ZN(n443) );
  XNOR2_X1 U444 ( .A(n458), .B(n457), .ZN(n519) );
  XNOR2_X1 U445 ( .A(n456), .B(KEYINPUT69), .ZN(n458) );
  NAND2_X1 U446 ( .A1(n487), .A2(G234), .ZN(n456) );
  XOR2_X1 U447 ( .A(KEYINPUT104), .B(KEYINPUT9), .Z(n461) );
  NAND2_X1 U448 ( .A1(n402), .A2(n670), .ZN(n401) );
  XNOR2_X1 U449 ( .A(n493), .B(KEYINPUT83), .ZN(n494) );
  INV_X1 U450 ( .A(KEYINPUT39), .ZN(n584) );
  NAND2_X1 U451 ( .A1(n417), .A2(n415), .ZN(n616) );
  NOR2_X1 U452 ( .A1(n610), .A2(n416), .ZN(n415) );
  XNOR2_X1 U453 ( .A(n609), .B(KEYINPUT109), .ZN(n417) );
  INV_X1 U454 ( .A(n686), .ZN(n416) );
  BUF_X1 U455 ( .A(n591), .Z(n394) );
  XNOR2_X1 U456 ( .A(n400), .B(n375), .ZN(n566) );
  XNOR2_X1 U457 ( .A(n399), .B(n420), .ZN(n375) );
  INV_X1 U458 ( .A(G478), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n669), .B(n388), .ZN(n387) );
  INV_X1 U460 ( .A(KEYINPUT86), .ZN(n388) );
  AND2_X1 U461 ( .A1(n606), .A2(n605), .ZN(n411) );
  INV_X1 U462 ( .A(KEYINPUT72), .ZN(n479) );
  XNOR2_X1 U463 ( .A(G101), .B(G131), .ZN(n529) );
  INV_X1 U464 ( .A(KEYINPUT5), .ZN(n528) );
  XOR2_X1 U465 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n527) );
  XNOR2_X1 U466 ( .A(KEYINPUT16), .B(G122), .ZN(n423) );
  XOR2_X1 U467 ( .A(G104), .B(G122), .Z(n467) );
  XNOR2_X1 U468 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n468) );
  XOR2_X1 U469 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n469) );
  XNOR2_X1 U470 ( .A(n433), .B(n488), .ZN(n491) );
  XNOR2_X1 U471 ( .A(n486), .B(n434), .ZN(n433) );
  XNOR2_X1 U472 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n434) );
  OR2_X1 U473 ( .A1(G237), .A2(G902), .ZN(n492) );
  INV_X1 U474 ( .A(KEYINPUT93), .ZN(n413) );
  XNOR2_X1 U475 ( .A(KEYINPUT15), .B(G902), .ZN(n414) );
  NAND2_X1 U476 ( .A1(n687), .A2(n686), .ZN(n690) );
  INV_X1 U477 ( .A(KEYINPUT105), .ZN(n420) );
  NAND2_X1 U478 ( .A1(n431), .A2(n429), .ZN(n575) );
  INV_X1 U479 ( .A(KEYINPUT73), .ZN(n389) );
  NAND2_X1 U480 ( .A1(n354), .A2(n378), .ZN(n543) );
  NOR2_X1 U481 ( .A1(n689), .A2(n379), .ZN(n378) );
  INV_X1 U482 ( .A(KEYINPUT77), .ZN(n582) );
  XNOR2_X1 U483 ( .A(n520), .B(n522), .ZN(n370) );
  XNOR2_X1 U484 ( .A(n445), .B(n442), .ZN(n520) );
  XNOR2_X1 U485 ( .A(n374), .B(n464), .ZN(n716) );
  XNOR2_X1 U486 ( .A(n463), .B(n465), .ZN(n374) );
  INV_X1 U487 ( .A(KEYINPUT40), .ZN(n395) );
  NOR2_X1 U488 ( .A1(n616), .A2(n355), .ZN(n612) );
  XNOR2_X1 U489 ( .A(n562), .B(n561), .ZN(n657) );
  XNOR2_X1 U490 ( .A(n560), .B(KEYINPUT100), .ZN(n561) );
  INV_X1 U491 ( .A(n602), .ZN(n650) );
  NOR2_X1 U492 ( .A1(n559), .A2(n394), .ZN(n555) );
  NAND2_X1 U493 ( .A1(n381), .A2(n426), .ZN(n372) );
  XNOR2_X1 U494 ( .A(n637), .B(n636), .ZN(n381) );
  INV_X1 U495 ( .A(KEYINPUT60), .ZN(n376) );
  NAND2_X1 U496 ( .A1(n383), .A2(n426), .ZN(n377) );
  XNOR2_X1 U497 ( .A(n714), .B(n365), .ZN(n383) );
  XNOR2_X1 U498 ( .A(n710), .B(n709), .ZN(n711) );
  INV_X1 U499 ( .A(KEYINPUT56), .ZN(n424) );
  NAND2_X1 U500 ( .A1(n427), .A2(n426), .ZN(n425) );
  XNOR2_X1 U501 ( .A(n428), .B(n364), .ZN(n427) );
  NOR2_X1 U502 ( .A1(n704), .A2(G953), .ZN(n386) );
  XNOR2_X1 U503 ( .A(KEYINPUT113), .B(KEYINPUT42), .ZN(n357) );
  XOR2_X1 U504 ( .A(n491), .B(n490), .Z(n358) );
  XOR2_X1 U505 ( .A(n532), .B(n533), .Z(n359) );
  AND2_X1 U506 ( .A1(n672), .A2(n671), .ZN(n361) );
  XOR2_X1 U507 ( .A(G122), .B(KEYINPUT16), .Z(n362) );
  XNOR2_X1 U508 ( .A(KEYINPUT74), .B(KEYINPUT34), .ZN(n363) );
  XOR2_X1 U509 ( .A(n706), .B(n455), .Z(n364) );
  XNOR2_X1 U510 ( .A(n370), .B(n521), .ZN(n718) );
  XNOR2_X1 U511 ( .A(n712), .B(KEYINPUT59), .ZN(n365) );
  XNOR2_X1 U512 ( .A(n414), .B(n413), .ZN(n625) );
  XNOR2_X1 U513 ( .A(KEYINPUT48), .B(KEYINPUT70), .ZN(n366) );
  NOR2_X1 U514 ( .A1(G952), .A2(n487), .ZN(n722) );
  INV_X1 U515 ( .A(n722), .ZN(n426) );
  NAND2_X1 U516 ( .A1(n367), .A2(n654), .ZN(n396) );
  XNOR2_X1 U517 ( .A(n585), .B(n584), .ZN(n367) );
  NAND2_X1 U518 ( .A1(n367), .A2(n658), .ZN(n663) );
  XNOR2_X1 U519 ( .A(n368), .B(n514), .ZN(n708) );
  XNOR2_X1 U520 ( .A(n368), .B(n359), .ZN(n633) );
  XNOR2_X2 U521 ( .A(n739), .B(G146), .ZN(n368) );
  AND2_X1 U522 ( .A1(n571), .A2(n638), .ZN(n432) );
  XNOR2_X2 U523 ( .A(n369), .B(n358), .ZN(n706) );
  XNOR2_X2 U524 ( .A(n731), .B(n513), .ZN(n369) );
  NOR2_X1 U525 ( .A1(n727), .A2(n625), .ZN(n451) );
  NOR2_X1 U526 ( .A1(n394), .A2(n590), .ZN(n593) );
  NAND2_X1 U527 ( .A1(n625), .A2(G234), .ZN(n412) );
  XNOR2_X1 U528 ( .A(n372), .B(KEYINPUT63), .ZN(G57) );
  NOR2_X2 U529 ( .A1(n690), .A2(n689), .ZN(n390) );
  NAND2_X1 U530 ( .A1(n553), .A2(n554), .ZN(n380) );
  XNOR2_X1 U531 ( .A(n377), .B(n376), .ZN(G60) );
  NAND2_X1 U532 ( .A1(n380), .A2(KEYINPUT44), .ZN(n393) );
  INV_X1 U533 ( .A(n382), .ZN(n408) );
  NOR2_X1 U534 ( .A1(n750), .A2(n409), .ZN(n382) );
  XNOR2_X1 U535 ( .A(n437), .B(n436), .ZN(n435) );
  NAND2_X1 U536 ( .A1(n361), .A2(n386), .ZN(n705) );
  NAND2_X1 U537 ( .A1(n387), .A2(n670), .ZN(n671) );
  XNOR2_X2 U538 ( .A(n507), .B(n508), .ZN(n739) );
  INV_X1 U539 ( .A(n533), .ZN(n392) );
  XNOR2_X2 U540 ( .A(n483), .B(n482), .ZN(n533) );
  NAND2_X1 U541 ( .A1(n392), .A2(n362), .ZN(n391) );
  NOR2_X1 U542 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X2 U543 ( .A(n396), .B(n395), .ZN(n750) );
  XNOR2_X2 U544 ( .A(n397), .B(n496), .ZN(n594) );
  NAND2_X1 U545 ( .A1(n621), .A2(n686), .ZN(n397) );
  NAND2_X1 U546 ( .A1(n706), .A2(n625), .ZN(n418) );
  XNOR2_X1 U547 ( .A(n540), .B(KEYINPUT67), .ZN(n430) );
  NAND2_X1 U548 ( .A1(n615), .A2(n614), .ZN(n398) );
  NOR2_X1 U549 ( .A1(n716), .A2(G902), .ZN(n400) );
  XNOR2_X2 U550 ( .A(n401), .B(KEYINPUT65), .ZN(n713) );
  NAND2_X1 U551 ( .A1(n403), .A2(n627), .ZN(n402) );
  NAND2_X1 U552 ( .A1(n449), .A2(n451), .ZN(n403) );
  NAND2_X1 U553 ( .A1(n408), .A2(n406), .ZN(n405) );
  NAND2_X1 U554 ( .A1(n749), .A2(KEYINPUT46), .ZN(n407) );
  NAND2_X1 U555 ( .A1(n410), .A2(n592), .ZN(n409) );
  INV_X1 U556 ( .A(n749), .ZN(n410) );
  XNOR2_X2 U557 ( .A(n418), .B(n494), .ZN(n621) );
  INV_X1 U558 ( .A(n687), .ZN(n586) );
  XNOR2_X2 U559 ( .A(n611), .B(KEYINPUT38), .ZN(n687) );
  XNOR2_X2 U560 ( .A(n421), .B(n357), .ZN(n749) );
  NAND2_X1 U561 ( .A1(n533), .A2(n423), .ZN(n422) );
  INV_X2 U562 ( .A(n621), .ZN(n611) );
  XNOR2_X2 U563 ( .A(n515), .B(G469), .ZN(n591) );
  XNOR2_X1 U564 ( .A(n425), .B(n424), .ZN(G51) );
  NAND2_X1 U565 ( .A1(n713), .A2(G210), .ZN(n428) );
  NAND2_X1 U566 ( .A1(n430), .A2(n553), .ZN(n429) );
  NAND2_X1 U567 ( .A1(n438), .A2(n435), .ZN(n583) );
  XNOR2_X1 U568 ( .A(n581), .B(KEYINPUT112), .ZN(n436) );
  NAND2_X1 U569 ( .A1(n541), .A2(n686), .ZN(n437) );
  XNOR2_X1 U570 ( .A(n440), .B(n439), .ZN(n438) );
  INV_X1 U571 ( .A(KEYINPUT78), .ZN(n439) );
  NAND2_X1 U572 ( .A1(n441), .A2(n542), .ZN(n440) );
  NOR2_X1 U573 ( .A1(n591), .A2(n588), .ZN(n441) );
  XNOR2_X2 U574 ( .A(n454), .B(n452), .ZN(n542) );
  XNOR2_X2 U575 ( .A(G113), .B(G119), .ZN(n480) );
  XNOR2_X1 U576 ( .A(n583), .B(n582), .ZN(n597) );
  XNOR2_X1 U577 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n455) );
  XNOR2_X1 U578 ( .A(n529), .B(n528), .ZN(n530) );
  INV_X1 U579 ( .A(KEYINPUT46), .ZN(n592) );
  XNOR2_X1 U580 ( .A(n531), .B(n530), .ZN(n532) );
  INV_X1 U581 ( .A(KEYINPUT30), .ZN(n581) );
  INV_X1 U582 ( .A(KEYINPUT79), .ZN(n495) );
  INV_X1 U583 ( .A(n747), .ZN(n623) );
  XNOR2_X1 U584 ( .A(n495), .B(KEYINPUT19), .ZN(n496) );
  NAND2_X1 U585 ( .A1(n623), .A2(n663), .ZN(n624) );
  XNOR2_X1 U586 ( .A(n512), .B(n513), .ZN(n514) );
  XNOR2_X1 U587 ( .A(n708), .B(n707), .ZN(n709) );
  INV_X1 U588 ( .A(KEYINPUT35), .ZN(n538) );
  INV_X1 U589 ( .A(n507), .ZN(n465) );
  XOR2_X1 U590 ( .A(KEYINPUT87), .B(KEYINPUT8), .Z(n457) );
  NAND2_X1 U591 ( .A1(n519), .A2(G217), .ZN(n464) );
  XOR2_X1 U592 ( .A(KEYINPUT7), .B(G107), .Z(n460) );
  XNOR2_X1 U593 ( .A(G116), .B(G122), .ZN(n459) );
  XNOR2_X1 U594 ( .A(n460), .B(n459), .ZN(n462) );
  XNOR2_X1 U595 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U596 ( .A(KEYINPUT13), .B(G475), .ZN(n477) );
  XNOR2_X1 U597 ( .A(n467), .B(n466), .ZN(n471) );
  XNOR2_X1 U598 ( .A(n469), .B(n468), .ZN(n470) );
  XOR2_X1 U599 ( .A(n471), .B(n470), .Z(n473) );
  NAND2_X1 U600 ( .A1(G214), .A2(n525), .ZN(n472) );
  XNOR2_X1 U601 ( .A(n473), .B(n472), .ZN(n475) );
  XNOR2_X1 U602 ( .A(n486), .B(KEYINPUT10), .ZN(n522) );
  INV_X1 U603 ( .A(n522), .ZN(n474) );
  XNOR2_X1 U604 ( .A(n474), .B(n509), .ZN(n738) );
  XNOR2_X1 U605 ( .A(n475), .B(n738), .ZN(n712) );
  NOR2_X1 U606 ( .A1(G902), .A2(n712), .ZN(n476) );
  XNOR2_X1 U607 ( .A(n477), .B(n476), .ZN(n564) );
  NAND2_X1 U608 ( .A1(n566), .A2(n564), .ZN(n478) );
  XNOR2_X1 U609 ( .A(n478), .B(KEYINPUT108), .ZN(n599) );
  NAND2_X1 U610 ( .A1(G214), .A2(n492), .ZN(n686) );
  XNOR2_X2 U611 ( .A(G116), .B(KEYINPUT71), .ZN(n481) );
  XNOR2_X1 U612 ( .A(G101), .B(G104), .ZN(n484) );
  NAND2_X1 U613 ( .A1(G224), .A2(n487), .ZN(n488) );
  XNOR2_X1 U614 ( .A(n489), .B(n506), .ZN(n490) );
  NAND2_X1 U615 ( .A1(n492), .A2(G210), .ZN(n493) );
  NAND2_X1 U616 ( .A1(G234), .A2(G237), .ZN(n497) );
  XNOR2_X1 U617 ( .A(n497), .B(KEYINPUT14), .ZN(n701) );
  NOR2_X1 U618 ( .A1(G902), .A2(n487), .ZN(n499) );
  NOR2_X1 U619 ( .A1(G953), .A2(G952), .ZN(n498) );
  NOR2_X1 U620 ( .A1(n499), .A2(n498), .ZN(n500) );
  AND2_X1 U621 ( .A1(n701), .A2(n500), .ZN(n577) );
  NAND2_X1 U622 ( .A1(G898), .A2(G953), .ZN(n501) );
  AND2_X1 U623 ( .A1(n577), .A2(n501), .ZN(n502) );
  NAND2_X1 U624 ( .A1(n594), .A2(n502), .ZN(n505) );
  XNOR2_X1 U625 ( .A(KEYINPUT0), .B(KEYINPUT66), .ZN(n503) );
  XNOR2_X1 U626 ( .A(n503), .B(KEYINPUT92), .ZN(n504) );
  XNOR2_X1 U627 ( .A(n506), .B(G137), .ZN(n508) );
  XOR2_X1 U628 ( .A(n509), .B(KEYINPUT94), .Z(n511) );
  NAND2_X1 U629 ( .A1(G227), .A2(n487), .ZN(n510) );
  XNOR2_X1 U630 ( .A(n511), .B(n510), .ZN(n512) );
  NOR2_X1 U631 ( .A1(n708), .A2(G902), .ZN(n515) );
  XOR2_X1 U632 ( .A(KEYINPUT96), .B(KEYINPUT21), .Z(n518) );
  XOR2_X1 U633 ( .A(KEYINPUT20), .B(KEYINPUT95), .Z(n516) );
  NAND2_X1 U634 ( .A1(n523), .A2(G221), .ZN(n517) );
  NAND2_X1 U635 ( .A1(G221), .A2(n519), .ZN(n521) );
  NAND2_X1 U636 ( .A1(n523), .A2(G217), .ZN(n524) );
  NAND2_X1 U637 ( .A1(n676), .A2(n542), .ZN(n673) );
  NOR2_X1 U638 ( .A1(n674), .A2(n673), .ZN(n558) );
  NAND2_X1 U639 ( .A1(n525), .A2(G210), .ZN(n526) );
  XNOR2_X1 U640 ( .A(n527), .B(n526), .ZN(n531) );
  INV_X1 U641 ( .A(G472), .ZN(n534) );
  NAND2_X1 U642 ( .A1(n354), .A2(n696), .ZN(n536) );
  XNOR2_X1 U643 ( .A(n536), .B(n363), .ZN(n537) );
  INV_X1 U644 ( .A(n542), .ZN(n580) );
  INV_X1 U645 ( .A(n674), .ZN(n617) );
  NAND2_X1 U646 ( .A1(n580), .A2(n570), .ZN(n544) );
  NOR2_X2 U647 ( .A1(n679), .A2(n544), .ZN(n646) );
  XNOR2_X1 U648 ( .A(n608), .B(KEYINPUT82), .ZN(n547) );
  NOR2_X1 U649 ( .A1(n674), .A2(n542), .ZN(n545) );
  XNOR2_X1 U650 ( .A(n545), .B(KEYINPUT107), .ZN(n546) );
  NOR2_X1 U651 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U652 ( .A(n548), .B(KEYINPUT81), .ZN(n549) );
  INV_X1 U653 ( .A(KEYINPUT91), .ZN(n552) );
  NAND2_X1 U654 ( .A1(n552), .A2(n748), .ZN(n554) );
  NOR2_X1 U655 ( .A1(n679), .A2(n673), .ZN(n556) );
  NAND2_X1 U656 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U657 ( .A1(n679), .A2(n558), .ZN(n682) );
  NOR2_X1 U658 ( .A1(n559), .A2(n682), .ZN(n562) );
  INV_X1 U659 ( .A(KEYINPUT31), .ZN(n560) );
  XNOR2_X1 U660 ( .A(n563), .B(KEYINPUT101), .ZN(n568) );
  INV_X1 U661 ( .A(n564), .ZN(n565) );
  AND2_X1 U662 ( .A1(n566), .A2(n565), .ZN(n658) );
  INV_X1 U663 ( .A(n691), .ZN(n567) );
  NAND2_X1 U664 ( .A1(n568), .A2(n567), .ZN(n571) );
  NOR2_X1 U665 ( .A1(n608), .A2(n580), .ZN(n569) );
  NAND2_X1 U666 ( .A1(n570), .A2(n569), .ZN(n638) );
  NAND2_X1 U667 ( .A1(n748), .A2(KEYINPUT44), .ZN(n572) );
  NAND2_X1 U668 ( .A1(n572), .A2(KEYINPUT91), .ZN(n573) );
  XOR2_X1 U669 ( .A(KEYINPUT45), .B(KEYINPUT64), .Z(n574) );
  XNOR2_X2 U670 ( .A(n575), .B(n574), .ZN(n727) );
  NAND2_X1 U671 ( .A1(G953), .A2(G900), .ZN(n576) );
  NAND2_X1 U672 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U673 ( .A(KEYINPUT84), .B(n578), .Z(n579) );
  NAND2_X1 U674 ( .A1(n676), .A2(n579), .ZN(n588) );
  INV_X1 U675 ( .A(KEYINPUT41), .ZN(n587) );
  NOR2_X1 U676 ( .A1(n542), .A2(n588), .ZN(n607) );
  AND2_X1 U677 ( .A1(n607), .A2(n679), .ZN(n589) );
  XOR2_X1 U678 ( .A(KEYINPUT28), .B(n589), .Z(n590) );
  NOR2_X1 U679 ( .A1(n691), .A2(KEYINPUT75), .ZN(n595) );
  NAND2_X1 U680 ( .A1(n594), .A2(n593), .ZN(n602) );
  NAND2_X1 U681 ( .A1(n595), .A2(n650), .ZN(n596) );
  NAND2_X1 U682 ( .A1(n596), .A2(KEYINPUT47), .ZN(n606) );
  OR2_X1 U683 ( .A1(n355), .A2(n597), .ZN(n598) );
  NOR2_X1 U684 ( .A1(n599), .A2(n598), .ZN(n649) );
  XNOR2_X1 U685 ( .A(n691), .B(KEYINPUT75), .ZN(n601) );
  INV_X1 U686 ( .A(KEYINPUT47), .ZN(n600) );
  NAND2_X1 U687 ( .A1(n601), .A2(n600), .ZN(n603) );
  NOR2_X1 U688 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U689 ( .A1(n649), .A2(n604), .ZN(n605) );
  INV_X1 U690 ( .A(n654), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U692 ( .A(n612), .B(KEYINPUT36), .ZN(n613) );
  NAND2_X1 U693 ( .A1(n613), .A2(n617), .ZN(n662) );
  NOR2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n619) );
  XNOR2_X1 U695 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n618) );
  XNOR2_X1 U696 ( .A(n619), .B(n618), .ZN(n620) );
  NOR2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U698 ( .A(KEYINPUT111), .B(n622), .Z(n747) );
  XNOR2_X1 U699 ( .A(n625), .B(KEYINPUT89), .ZN(n626) );
  NAND2_X1 U700 ( .A1(n626), .A2(KEYINPUT2), .ZN(n627) );
  NOR2_X1 U701 ( .A1(n747), .A2(n628), .ZN(n632) );
  NAND2_X1 U702 ( .A1(KEYINPUT2), .A2(n663), .ZN(n629) );
  XOR2_X1 U703 ( .A(KEYINPUT85), .B(n629), .Z(n630) );
  NOR2_X1 U704 ( .A1(n727), .A2(n630), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n632), .A2(n631), .ZN(n670) );
  NAND2_X1 U706 ( .A1(n713), .A2(G472), .ZN(n637) );
  XOR2_X1 U707 ( .A(KEYINPUT115), .B(KEYINPUT62), .Z(n635) );
  XOR2_X1 U708 ( .A(n633), .B(KEYINPUT114), .Z(n634) );
  XNOR2_X1 U709 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U710 ( .A(G101), .B(n638), .ZN(G3) );
  XNOR2_X1 U711 ( .A(G104), .B(KEYINPUT116), .ZN(n640) );
  NAND2_X1 U712 ( .A1(n654), .A2(n641), .ZN(n639) );
  XNOR2_X1 U713 ( .A(n640), .B(n639), .ZN(G6) );
  XOR2_X1 U714 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n643) );
  NAND2_X1 U715 ( .A1(n641), .A2(n658), .ZN(n642) );
  XNOR2_X1 U716 ( .A(n643), .B(n642), .ZN(n645) );
  XOR2_X1 U717 ( .A(G107), .B(KEYINPUT117), .Z(n644) );
  XNOR2_X1 U718 ( .A(n645), .B(n644), .ZN(G9) );
  XOR2_X1 U719 ( .A(n646), .B(G110), .Z(G12) );
  XOR2_X1 U720 ( .A(G128), .B(KEYINPUT29), .Z(n648) );
  NAND2_X1 U721 ( .A1(n650), .A2(n658), .ZN(n647) );
  XNOR2_X1 U722 ( .A(n648), .B(n647), .ZN(G30) );
  XOR2_X1 U723 ( .A(G143), .B(n649), .Z(G45) );
  XOR2_X1 U724 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n652) );
  NAND2_X1 U725 ( .A1(n650), .A2(n654), .ZN(n651) );
  XNOR2_X1 U726 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U727 ( .A(G146), .B(n653), .ZN(G48) );
  NAND2_X1 U728 ( .A1(n657), .A2(n654), .ZN(n655) );
  XNOR2_X1 U729 ( .A(n655), .B(KEYINPUT120), .ZN(n656) );
  XNOR2_X1 U730 ( .A(G113), .B(n656), .ZN(G15) );
  XOR2_X1 U731 ( .A(G116), .B(KEYINPUT121), .Z(n660) );
  NAND2_X1 U732 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U733 ( .A(n660), .B(n659), .ZN(G18) );
  XOR2_X1 U734 ( .A(G125), .B(KEYINPUT37), .Z(n661) );
  XNOR2_X1 U735 ( .A(n662), .B(n661), .ZN(G27) );
  XNOR2_X1 U736 ( .A(G134), .B(n663), .ZN(G36) );
  NAND2_X1 U737 ( .A1(n696), .A2(n664), .ZN(n672) );
  INV_X1 U738 ( .A(KEYINPUT2), .ZN(n666) );
  NAND2_X1 U739 ( .A1(n356), .A2(n666), .ZN(n665) );
  XNOR2_X1 U740 ( .A(n665), .B(KEYINPUT88), .ZN(n668) );
  NAND2_X1 U741 ( .A1(n727), .A2(n666), .ZN(n667) );
  NAND2_X1 U742 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U743 ( .A(KEYINPUT52), .B(KEYINPUT123), .ZN(n700) );
  NAND2_X1 U744 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U745 ( .A(n675), .B(KEYINPUT50), .ZN(n681) );
  NOR2_X1 U746 ( .A1(n542), .A2(n676), .ZN(n677) );
  XOR2_X1 U747 ( .A(KEYINPUT49), .B(n677), .Z(n678) );
  NOR2_X1 U748 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U749 ( .A1(n681), .A2(n680), .ZN(n683) );
  NAND2_X1 U750 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U751 ( .A(KEYINPUT51), .B(n684), .Z(n685) );
  NAND2_X1 U752 ( .A1(n664), .A2(n685), .ZN(n698) );
  NOR2_X1 U753 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U754 ( .A1(n689), .A2(n688), .ZN(n694) );
  NOR2_X1 U755 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U756 ( .A(KEYINPUT122), .B(n692), .ZN(n693) );
  OR2_X1 U757 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U758 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U759 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U760 ( .A(n700), .B(n699), .ZN(n703) );
  NAND2_X1 U761 ( .A1(n701), .A2(G952), .ZN(n702) );
  NOR2_X1 U762 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U763 ( .A(KEYINPUT53), .B(n705), .Z(G75) );
  BUF_X2 U764 ( .A(n713), .Z(n719) );
  NAND2_X1 U765 ( .A1(n719), .A2(G469), .ZN(n710) );
  XOR2_X1 U766 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n707) );
  NOR2_X1 U767 ( .A1(n722), .A2(n711), .ZN(G54) );
  NAND2_X1 U768 ( .A1(n713), .A2(G475), .ZN(n714) );
  NAND2_X1 U769 ( .A1(G478), .A2(n719), .ZN(n715) );
  NAND2_X1 U770 ( .A1(G217), .A2(n719), .ZN(n720) );
  NAND2_X1 U771 ( .A1(G224), .A2(G953), .ZN(n723) );
  XNOR2_X1 U772 ( .A(n723), .B(KEYINPUT61), .ZN(n724) );
  XNOR2_X1 U773 ( .A(KEYINPUT124), .B(n724), .ZN(n725) );
  NAND2_X1 U774 ( .A1(n725), .A2(G898), .ZN(n726) );
  XNOR2_X1 U775 ( .A(KEYINPUT125), .B(n726), .ZN(n730) );
  NOR2_X1 U776 ( .A1(G953), .A2(n727), .ZN(n728) );
  XNOR2_X1 U777 ( .A(n728), .B(KEYINPUT126), .ZN(n729) );
  NOR2_X1 U778 ( .A1(n730), .A2(n729), .ZN(n737) );
  XNOR2_X1 U779 ( .A(n731), .B(n732), .ZN(n733) );
  XNOR2_X1 U780 ( .A(n733), .B(KEYINPUT127), .ZN(n735) );
  NOR2_X1 U781 ( .A1(G898), .A2(n487), .ZN(n734) );
  NOR2_X1 U782 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U783 ( .A(n737), .B(n736), .Z(G69) );
  XNOR2_X1 U784 ( .A(n739), .B(n738), .ZN(n743) );
  XNOR2_X1 U785 ( .A(G227), .B(n743), .ZN(n740) );
  NAND2_X1 U786 ( .A1(G900), .A2(n740), .ZN(n741) );
  NAND2_X1 U787 ( .A1(n741), .A2(G953), .ZN(n746) );
  XNOR2_X1 U788 ( .A(n743), .B(n356), .ZN(n744) );
  NAND2_X1 U789 ( .A1(n744), .A2(n487), .ZN(n745) );
  NAND2_X1 U790 ( .A1(n746), .A2(n745), .ZN(G72) );
  XOR2_X1 U791 ( .A(G140), .B(n747), .Z(G42) );
  XOR2_X1 U792 ( .A(G122), .B(n748), .Z(G24) );
  XOR2_X1 U793 ( .A(G137), .B(n749), .Z(G39) );
  XOR2_X1 U794 ( .A(n750), .B(G131), .Z(G33) );
  XOR2_X1 U795 ( .A(n751), .B(G119), .Z(G21) );
endmodule

