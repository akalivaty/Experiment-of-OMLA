//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 1 0 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  OR2_X1    g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  AOI21_X1  g035(.A(G2105), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT67), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n465), .A2(new_n462), .A3(G101), .A4(G2104), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n461), .A2(G137), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n468), .B1(new_n459), .B2(new_n460), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(G2105), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n473), .B(KEYINPUT68), .ZN(G160));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G112), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  AND2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n462), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n461), .A2(KEYINPUT69), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n485), .B1(new_n480), .B2(G2105), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AOI211_X1 g062(.A(new_n477), .B(new_n483), .C1(G136), .C2(new_n487), .ZN(G162));
  OAI211_X1 g063(.A(G126), .B(G2105), .C1(new_n478), .C2(new_n479), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n478), .B2(new_n479), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n495), .B(new_n498), .C1(new_n479), .C2(new_n478), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n493), .B1(new_n497), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(G651), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n503), .A2(new_n505), .B1(new_n502), .B2(G651), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(G50), .A3(G543), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(KEYINPUT71), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT5), .A3(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n503), .A2(new_n505), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n502), .A2(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n507), .B1(new_n508), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n519), .A2(new_n504), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n518), .A2(new_n520), .ZN(G166));
  AND2_X1   g096(.A1(G63), .A2(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n514), .A2(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n515), .A2(G543), .A3(new_n516), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  INV_X1    g103(.A(G89), .ZN(new_n529));
  OAI221_X1 g104(.A(new_n526), .B1(new_n527), .B2(new_n528), .C1(new_n529), .C2(new_n517), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  INV_X1    g106(.A(new_n517), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G90), .ZN(new_n533));
  INV_X1    g108(.A(new_n527), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G52), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n514), .A2(G64), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n533), .A2(new_n535), .A3(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  AOI22_X1  g116(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n504), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n532), .A2(G81), .ZN(new_n544));
  XOR2_X1   g119(.A(KEYINPUT72), .B(G43), .Z(new_n545));
  NAND2_X1  g120(.A1(new_n534), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g124(.A1(new_n543), .A2(new_n544), .A3(KEYINPUT73), .A4(new_n546), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n527), .B2(new_n558), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n506), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n506), .A2(G91), .A3(new_n514), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(new_n511), .B2(new_n513), .ZN(new_n563));
  AND2_X1   g138(.A1(G78), .A2(G543), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n559), .A2(new_n560), .A3(new_n561), .A4(new_n565), .ZN(G299));
  OAI221_X1 g141(.A(new_n507), .B1(new_n517), .B2(new_n508), .C1(new_n504), .C2(new_n519), .ZN(G303));
  NAND3_X1  g142(.A1(new_n506), .A2(G87), .A3(new_n514), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n515), .A2(G49), .A3(G543), .A4(new_n516), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  INV_X1    g146(.A(G61), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n572), .B1(new_n511), .B2(new_n513), .ZN(new_n573));
  AND2_X1   g148(.A1(G73), .A2(G543), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n506), .A2(G86), .A3(new_n514), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n506), .A2(G48), .A3(G543), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n579), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(new_n504), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  INV_X1    g161(.A(G47), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n517), .A2(new_n586), .B1(new_n527), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT75), .ZN(new_n589));
  AND2_X1   g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n588), .A2(new_n589), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n585), .B1(new_n590), .B2(new_n591), .ZN(G290));
  XNOR2_X1  g167(.A(KEYINPUT76), .B(KEYINPUT10), .ZN(new_n593));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n517), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n593), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n506), .A2(G92), .A3(new_n596), .A4(new_n514), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(new_n511), .B2(new_n513), .ZN(new_n599));
  AND2_X1   g174(.A1(G79), .A2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n506), .A2(G54), .A3(G543), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n595), .A2(new_n597), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G171), .B2(new_n604), .ZN(G284));
  OAI21_X1  g181(.A(new_n605), .B1(G171), .B2(new_n604), .ZN(G321));
  NAND2_X1  g182(.A1(G286), .A2(G868), .ZN(new_n608));
  INV_X1    g183(.A(G299), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(G297));
  OAI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(G280));
  INV_X1    g186(.A(new_n603), .ZN(new_n612));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(new_n551), .B2(G868), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT77), .Z(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g194(.A(KEYINPUT3), .B(G2104), .ZN(new_n620));
  INV_X1    g195(.A(G2104), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n621), .A2(G2105), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(G111), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n627), .A2(KEYINPUT78), .A3(G2105), .ZN(new_n628));
  AOI21_X1  g203(.A(KEYINPUT78), .B1(new_n627), .B2(G2105), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI22_X1  g206(.A1(new_n481), .A2(G123), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n484), .A2(new_n486), .ZN(new_n633));
  INV_X1    g208(.A(G135), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI22_X1  g210(.A1(new_n626), .A2(G2100), .B1(G2096), .B2(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(G2096), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n636), .B(new_n637), .C1(G2100), .C2(new_n626), .ZN(G156));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n646), .A2(new_n648), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT79), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n649), .A2(new_n654), .A3(new_n650), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G401));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT80), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2072), .B(G2078), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT81), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  NAND3_X1  g240(.A1(new_n662), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT18), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n664), .B(KEYINPUT17), .Z(new_n668));
  INV_X1    g243(.A(new_n665), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n662), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n667), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n669), .B1(new_n662), .B2(new_n664), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n672), .A2(KEYINPUT82), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(KEYINPUT82), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n673), .B(new_n674), .C1(new_n668), .C2(new_n661), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2096), .B(G2100), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n671), .A2(new_n675), .A3(new_n677), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n682), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n682), .B2(new_n688), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT83), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n694), .A2(new_n696), .ZN(new_n699));
  AND3_X1   g274(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n698), .B1(new_n697), .B2(new_n699), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(G229));
  NAND3_X1  g277(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT96), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT26), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n622), .A2(G105), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n481), .B2(G129), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n487), .A2(G141), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n708), .A2(KEYINPUT95), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(KEYINPUT95), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n705), .B(new_n707), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G29), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G32), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT27), .B(G1996), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n712), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT97), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n715), .B1(new_n712), .B2(new_n714), .ZN(new_n719));
  NAND2_X1  g294(.A1(G160), .A2(G29), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT84), .B(G29), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT24), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n722), .A2(G34), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(G34), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n721), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G2084), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G16), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G21), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G168), .B2(new_n729), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(G1966), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n729), .A2(G5), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G171), .B2(new_n729), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G1961), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n720), .A2(G2084), .A3(new_n725), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n728), .A2(new_n732), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT31), .B(G11), .Z(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT98), .B(G28), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(KEYINPUT30), .ZN(new_n741));
  AOI21_X1  g316(.A(G29), .B1(new_n740), .B2(KEYINPUT30), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n738), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n635), .B2(new_n721), .ZN(new_n744));
  NOR2_X1   g319(.A1(G164), .A2(new_n721), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G27), .B2(new_n721), .ZN(new_n746));
  INV_X1    g321(.A(G2078), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n744), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n731), .A2(G1966), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n748), .B(new_n749), .C1(new_n747), .C2(new_n746), .ZN(new_n750));
  NOR3_X1   g325(.A1(new_n719), .A2(new_n737), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(G115), .A2(G2104), .ZN(new_n752));
  INV_X1    g327(.A(G127), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n480), .B2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT94), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n462), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n755), .B2(new_n754), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n487), .A2(G139), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT25), .Z(new_n760));
  NAND3_X1  g335(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  MUX2_X1   g336(.A(G33), .B(new_n761), .S(G29), .Z(new_n762));
  OAI22_X1  g337(.A1(new_n762), .A2(G2072), .B1(new_n734), .B2(G1961), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G2072), .B2(new_n762), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n718), .A2(new_n751), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(KEYINPUT99), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT99), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n718), .A2(new_n751), .A3(new_n767), .A4(new_n764), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n721), .ZN(new_n770));
  NAND2_X1  g345(.A1(G162), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G35), .B2(new_n770), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT29), .ZN(new_n773));
  INV_X1    g348(.A(G2090), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n729), .A2(G20), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT23), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n609), .B2(new_n729), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT100), .ZN(new_n779));
  INV_X1    g354(.A(G1956), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n779), .A2(new_n780), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n775), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(KEYINPUT101), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(KEYINPUT101), .ZN(new_n785));
  INV_X1    g360(.A(G19), .ZN(new_n786));
  OR3_X1    g361(.A1(new_n786), .A2(KEYINPUT89), .A3(G16), .ZN(new_n787));
  OAI21_X1  g362(.A(KEYINPUT89), .B1(new_n786), .B2(G16), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n787), .B(new_n788), .C1(new_n551), .C2(new_n729), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT90), .B(G1341), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G1348), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n612), .A2(new_n729), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G4), .B2(new_n729), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n773), .A2(new_n774), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n721), .A2(G26), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n487), .A2(G140), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT91), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G116), .B2(new_n462), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n481), .A2(G128), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT92), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n801), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n798), .B1(new_n807), .B2(G29), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G2067), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n794), .A2(new_n792), .ZN(new_n810));
  AND4_X1   g385(.A1(new_n791), .A2(new_n795), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n769), .A2(new_n784), .A3(new_n785), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(G6), .A2(G16), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n582), .B2(G16), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT32), .B(G1981), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n814), .B(new_n815), .Z(new_n816));
  NAND2_X1  g391(.A1(G288), .A2(KEYINPUT86), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT86), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n568), .A2(new_n569), .A3(new_n570), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G16), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G16), .B2(G23), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT33), .B(G1976), .Z(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n729), .A2(G22), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(G166), .B2(new_n729), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G1971), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n825), .B2(new_n823), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n816), .A2(new_n826), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT34), .ZN(new_n832));
  MUX2_X1   g407(.A(G24), .B(G290), .S(G16), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G1986), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n770), .A2(G25), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n481), .A2(G119), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n462), .A2(G107), .ZN(new_n838));
  OAI21_X1  g413(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n839));
  INV_X1    g414(.A(G131), .ZN(new_n840));
  OAI221_X1 g415(.A(new_n837), .B1(new_n838), .B2(new_n839), .C1(new_n633), .C2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT85), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n836), .B1(new_n842), .B2(new_n721), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT35), .B(G1991), .Z(new_n844));
  AND2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n834), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT87), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT34), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n816), .A2(new_n849), .A3(new_n826), .A4(new_n830), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n848), .B1(new_n847), .B2(new_n850), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n832), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n854), .A2(KEYINPUT88), .A3(KEYINPUT36), .ZN(new_n855));
  NAND2_X1  g430(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n832), .B(new_n856), .C1(new_n852), .C2(new_n853), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n812), .B1(new_n855), .B2(new_n857), .ZN(G311));
  INV_X1    g433(.A(new_n812), .ZN(new_n859));
  INV_X1    g434(.A(new_n853), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n851), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n856), .B1(new_n861), .B2(new_n832), .ZN(new_n862));
  INV_X1    g437(.A(new_n857), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(G150));
  AOI22_X1  g439(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n865), .A2(new_n504), .ZN(new_n866));
  XOR2_X1   g441(.A(KEYINPUT102), .B(G93), .Z(new_n867));
  NAND3_X1  g442(.A1(new_n506), .A2(new_n514), .A3(new_n867), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n515), .A2(G55), .A3(G543), .A4(new_n516), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n868), .A2(KEYINPUT103), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT103), .B1(new_n868), .B2(new_n869), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n866), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g449(.A(KEYINPUT104), .B(new_n866), .C1(new_n870), .C2(new_n871), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n547), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n549), .A2(new_n550), .A3(new_n872), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n603), .A2(new_n613), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT38), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n878), .B(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT39), .ZN(new_n882));
  AOI21_X1  g457(.A(G860), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(new_n882), .B2(new_n881), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT105), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n874), .A2(new_n875), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(G860), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT106), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT37), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n885), .A2(new_n889), .ZN(G145));
  INV_X1    g465(.A(KEYINPUT40), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n807), .A2(new_n711), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n807), .A2(new_n711), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n487), .A2(G142), .ZN(new_n895));
  OAI21_X1  g470(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n896));
  INV_X1    g471(.A(G118), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n896), .B1(new_n897), .B2(G2105), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n898), .B1(new_n481), .B2(G130), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n895), .A2(new_n899), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n892), .A2(new_n901), .A3(new_n893), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n841), .B(KEYINPUT108), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n624), .ZN(new_n905));
  XNOR2_X1  g480(.A(G164), .B(KEYINPUT107), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(new_n761), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n907), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n903), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(G160), .B(new_n635), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(G162), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n900), .A2(new_n908), .A3(new_n902), .A4(new_n909), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G37), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n913), .B1(new_n911), .B2(new_n914), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n891), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n918), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n920), .A2(KEYINPUT40), .A3(new_n916), .A4(new_n915), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n919), .A2(new_n921), .ZN(G395));
  XNOR2_X1  g497(.A(new_n878), .B(new_n615), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n612), .A2(G299), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n609), .A2(new_n603), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n609), .A2(new_n930), .A3(new_n603), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n924), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n930), .B1(new_n609), .B2(new_n603), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT110), .B1(new_n926), .B2(new_n929), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n924), .A2(new_n925), .A3(new_n936), .A4(KEYINPUT41), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n923), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n928), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT42), .ZN(new_n941));
  NAND2_X1  g516(.A1(G290), .A2(G166), .ZN(new_n942));
  OAI211_X1 g517(.A(G303), .B(new_n585), .C1(new_n590), .C2(new_n591), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n582), .A2(new_n821), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n820), .A2(new_n580), .A3(new_n581), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n944), .A2(new_n947), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n928), .A2(new_n951), .A3(new_n939), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n941), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n950), .B1(new_n941), .B2(new_n952), .ZN(new_n954));
  OAI21_X1  g529(.A(G868), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n886), .A2(new_n604), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(G295));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n956), .ZN(G331));
  NAND2_X1  g533(.A1(new_n925), .A2(KEYINPUT109), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n959), .A2(KEYINPUT41), .A3(new_n931), .A4(new_n924), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n931), .A2(new_n924), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n963), .A2(KEYINPUT111), .A3(KEYINPUT41), .A4(new_n959), .ZN(new_n964));
  XNOR2_X1  g539(.A(G301), .B(G286), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n876), .A2(new_n965), .A3(new_n877), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n965), .B1(new_n876), .B2(new_n877), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n962), .B(new_n964), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n965), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n878), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n876), .A2(new_n965), .A3(new_n877), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n929), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n968), .B1(new_n972), .B2(new_n927), .ZN(new_n973));
  INV_X1    g548(.A(new_n950), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n938), .B1(new_n966), .B2(new_n967), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n970), .A2(new_n926), .A3(new_n971), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n950), .A3(new_n978), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n975), .A2(new_n976), .A3(new_n916), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT112), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n979), .A2(new_n916), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n982), .A2(new_n983), .A3(new_n976), .A4(new_n975), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n979), .A2(new_n916), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n950), .B1(new_n977), .B2(new_n978), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT43), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n981), .A2(new_n984), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n982), .A2(KEYINPUT43), .A3(new_n975), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n976), .B1(new_n985), .B2(new_n986), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT44), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n990), .A2(new_n994), .ZN(G397));
  NAND2_X1  g570(.A1(new_n497), .A2(new_n499), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n489), .A2(new_n492), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n998), .A2(KEYINPUT45), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n464), .A2(new_n466), .ZN(new_n1000));
  OAI211_X1 g575(.A(G137), .B(new_n462), .C1(new_n478), .C2(new_n479), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(G125), .B1(new_n478), .B2(new_n479), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n462), .B1(new_n1003), .B2(new_n470), .ZN(new_n1004));
  INV_X1    g579(.A(G40), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n999), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n807), .B(G2067), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1008), .B1(new_n1009), .B2(new_n711), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1007), .A2(G1996), .ZN(new_n1011));
  XOR2_X1   g586(.A(new_n1011), .B(KEYINPUT46), .Z(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1013), .A2(KEYINPUT47), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1013), .A2(KEYINPUT47), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n711), .B(G1996), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1008), .B1(new_n1009), .B2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n841), .B(new_n844), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1017), .B1(new_n1007), .B2(new_n1018), .ZN(new_n1019));
  NOR3_X1   g594(.A1(G290), .A2(new_n1007), .A3(G1986), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(KEYINPUT48), .ZN(new_n1021));
  OAI22_X1  g596(.A1(new_n1014), .A2(new_n1015), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n807), .A2(G2067), .ZN(new_n1023));
  INV_X1    g598(.A(new_n844), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n842), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1023), .B1(new_n1017), .B2(new_n1025), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1026), .A2(KEYINPUT126), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1007), .B1(new_n1026), .B2(KEYINPUT126), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1022), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n998), .B2(KEYINPUT45), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n467), .A2(new_n472), .A3(G40), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(new_n998), .B2(KEYINPUT45), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n1034));
  OAI211_X1 g609(.A(KEYINPUT113), .B(new_n1034), .C1(G164), .C2(G1384), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1031), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1971), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1006), .B1(G164), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n1042));
  INV_X1    g617(.A(new_n499), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n498), .B1(new_n620), .B2(new_n495), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n489), .B(new_n492), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1384), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1042), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1041), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n774), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1038), .A2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT55), .B(G8), .C1(new_n518), .C2(new_n520), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT114), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n1053));
  INV_X1    g628(.A(G8), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1053), .B1(G166), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT114), .ZN(new_n1056));
  NAND4_X1  g631(.A1(G303), .A2(new_n1056), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1052), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1050), .A2(G8), .A3(new_n1058), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1052), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1036), .A2(new_n1037), .B1(new_n1048), .B2(new_n774), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(new_n1061), .B2(new_n1054), .ZN(new_n1062));
  AND2_X1   g637(.A1(KEYINPUT115), .A2(G86), .ZN(new_n1063));
  NOR2_X1   g638(.A1(KEYINPUT115), .A2(G86), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n514), .A2(new_n515), .A3(new_n516), .A4(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n575), .A2(new_n577), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(G1981), .ZN(new_n1068));
  INV_X1    g643(.A(G1981), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n576), .A2(new_n575), .A3(new_n577), .A4(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT49), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1054), .B1(new_n998), .B2(new_n1006), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1068), .A2(KEYINPUT49), .A3(new_n1070), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n817), .A2(G1976), .A3(new_n819), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n1074), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT52), .ZN(new_n1079));
  INV_X1    g654(.A(G1976), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT52), .B1(G288), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1077), .A2(new_n1074), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1076), .A2(new_n1079), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1059), .A2(new_n1062), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1031), .A2(new_n1033), .A3(new_n747), .A4(new_n1035), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1032), .B1(new_n1045), .B2(new_n1039), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1091));
  AOI21_X1  g666(.A(G1961), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT124), .B1(new_n999), .B2(new_n1032), .ZN(new_n1094));
  AOI211_X1 g669(.A(new_n1088), .B(G2078), .C1(new_n998), .C2(KEYINPUT45), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1034), .B1(G164), .B2(G1384), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(new_n1097), .A3(new_n1006), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1094), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1099));
  AND4_X1   g674(.A1(G301), .A2(new_n1089), .A3(new_n1093), .A4(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1092), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1095), .A2(new_n1096), .A3(new_n1006), .ZN(new_n1102));
  AOI21_X1  g677(.A(G301), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1086), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1089), .A2(new_n1099), .A3(new_n1093), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(G171), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1101), .A2(G301), .A3(new_n1102), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(KEYINPUT54), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G1966), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1045), .A2(KEYINPUT45), .A3(new_n1046), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n1006), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1109), .B1(new_n1111), .B2(new_n999), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT119), .B(G2084), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1090), .A2(new_n1091), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1054), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(G286), .A2(G8), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT51), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1090), .A2(new_n1091), .A3(new_n1113), .ZN(new_n1120));
  AOI21_X1  g695(.A(G1966), .B1(new_n1033), .B2(new_n1096), .ZN(new_n1121));
  OAI21_X1  g696(.A(G8), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1116), .B(KEYINPUT123), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1117), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g699(.A(G8), .B(G286), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1119), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AND4_X1   g701(.A1(new_n1085), .A2(new_n1104), .A3(new_n1108), .A4(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT56), .B(G2072), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1031), .A2(new_n1033), .A3(new_n1035), .A4(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n1130));
  NAND2_X1  g705(.A1(G299), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT57), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(G299), .A2(new_n1130), .A3(KEYINPUT57), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n780), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1129), .A2(new_n1133), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(G1348), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n1138));
  INV_X1    g713(.A(G2067), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n998), .A2(new_n1006), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1137), .A2(new_n1138), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n792), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT122), .B1(new_n1143), .B2(new_n1140), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n1142), .A2(new_n1144), .A3(new_n603), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1129), .A2(new_n1135), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1136), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT60), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1138), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1143), .A2(KEYINPUT122), .A3(new_n1140), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1148), .A2(new_n612), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1136), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1154), .B1(new_n1155), .B2(new_n1146), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1146), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1157), .A2(new_n1136), .A3(KEYINPUT61), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1153), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n998), .A2(new_n1006), .ZN(new_n1160));
  XOR2_X1   g735(.A(KEYINPUT58), .B(G1341), .Z(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1162), .B1(new_n1036), .B2(G1996), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n551), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT59), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1163), .A2(KEYINPUT59), .A3(new_n551), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1166), .B(new_n1167), .C1(new_n612), .C2(new_n1148), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1147), .B1(new_n1159), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1127), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT63), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1059), .A2(new_n1062), .A3(new_n1084), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1115), .A2(G168), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1061), .A2(new_n1060), .A3(new_n1054), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1175), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT116), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1083), .A2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1076), .A2(new_n1079), .A3(KEYINPUT116), .A4(new_n1082), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1050), .A2(G8), .ZN(new_n1180));
  AOI22_X1  g755(.A1(new_n1178), .A2(new_n1179), .B1(new_n1180), .B2(new_n1060), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1176), .B1(new_n1181), .B2(KEYINPUT120), .ZN(new_n1182));
  AOI21_X1  g757(.A(KEYINPUT49), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1160), .A2(G8), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1185), .A2(new_n1075), .B1(KEYINPUT52), .B2(new_n1078), .ZN(new_n1186));
  AOI21_X1  g761(.A(KEYINPUT116), .B1(new_n1186), .B2(new_n1082), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1179), .ZN(new_n1188));
  OAI211_X1 g763(.A(KEYINPUT120), .B(new_n1062), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1174), .B1(new_n1182), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1175), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1192));
  NOR2_X1   g767(.A1(G288), .A2(G1976), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1193), .B(KEYINPUT118), .ZN(new_n1194));
  AND2_X1   g769(.A1(new_n1076), .A2(new_n1194), .ZN(new_n1195));
  XOR2_X1   g770(.A(new_n1070), .B(KEYINPUT117), .Z(new_n1196));
  OAI21_X1  g771(.A(new_n1074), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1192), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT123), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1116), .B(new_n1199), .ZN(new_n1200));
  OAI211_X1 g775(.A(new_n1125), .B(KEYINPUT51), .C1(new_n1115), .C2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1122), .A2(new_n1117), .A3(new_n1116), .ZN(new_n1202));
  AOI21_X1  g777(.A(KEYINPUT62), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND4_X1  g778(.A1(new_n1059), .A2(new_n1103), .A3(new_n1062), .A4(new_n1084), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1126), .A2(KEYINPUT62), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1198), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1170), .A2(new_n1191), .A3(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT125), .ZN(new_n1209));
  XNOR2_X1  g784(.A(G290), .B(G1986), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1019), .B1(new_n1008), .B2(new_n1210), .ZN(new_n1211));
  AND3_X1   g786(.A1(new_n1208), .A2(new_n1209), .A3(new_n1211), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1209), .B1(new_n1208), .B2(new_n1211), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1029), .B1(new_n1212), .B2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g789(.A1(new_n920), .A2(new_n916), .A3(new_n915), .ZN(new_n1216));
  AND3_X1   g790(.A1(new_n678), .A2(G319), .A3(new_n679), .ZN(new_n1217));
  NAND2_X1  g791(.A1(new_n1217), .A2(new_n658), .ZN(new_n1218));
  INV_X1    g792(.A(KEYINPUT127), .ZN(new_n1219));
  NAND2_X1  g793(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g794(.A1(new_n1217), .A2(KEYINPUT127), .A3(new_n658), .ZN(new_n1221));
  AOI21_X1  g795(.A(G229), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  AND3_X1   g796(.A1(new_n988), .A2(new_n1216), .A3(new_n1222), .ZN(G308));
  NAND3_X1  g797(.A1(new_n988), .A2(new_n1216), .A3(new_n1222), .ZN(G225));
endmodule


