

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U554 ( .A(n524), .B(KEYINPUT17), .ZN(n525) );
  BUF_X2 U555 ( .A(n902), .Z(n521) );
  NOR2_X1 U556 ( .A1(G2104), .A2(n529), .ZN(n902) );
  INV_X1 U557 ( .A(KEYINPUT103), .ZN(n768) );
  INV_X1 U558 ( .A(KEYINPUT23), .ZN(n522) );
  INV_X1 U559 ( .A(KEYINPUT97), .ZN(n690) );
  NOR2_X1 U560 ( .A1(n692), .A2(n927), .ZN(n693) );
  INV_X1 U561 ( .A(KEYINPUT100), .ZN(n708) );
  NOR2_X1 U562 ( .A1(G164), .A2(G1384), .ZN(n684) );
  INV_X1 U563 ( .A(n945), .ZN(n761) );
  XNOR2_X1 U564 ( .A(KEYINPUT87), .B(n682), .ZN(n781) );
  INV_X1 U565 ( .A(KEYINPUT66), .ZN(n524) );
  INV_X1 U566 ( .A(KEYINPUT104), .ZN(n778) );
  INV_X1 U567 ( .A(G2105), .ZN(n529) );
  AND2_X2 U568 ( .A1(n529), .A2(G2104), .ZN(n899) );
  XNOR2_X1 U569 ( .A(n523), .B(n522), .ZN(n528) );
  NAND2_X1 U570 ( .A1(G101), .A2(n899), .ZN(n523) );
  NOR2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XNOR2_X2 U572 ( .A(n526), .B(n525), .ZN(n604) );
  NAND2_X1 U573 ( .A1(G137), .A2(n604), .ZN(n527) );
  NAND2_X1 U574 ( .A1(n528), .A2(n527), .ZN(n533) );
  NAND2_X1 U575 ( .A1(G125), .A2(n521), .ZN(n531) );
  AND2_X1 U576 ( .A1(G2104), .A2(G2105), .ZN(n904) );
  NAND2_X1 U577 ( .A1(G113), .A2(n904), .ZN(n530) );
  NAND2_X1 U578 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X2 U579 ( .A1(n533), .A2(n532), .ZN(G160) );
  INV_X1 U580 ( .A(G651), .ZN(n539) );
  NOR2_X1 U581 ( .A1(G543), .A2(n539), .ZN(n534) );
  XOR2_X1 U582 ( .A(KEYINPUT1), .B(n534), .Z(n643) );
  NAND2_X1 U583 ( .A1(G64), .A2(n643), .ZN(n538) );
  XNOR2_X1 U584 ( .A(G543), .B(KEYINPUT0), .ZN(n535) );
  XNOR2_X1 U585 ( .A(n535), .B(KEYINPUT67), .ZN(n621) );
  NOR2_X1 U586 ( .A1(G651), .A2(n621), .ZN(n536) );
  XOR2_X2 U587 ( .A(KEYINPUT65), .B(n536), .Z(n650) );
  NAND2_X1 U588 ( .A1(G52), .A2(n650), .ZN(n537) );
  NAND2_X1 U589 ( .A1(n538), .A2(n537), .ZN(n545) );
  NOR2_X1 U590 ( .A1(n621), .A2(n539), .ZN(n646) );
  NAND2_X1 U591 ( .A1(n646), .A2(G77), .ZN(n540) );
  XNOR2_X1 U592 ( .A(n540), .B(KEYINPUT70), .ZN(n542) );
  NOR2_X1 U593 ( .A1(G651), .A2(G543), .ZN(n642) );
  NAND2_X1 U594 ( .A1(G90), .A2(n642), .ZN(n541) );
  NAND2_X1 U595 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U596 ( .A(KEYINPUT9), .B(n543), .Z(n544) );
  NOR2_X1 U597 ( .A1(n545), .A2(n544), .ZN(G171) );
  INV_X1 U598 ( .A(G171), .ZN(G301) );
  AND2_X1 U599 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U600 ( .A1(G126), .A2(n521), .ZN(n547) );
  NAND2_X1 U601 ( .A1(G114), .A2(n904), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U603 ( .A(KEYINPUT86), .B(n548), .ZN(n552) );
  NAND2_X1 U604 ( .A1(n899), .A2(G102), .ZN(n550) );
  NAND2_X1 U605 ( .A1(G138), .A2(n604), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U607 ( .A1(n552), .A2(n551), .ZN(G164) );
  INV_X1 U608 ( .A(G57), .ZN(G237) );
  INV_X1 U609 ( .A(G132), .ZN(G219) );
  INV_X1 U610 ( .A(G82), .ZN(G220) );
  NAND2_X1 U611 ( .A1(n642), .A2(G89), .ZN(n553) );
  XNOR2_X1 U612 ( .A(n553), .B(KEYINPUT4), .ZN(n555) );
  NAND2_X1 U613 ( .A1(G76), .A2(n646), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U615 ( .A(n556), .B(KEYINPUT5), .ZN(n561) );
  NAND2_X1 U616 ( .A1(G63), .A2(n643), .ZN(n558) );
  NAND2_X1 U617 ( .A1(G51), .A2(n650), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U619 ( .A(KEYINPUT6), .B(n559), .Z(n560) );
  NAND2_X1 U620 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U621 ( .A(n562), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U622 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U623 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n565) );
  NAND2_X1 U624 ( .A1(G7), .A2(G661), .ZN(n563) );
  XOR2_X1 U625 ( .A(n563), .B(KEYINPUT10), .Z(n835) );
  NAND2_X1 U626 ( .A1(G567), .A2(n835), .ZN(n564) );
  XNOR2_X1 U627 ( .A(n565), .B(n564), .ZN(G234) );
  NAND2_X1 U628 ( .A1(n643), .A2(G56), .ZN(n566) );
  XOR2_X1 U629 ( .A(KEYINPUT14), .B(n566), .Z(n574) );
  NAND2_X1 U630 ( .A1(G68), .A2(n646), .ZN(n570) );
  XOR2_X1 U631 ( .A(KEYINPUT73), .B(KEYINPUT12), .Z(n568) );
  NAND2_X1 U632 ( .A1(G81), .A2(n642), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U635 ( .A(n571), .B(KEYINPUT74), .ZN(n572) );
  XOR2_X1 U636 ( .A(KEYINPUT13), .B(n572), .Z(n573) );
  NOR2_X1 U637 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U638 ( .A1(n650), .A2(G43), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n927) );
  XNOR2_X1 U640 ( .A(G860), .B(KEYINPUT75), .ZN(n595) );
  OR2_X1 U641 ( .A1(n927), .A2(n595), .ZN(G153) );
  NAND2_X1 U642 ( .A1(G868), .A2(G301), .ZN(n585) );
  NAND2_X1 U643 ( .A1(G79), .A2(n646), .ZN(n578) );
  NAND2_X1 U644 ( .A1(G66), .A2(n643), .ZN(n577) );
  NAND2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n582) );
  NAND2_X1 U646 ( .A1(G92), .A2(n642), .ZN(n580) );
  NAND2_X1 U647 ( .A1(G54), .A2(n650), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U649 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U650 ( .A(KEYINPUT15), .B(n583), .Z(n926) );
  OR2_X1 U651 ( .A1(n926), .A2(G868), .ZN(n584) );
  NAND2_X1 U652 ( .A1(n585), .A2(n584), .ZN(G284) );
  NAND2_X1 U653 ( .A1(G78), .A2(n646), .ZN(n587) );
  NAND2_X1 U654 ( .A1(G65), .A2(n643), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U656 ( .A1(G91), .A2(n642), .ZN(n588) );
  XNOR2_X1 U657 ( .A(KEYINPUT71), .B(n588), .ZN(n589) );
  NOR2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U659 ( .A1(n650), .A2(G53), .ZN(n591) );
  NAND2_X1 U660 ( .A1(n592), .A2(n591), .ZN(G299) );
  INV_X1 U661 ( .A(G868), .ZN(n661) );
  NOR2_X1 U662 ( .A1(G286), .A2(n661), .ZN(n594) );
  NOR2_X1 U663 ( .A1(G868), .A2(G299), .ZN(n593) );
  NOR2_X1 U664 ( .A1(n594), .A2(n593), .ZN(G297) );
  NAND2_X1 U665 ( .A1(n595), .A2(G559), .ZN(n596) );
  NAND2_X1 U666 ( .A1(n596), .A2(n926), .ZN(n597) );
  XNOR2_X1 U667 ( .A(n597), .B(KEYINPUT16), .ZN(n598) );
  XNOR2_X1 U668 ( .A(KEYINPUT76), .B(n598), .ZN(G148) );
  NOR2_X1 U669 ( .A1(G868), .A2(n927), .ZN(n601) );
  NAND2_X1 U670 ( .A1(n926), .A2(G868), .ZN(n599) );
  NOR2_X1 U671 ( .A1(G559), .A2(n599), .ZN(n600) );
  NOR2_X1 U672 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U673 ( .A1(G123), .A2(n521), .ZN(n602) );
  XOR2_X1 U674 ( .A(KEYINPUT18), .B(n602), .Z(n603) );
  XNOR2_X1 U675 ( .A(n603), .B(KEYINPUT77), .ZN(n606) );
  NAND2_X1 U676 ( .A1(G135), .A2(n604), .ZN(n605) );
  NAND2_X1 U677 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U678 ( .A(KEYINPUT78), .B(n607), .ZN(n611) );
  NAND2_X1 U679 ( .A1(G111), .A2(n904), .ZN(n609) );
  NAND2_X1 U680 ( .A1(G99), .A2(n899), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U682 ( .A1(n611), .A2(n610), .ZN(n988) );
  XNOR2_X1 U683 ( .A(n988), .B(G2096), .ZN(n612) );
  INV_X1 U684 ( .A(G2100), .ZN(n857) );
  NAND2_X1 U685 ( .A1(n612), .A2(n857), .ZN(G156) );
  NAND2_X1 U686 ( .A1(G80), .A2(n646), .ZN(n614) );
  NAND2_X1 U687 ( .A1(G67), .A2(n643), .ZN(n613) );
  NAND2_X1 U688 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U689 ( .A1(G93), .A2(n642), .ZN(n616) );
  NAND2_X1 U690 ( .A1(G55), .A2(n650), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n617) );
  OR2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n662) );
  NAND2_X1 U693 ( .A1(G559), .A2(n926), .ZN(n619) );
  XNOR2_X1 U694 ( .A(n927), .B(n619), .ZN(n658) );
  NOR2_X1 U695 ( .A1(G860), .A2(n658), .ZN(n620) );
  XOR2_X1 U696 ( .A(n662), .B(n620), .Z(G145) );
  NAND2_X1 U697 ( .A1(G49), .A2(n650), .ZN(n623) );
  NAND2_X1 U698 ( .A1(G87), .A2(n621), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U700 ( .A1(n643), .A2(n624), .ZN(n626) );
  NAND2_X1 U701 ( .A1(G651), .A2(G74), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n626), .A2(n625), .ZN(G288) );
  NAND2_X1 U703 ( .A1(G88), .A2(n642), .ZN(n628) );
  NAND2_X1 U704 ( .A1(G62), .A2(n643), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U706 ( .A1(G75), .A2(n646), .ZN(n629) );
  XNOR2_X1 U707 ( .A(KEYINPUT79), .B(n629), .ZN(n630) );
  NOR2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n650), .A2(G50), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(G303) );
  NAND2_X1 U711 ( .A1(n643), .A2(G60), .ZN(n640) );
  NAND2_X1 U712 ( .A1(G72), .A2(n646), .ZN(n635) );
  NAND2_X1 U713 ( .A1(G85), .A2(n642), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U715 ( .A1(G47), .A2(n650), .ZN(n636) );
  XOR2_X1 U716 ( .A(KEYINPUT68), .B(n636), .Z(n637) );
  NOR2_X1 U717 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U719 ( .A(KEYINPUT69), .B(n641), .Z(G290) );
  NAND2_X1 U720 ( .A1(G86), .A2(n642), .ZN(n645) );
  NAND2_X1 U721 ( .A1(G61), .A2(n643), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(n649) );
  NAND2_X1 U723 ( .A1(n646), .A2(G73), .ZN(n647) );
  XOR2_X1 U724 ( .A(KEYINPUT2), .B(n647), .Z(n648) );
  NOR2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U726 ( .A1(n650), .A2(G48), .ZN(n651) );
  NAND2_X1 U727 ( .A1(n652), .A2(n651), .ZN(G305) );
  XNOR2_X1 U728 ( .A(KEYINPUT19), .B(G288), .ZN(n657) );
  XOR2_X1 U729 ( .A(G303), .B(G290), .Z(n653) );
  XNOR2_X1 U730 ( .A(n653), .B(G305), .ZN(n654) );
  XOR2_X1 U731 ( .A(n662), .B(n654), .Z(n655) );
  XNOR2_X1 U732 ( .A(n655), .B(G299), .ZN(n656) );
  XNOR2_X1 U733 ( .A(n657), .B(n656), .ZN(n915) );
  XOR2_X1 U734 ( .A(n658), .B(n915), .Z(n659) );
  XNOR2_X1 U735 ( .A(KEYINPUT80), .B(n659), .ZN(n660) );
  NOR2_X1 U736 ( .A1(n661), .A2(n660), .ZN(n664) );
  NOR2_X1 U737 ( .A1(G868), .A2(n662), .ZN(n663) );
  NOR2_X1 U738 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U739 ( .A1(G2078), .A2(G2084), .ZN(n665) );
  XNOR2_X1 U740 ( .A(n665), .B(KEYINPUT20), .ZN(n666) );
  XNOR2_X1 U741 ( .A(n666), .B(KEYINPUT81), .ZN(n667) );
  NAND2_X1 U742 ( .A1(n667), .A2(G2090), .ZN(n668) );
  XNOR2_X1 U743 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U744 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U745 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U746 ( .A1(G220), .A2(G219), .ZN(n670) );
  XOR2_X1 U747 ( .A(KEYINPUT22), .B(n670), .Z(n671) );
  NOR2_X1 U748 ( .A1(G218), .A2(n671), .ZN(n672) );
  NAND2_X1 U749 ( .A1(G96), .A2(n672), .ZN(n839) );
  NAND2_X1 U750 ( .A1(G2106), .A2(n839), .ZN(n673) );
  XNOR2_X1 U751 ( .A(n673), .B(KEYINPUT82), .ZN(n677) );
  NAND2_X1 U752 ( .A1(G69), .A2(G120), .ZN(n674) );
  NOR2_X1 U753 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U754 ( .A1(G108), .A2(n675), .ZN(n840) );
  NAND2_X1 U755 ( .A1(G567), .A2(n840), .ZN(n676) );
  NAND2_X1 U756 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U757 ( .A(KEYINPUT83), .B(n678), .Z(n925) );
  NAND2_X1 U758 ( .A1(G661), .A2(G483), .ZN(n679) );
  XNOR2_X1 U759 ( .A(KEYINPUT84), .B(n679), .ZN(n680) );
  NOR2_X1 U760 ( .A1(n925), .A2(n680), .ZN(n838) );
  NAND2_X1 U761 ( .A1(n838), .A2(G36), .ZN(n681) );
  XOR2_X1 U762 ( .A(KEYINPUT85), .B(n681), .Z(G176) );
  NAND2_X1 U763 ( .A1(G1976), .A2(G288), .ZN(n935) );
  NAND2_X1 U764 ( .A1(G40), .A2(G160), .ZN(n682) );
  XNOR2_X1 U765 ( .A(n684), .B(KEYINPUT64), .ZN(n780) );
  NAND2_X1 U766 ( .A1(n781), .A2(n780), .ZN(n687) );
  INV_X1 U767 ( .A(n687), .ZN(n685) );
  NAND2_X1 U768 ( .A1(n685), .A2(G1996), .ZN(n686) );
  XNOR2_X1 U769 ( .A(n686), .B(KEYINPUT26), .ZN(n689) );
  BUF_X2 U770 ( .A(n687), .Z(n732) );
  NAND2_X1 U771 ( .A1(G1341), .A2(n732), .ZN(n688) );
  NAND2_X1 U772 ( .A1(n689), .A2(n688), .ZN(n691) );
  XNOR2_X1 U773 ( .A(n691), .B(n690), .ZN(n692) );
  OR2_X1 U774 ( .A1(n926), .A2(n693), .ZN(n701) );
  NAND2_X1 U775 ( .A1(n693), .A2(n926), .ZN(n699) );
  NAND2_X1 U776 ( .A1(n732), .A2(G1348), .ZN(n694) );
  XNOR2_X1 U777 ( .A(n694), .B(KEYINPUT98), .ZN(n697) );
  INV_X1 U778 ( .A(n732), .ZN(n695) );
  NAND2_X1 U779 ( .A1(n695), .A2(G2067), .ZN(n696) );
  NAND2_X1 U780 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U781 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U782 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U783 ( .A(n702), .B(KEYINPUT99), .ZN(n707) );
  NAND2_X1 U784 ( .A1(n695), .A2(G2072), .ZN(n703) );
  XOR2_X1 U785 ( .A(KEYINPUT27), .B(n703), .Z(n705) );
  NAND2_X1 U786 ( .A1(G1956), .A2(n732), .ZN(n704) );
  NAND2_X1 U787 ( .A1(n705), .A2(n704), .ZN(n710) );
  NOR2_X1 U788 ( .A1(G299), .A2(n710), .ZN(n706) );
  NOR2_X2 U789 ( .A1(n707), .A2(n706), .ZN(n709) );
  XNOR2_X1 U790 ( .A(n709), .B(n708), .ZN(n714) );
  NAND2_X1 U791 ( .A1(n710), .A2(G299), .ZN(n712) );
  XNOR2_X1 U792 ( .A(KEYINPUT28), .B(KEYINPUT96), .ZN(n711) );
  XNOR2_X1 U793 ( .A(n712), .B(n711), .ZN(n713) );
  NAND2_X1 U794 ( .A1(n714), .A2(n713), .ZN(n716) );
  XNOR2_X1 U795 ( .A(KEYINPUT29), .B(KEYINPUT101), .ZN(n715) );
  XNOR2_X1 U796 ( .A(n716), .B(n715), .ZN(n720) );
  INV_X1 U797 ( .A(G1961), .ZN(n932) );
  NAND2_X1 U798 ( .A1(n732), .A2(n932), .ZN(n718) );
  XNOR2_X1 U799 ( .A(G2078), .B(KEYINPUT25), .ZN(n958) );
  NAND2_X1 U800 ( .A1(n695), .A2(n958), .ZN(n717) );
  NAND2_X1 U801 ( .A1(n718), .A2(n717), .ZN(n726) );
  NAND2_X1 U802 ( .A1(n726), .A2(G171), .ZN(n719) );
  NAND2_X1 U803 ( .A1(n720), .A2(n719), .ZN(n731) );
  NAND2_X1 U804 ( .A1(G8), .A2(n732), .ZN(n773) );
  NOR2_X1 U805 ( .A1(G1966), .A2(n773), .ZN(n744) );
  NOR2_X1 U806 ( .A1(G2084), .A2(n732), .ZN(n721) );
  XOR2_X1 U807 ( .A(KEYINPUT95), .B(n721), .Z(n741) );
  INV_X1 U808 ( .A(n741), .ZN(n722) );
  NAND2_X1 U809 ( .A1(G8), .A2(n722), .ZN(n723) );
  NOR2_X1 U810 ( .A1(n744), .A2(n723), .ZN(n724) );
  XOR2_X1 U811 ( .A(KEYINPUT30), .B(n724), .Z(n725) );
  NOR2_X1 U812 ( .A1(G168), .A2(n725), .ZN(n728) );
  NOR2_X1 U813 ( .A1(G171), .A2(n726), .ZN(n727) );
  NOR2_X1 U814 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U815 ( .A(KEYINPUT31), .B(n729), .Z(n730) );
  NAND2_X1 U816 ( .A1(n731), .A2(n730), .ZN(n742) );
  NAND2_X1 U817 ( .A1(n742), .A2(G286), .ZN(n739) );
  INV_X1 U818 ( .A(G8), .ZN(n737) );
  NOR2_X1 U819 ( .A1(G2090), .A2(n732), .ZN(n734) );
  NOR2_X1 U820 ( .A1(G1971), .A2(n773), .ZN(n733) );
  NOR2_X1 U821 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U822 ( .A1(n735), .A2(G303), .ZN(n736) );
  OR2_X1 U823 ( .A1(n737), .A2(n736), .ZN(n738) );
  AND2_X1 U824 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U825 ( .A(n740), .B(KEYINPUT32), .ZN(n748) );
  NAND2_X1 U826 ( .A1(G8), .A2(n741), .ZN(n746) );
  INV_X1 U827 ( .A(n742), .ZN(n743) );
  NOR2_X1 U828 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U829 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U830 ( .A1(n748), .A2(n747), .ZN(n767) );
  NOR2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n756) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n749) );
  NOR2_X1 U833 ( .A1(n756), .A2(n749), .ZN(n936) );
  NAND2_X1 U834 ( .A1(n767), .A2(n936), .ZN(n750) );
  NAND2_X1 U835 ( .A1(n935), .A2(n750), .ZN(n752) );
  INV_X1 U836 ( .A(KEYINPUT102), .ZN(n755) );
  OR2_X1 U837 ( .A1(n773), .A2(n755), .ZN(n751) );
  NOR2_X1 U838 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U839 ( .A1(KEYINPUT33), .A2(n753), .ZN(n754) );
  INV_X1 U840 ( .A(n754), .ZN(n764) );
  NAND2_X1 U841 ( .A1(n755), .A2(n756), .ZN(n759) );
  NAND2_X1 U842 ( .A1(n756), .A2(KEYINPUT33), .ZN(n757) );
  NAND2_X1 U843 ( .A1(n757), .A2(KEYINPUT102), .ZN(n758) );
  NAND2_X1 U844 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U845 ( .A1(n773), .A2(n760), .ZN(n762) );
  XOR2_X1 U846 ( .A(G1981), .B(G305), .Z(n945) );
  NOR2_X1 U847 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U848 ( .A1(n764), .A2(n763), .ZN(n777) );
  NOR2_X1 U849 ( .A1(G2090), .A2(G303), .ZN(n765) );
  NAND2_X1 U850 ( .A1(G8), .A2(n765), .ZN(n766) );
  NAND2_X1 U851 ( .A1(n767), .A2(n766), .ZN(n769) );
  XNOR2_X1 U852 ( .A(n769), .B(n768), .ZN(n770) );
  NAND2_X1 U853 ( .A1(n770), .A2(n773), .ZN(n775) );
  NOR2_X1 U854 ( .A1(G1981), .A2(G305), .ZN(n771) );
  XOR2_X1 U855 ( .A(n771), .B(KEYINPUT24), .Z(n772) );
  OR2_X1 U856 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U857 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U858 ( .A1(n777), .A2(n776), .ZN(n779) );
  XNOR2_X1 U859 ( .A(n779), .B(n778), .ZN(n818) );
  XNOR2_X1 U860 ( .A(G1986), .B(G290), .ZN(n943) );
  INV_X1 U861 ( .A(n780), .ZN(n782) );
  NAND2_X1 U862 ( .A1(n782), .A2(n781), .ZN(n812) );
  INV_X1 U863 ( .A(n812), .ZN(n829) );
  NAND2_X1 U864 ( .A1(n943), .A2(n829), .ZN(n816) );
  XNOR2_X1 U865 ( .A(G2067), .B(KEYINPUT37), .ZN(n827) );
  NAND2_X1 U866 ( .A1(n899), .A2(G104), .ZN(n784) );
  NAND2_X1 U867 ( .A1(G140), .A2(n604), .ZN(n783) );
  NAND2_X1 U868 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U869 ( .A(KEYINPUT34), .B(n785), .ZN(n791) );
  NAND2_X1 U870 ( .A1(G128), .A2(n521), .ZN(n787) );
  NAND2_X1 U871 ( .A1(G116), .A2(n904), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U873 ( .A(KEYINPUT88), .B(n788), .Z(n789) );
  XNOR2_X1 U874 ( .A(KEYINPUT35), .B(n789), .ZN(n790) );
  NOR2_X1 U875 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U876 ( .A(KEYINPUT36), .B(n792), .ZN(n912) );
  OR2_X1 U877 ( .A1(n827), .A2(n912), .ZN(n793) );
  XNOR2_X1 U878 ( .A(n793), .B(KEYINPUT89), .ZN(n1000) );
  NAND2_X1 U879 ( .A1(n829), .A2(n1000), .ZN(n825) );
  INV_X1 U880 ( .A(n825), .ZN(n814) );
  XOR2_X1 U881 ( .A(KEYINPUT90), .B(G1991), .Z(n953) );
  NAND2_X1 U882 ( .A1(n899), .A2(G95), .ZN(n795) );
  NAND2_X1 U883 ( .A1(G131), .A2(n604), .ZN(n794) );
  NAND2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n799) );
  NAND2_X1 U885 ( .A1(G119), .A2(n521), .ZN(n797) );
  NAND2_X1 U886 ( .A1(G107), .A2(n904), .ZN(n796) );
  NAND2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U888 ( .A1(n799), .A2(n798), .ZN(n882) );
  NOR2_X1 U889 ( .A1(n953), .A2(n882), .ZN(n810) );
  NAND2_X1 U890 ( .A1(G129), .A2(n521), .ZN(n801) );
  NAND2_X1 U891 ( .A1(G117), .A2(n904), .ZN(n800) );
  NAND2_X1 U892 ( .A1(n801), .A2(n800), .ZN(n804) );
  NAND2_X1 U893 ( .A1(n899), .A2(G105), .ZN(n802) );
  XOR2_X1 U894 ( .A(KEYINPUT38), .B(n802), .Z(n803) );
  NOR2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U896 ( .A(KEYINPUT91), .B(n805), .Z(n807) );
  NAND2_X1 U897 ( .A1(G141), .A2(n604), .ZN(n806) );
  NAND2_X1 U898 ( .A1(n807), .A2(n806), .ZN(n896) );
  NAND2_X1 U899 ( .A1(G1996), .A2(n896), .ZN(n808) );
  XOR2_X1 U900 ( .A(KEYINPUT92), .B(n808), .Z(n809) );
  NOR2_X1 U901 ( .A1(n810), .A2(n809), .ZN(n811) );
  XOR2_X1 U902 ( .A(KEYINPUT93), .B(n811), .Z(n998) );
  NOR2_X1 U903 ( .A1(n998), .A2(n812), .ZN(n813) );
  XNOR2_X1 U904 ( .A(KEYINPUT94), .B(n813), .ZN(n821) );
  NOR2_X1 U905 ( .A1(n814), .A2(n821), .ZN(n815) );
  AND2_X1 U906 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U907 ( .A1(n818), .A2(n817), .ZN(n832) );
  NOR2_X1 U908 ( .A1(G1996), .A2(n896), .ZN(n981) );
  AND2_X1 U909 ( .A1(n953), .A2(n882), .ZN(n979) );
  NOR2_X1 U910 ( .A1(G1986), .A2(G290), .ZN(n819) );
  NOR2_X1 U911 ( .A1(n979), .A2(n819), .ZN(n820) );
  NOR2_X1 U912 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U913 ( .A1(n981), .A2(n822), .ZN(n824) );
  XOR2_X1 U914 ( .A(KEYINPUT39), .B(KEYINPUT105), .Z(n823) );
  XNOR2_X1 U915 ( .A(n824), .B(n823), .ZN(n826) );
  NAND2_X1 U916 ( .A1(n826), .A2(n825), .ZN(n828) );
  NAND2_X1 U917 ( .A1(n912), .A2(n827), .ZN(n989) );
  NAND2_X1 U918 ( .A1(n828), .A2(n989), .ZN(n830) );
  NAND2_X1 U919 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U920 ( .A1(n832), .A2(n831), .ZN(n834) );
  XNOR2_X1 U921 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n833) );
  XNOR2_X1 U922 ( .A(n834), .B(n833), .ZN(G329) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n835), .ZN(G217) );
  INV_X1 U924 ( .A(n835), .ZN(G223) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U926 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U928 ( .A1(n838), .A2(n837), .ZN(G188) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  INV_X1 U932 ( .A(G69), .ZN(G235) );
  NOR2_X1 U933 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U935 ( .A(G2443), .B(G2438), .ZN(n850) );
  XOR2_X1 U936 ( .A(G2454), .B(G2430), .Z(n842) );
  XNOR2_X1 U937 ( .A(G2446), .B(KEYINPUT107), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U939 ( .A(G2451), .B(G2427), .Z(n844) );
  XNOR2_X1 U940 ( .A(G1341), .B(G1348), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U942 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U943 ( .A(G2435), .B(KEYINPUT108), .ZN(n847) );
  XNOR2_X1 U944 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U945 ( .A(n850), .B(n849), .ZN(n851) );
  NAND2_X1 U946 ( .A1(n851), .A2(G14), .ZN(n852) );
  XNOR2_X1 U947 ( .A(KEYINPUT109), .B(n852), .ZN(G401) );
  XOR2_X1 U948 ( .A(G2096), .B(G2090), .Z(n854) );
  XNOR2_X1 U949 ( .A(G2067), .B(G2072), .ZN(n853) );
  XNOR2_X1 U950 ( .A(n854), .B(n853), .ZN(n865) );
  XOR2_X1 U951 ( .A(KEYINPUT42), .B(KEYINPUT113), .Z(n856) );
  XNOR2_X1 U952 ( .A(G2678), .B(KEYINPUT110), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(n861) );
  XNOR2_X1 U954 ( .A(n857), .B(KEYINPUT43), .ZN(n859) );
  XNOR2_X1 U955 ( .A(KEYINPUT112), .B(KEYINPUT111), .ZN(n858) );
  XNOR2_X1 U956 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U957 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U958 ( .A(G2078), .B(G2084), .ZN(n862) );
  XNOR2_X1 U959 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U960 ( .A(n865), .B(n864), .Z(G227) );
  XNOR2_X1 U961 ( .A(G1981), .B(n932), .ZN(n867) );
  XNOR2_X1 U962 ( .A(G1966), .B(G1956), .ZN(n866) );
  XNOR2_X1 U963 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U964 ( .A(n868), .B(G2474), .Z(n870) );
  XNOR2_X1 U965 ( .A(G1996), .B(G1991), .ZN(n869) );
  XNOR2_X1 U966 ( .A(n870), .B(n869), .ZN(n874) );
  XOR2_X1 U967 ( .A(KEYINPUT41), .B(G1976), .Z(n872) );
  XNOR2_X1 U968 ( .A(G1986), .B(G1971), .ZN(n871) );
  XNOR2_X1 U969 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U970 ( .A(n874), .B(n873), .ZN(G229) );
  NAND2_X1 U971 ( .A1(n521), .A2(G124), .ZN(n875) );
  XNOR2_X1 U972 ( .A(n875), .B(KEYINPUT44), .ZN(n877) );
  NAND2_X1 U973 ( .A1(G112), .A2(n904), .ZN(n876) );
  NAND2_X1 U974 ( .A1(n877), .A2(n876), .ZN(n881) );
  NAND2_X1 U975 ( .A1(n899), .A2(G100), .ZN(n879) );
  NAND2_X1 U976 ( .A1(G136), .A2(n604), .ZN(n878) );
  NAND2_X1 U977 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U978 ( .A1(n881), .A2(n880), .ZN(G162) );
  XOR2_X1 U979 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n884) );
  XNOR2_X1 U980 ( .A(G164), .B(n882), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n884), .B(n883), .ZN(n894) );
  NAND2_X1 U982 ( .A1(G130), .A2(n521), .ZN(n886) );
  NAND2_X1 U983 ( .A1(G118), .A2(n904), .ZN(n885) );
  NAND2_X1 U984 ( .A1(n886), .A2(n885), .ZN(n892) );
  NAND2_X1 U985 ( .A1(n899), .A2(G106), .ZN(n887) );
  XNOR2_X1 U986 ( .A(n887), .B(KEYINPUT114), .ZN(n889) );
  NAND2_X1 U987 ( .A1(G142), .A2(n604), .ZN(n888) );
  NAND2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U989 ( .A(n890), .B(KEYINPUT45), .Z(n891) );
  NOR2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U991 ( .A(n894), .B(n893), .Z(n898) );
  XOR2_X1 U992 ( .A(G160), .B(G162), .Z(n895) );
  XNOR2_X1 U993 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U994 ( .A(n898), .B(n897), .Z(n911) );
  NAND2_X1 U995 ( .A1(n899), .A2(G103), .ZN(n901) );
  NAND2_X1 U996 ( .A1(G139), .A2(n604), .ZN(n900) );
  NAND2_X1 U997 ( .A1(n901), .A2(n900), .ZN(n909) );
  NAND2_X1 U998 ( .A1(n521), .A2(G127), .ZN(n903) );
  XOR2_X1 U999 ( .A(KEYINPUT115), .B(n903), .Z(n906) );
  NAND2_X1 U1000 ( .A1(n904), .A2(G115), .ZN(n905) );
  NAND2_X1 U1001 ( .A1(n906), .A2(n905), .ZN(n907) );
  XOR2_X1 U1002 ( .A(KEYINPUT47), .B(n907), .Z(n908) );
  NOR2_X1 U1003 ( .A1(n909), .A2(n908), .ZN(n991) );
  XNOR2_X1 U1004 ( .A(n991), .B(n988), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(n911), .B(n910), .ZN(n913) );
  XOR2_X1 U1006 ( .A(n913), .B(n912), .Z(n914) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n914), .ZN(G395) );
  XOR2_X1 U1008 ( .A(G301), .B(G286), .Z(n916) );
  XNOR2_X1 U1009 ( .A(n916), .B(n915), .ZN(n918) );
  XNOR2_X1 U1010 ( .A(n927), .B(n926), .ZN(n917) );
  XNOR2_X1 U1011 ( .A(n918), .B(n917), .ZN(n919) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n919), .ZN(G397) );
  OR2_X1 U1013 ( .A1(n925), .A2(G401), .ZN(n922) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n920) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n920), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(n922), .A2(n921), .ZN(n924) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1018 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G303), .ZN(G166) );
  INV_X1 U1021 ( .A(n925), .ZN(G319) );
  INV_X1 U1022 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1023 ( .A(G16), .B(KEYINPUT56), .Z(n952) );
  XNOR2_X1 U1024 ( .A(n926), .B(G1348), .ZN(n931) );
  XNOR2_X1 U1025 ( .A(G299), .B(G1956), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(n927), .B(G1341), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n934) );
  XOR2_X1 U1029 ( .A(n932), .B(G301), .Z(n933) );
  NOR2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n941) );
  NAND2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n938) );
  AND2_X1 U1032 ( .A1(G303), .A2(G1971), .ZN(n937) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1034 ( .A(KEYINPUT121), .B(n939), .Z(n940) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1036 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(KEYINPUT122), .B(n944), .ZN(n949) );
  XNOR2_X1 U1038 ( .A(G1966), .B(G168), .ZN(n946) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(KEYINPUT57), .B(n947), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(n950), .B(KEYINPUT123), .ZN(n951) );
  NOR2_X1 U1043 ( .A1(n952), .A2(n951), .ZN(n977) );
  XOR2_X1 U1044 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n1002) );
  XNOR2_X1 U1045 ( .A(G2090), .B(G35), .ZN(n968) );
  XNOR2_X1 U1046 ( .A(n953), .B(G25), .ZN(n956) );
  XOR2_X1 U1047 ( .A(G2072), .B(KEYINPUT120), .Z(n954) );
  XNOR2_X1 U1048 ( .A(G33), .B(n954), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n965) );
  XNOR2_X1 U1050 ( .A(KEYINPUT119), .B(G2067), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(n957), .B(G26), .ZN(n963) );
  XNOR2_X1 U1052 ( .A(G27), .B(n958), .ZN(n959) );
  NAND2_X1 U1053 ( .A1(n959), .A2(G28), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(G32), .B(G1996), .ZN(n960) );
  NOR2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(KEYINPUT53), .B(n966), .ZN(n967) );
  NOR2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n971) );
  XOR2_X1 U1060 ( .A(G2084), .B(G34), .Z(n969) );
  XNOR2_X1 U1061 ( .A(KEYINPUT54), .B(n969), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1063 ( .A(n1002), .B(n972), .ZN(n974) );
  INV_X1 U1064 ( .A(G29), .ZN(n973) );
  NAND2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1066 ( .A1(G11), .A2(n975), .ZN(n976) );
  NOR2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n1006) );
  XOR2_X1 U1068 ( .A(G160), .B(G2084), .Z(n978) );
  NOR2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n986) );
  XOR2_X1 U1070 ( .A(G2090), .B(G162), .Z(n980) );
  NOR2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1072 ( .A(KEYINPUT117), .B(n982), .Z(n984) );
  XOR2_X1 U1073 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n983) );
  XNOR2_X1 U1074 ( .A(n984), .B(n983), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n990) );
  NAND2_X1 U1077 ( .A1(n990), .A2(n989), .ZN(n996) );
  XOR2_X1 U1078 ( .A(G2072), .B(n991), .Z(n993) );
  XOR2_X1 U1079 ( .A(G164), .B(G2078), .Z(n992) );
  NOR2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1081 ( .A(KEYINPUT50), .B(n994), .Z(n995) );
  NOR2_X1 U1082 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1083 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1084 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1085 ( .A(KEYINPUT52), .B(n1001), .ZN(n1003) );
  NAND2_X1 U1086 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1087 ( .A1(n1004), .A2(G29), .ZN(n1005) );
  NAND2_X1 U1088 ( .A1(n1006), .A2(n1005), .ZN(n1032) );
  XOR2_X1 U1089 ( .A(G1976), .B(G23), .Z(n1008) );
  XOR2_X1 U1090 ( .A(G1971), .B(G22), .Z(n1007) );
  NAND2_X1 U1091 ( .A1(n1008), .A2(n1007), .ZN(n1010) );
  XNOR2_X1 U1092 ( .A(G24), .B(G1986), .ZN(n1009) );
  NOR2_X1 U1093 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1094 ( .A(KEYINPUT58), .B(n1011), .Z(n1028) );
  XOR2_X1 U1095 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n1021) );
  XNOR2_X1 U1096 ( .A(G1341), .B(G19), .ZN(n1013) );
  XNOR2_X1 U1097 ( .A(G6), .B(G1981), .ZN(n1012) );
  NOR2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1019) );
  XOR2_X1 U1099 ( .A(G4), .B(KEYINPUT124), .Z(n1015) );
  XNOR2_X1 U1100 ( .A(G1348), .B(KEYINPUT59), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(n1015), .B(n1014), .ZN(n1017) );
  XNOR2_X1 U1102 ( .A(G1956), .B(G20), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(n1021), .B(n1020), .ZN(n1025) );
  XOR2_X1 U1106 ( .A(G1966), .B(G21), .Z(n1023) );
  XOR2_X1 U1107 ( .A(G1961), .B(G5), .Z(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1110 ( .A(KEYINPUT126), .B(n1026), .Z(n1027) );
  NOR2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1112 ( .A(KEYINPUT61), .B(n1029), .Z(n1030) );
  NOR2_X1 U1113 ( .A1(G16), .A2(n1030), .ZN(n1031) );
  NOR2_X1 U1114 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1115 ( .A(n1033), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1116 ( .A(G150), .ZN(G311) );
endmodule

