//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n618,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1155, new_n1156;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n459), .A2(KEYINPUT68), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(KEYINPUT68), .ZN(new_n461));
  INV_X1    g036(.A(new_n454), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G567), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n460), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n466), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n467), .A2(new_n468), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(KEYINPUT69), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n470), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n480), .A2(new_n481), .A3(G125), .ZN(new_n482));
  NAND2_X1  g057(.A1(G113), .A2(G2104), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n476), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n473), .B1(new_n484), .B2(G2105), .ZN(G160));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G112), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n474), .A2(new_n466), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G124), .ZN(new_n490));
  AOI21_X1  g065(.A(G2105), .B1(new_n478), .B2(new_n479), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G136), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n492), .A2(KEYINPUT70), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n492), .A2(KEYINPUT70), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  INV_X1    g071(.A(KEYINPUT72), .ZN(new_n497));
  OR2_X1    g072(.A1(new_n466), .A2(G114), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(G126), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n502), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n501), .B1(new_n507), .B2(new_n474), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n506), .B1(new_n491), .B2(G138), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n497), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(G126), .A2(G2105), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n466), .A2(G138), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(new_n505), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(new_n480), .B1(new_n498), .B2(new_n500), .ZN(new_n514));
  OAI211_X1 g089(.A(G138), .B(new_n466), .C1(new_n467), .C2(new_n468), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(new_n505), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n514), .A2(KEYINPUT72), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n510), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(G164));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(G50), .A3(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT73), .A2(KEYINPUT5), .ZN(new_n522));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(new_n520), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n521), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n526), .A2(G62), .ZN(new_n531));
  NAND2_X1  g106(.A1(G75), .A2(G543), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n529), .A2(new_n533), .ZN(G166));
  INV_X1    g109(.A(new_n527), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n535), .A2(G89), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n520), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G51), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n537), .B(new_n539), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n536), .A2(new_n542), .ZN(G168));
  AOI22_X1  g118(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n530), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT74), .B(G90), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n527), .A2(new_n546), .B1(new_n540), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(G171));
  INV_X1    g124(.A(new_n540), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n535), .A2(G81), .B1(new_n550), .B2(G43), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n530), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT75), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OR3_X1    g136(.A1(new_n540), .A2(KEYINPUT9), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT9), .B1(new_n540), .B2(new_n561), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(new_n526), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n562), .A2(new_n563), .B1(G651), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(G91), .ZN(new_n569));
  OR3_X1    g144(.A1(new_n527), .A2(KEYINPUT76), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT76), .B1(new_n527), .B2(new_n569), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  INV_X1    g150(.A(new_n533), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n535), .A2(G88), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n576), .A2(new_n577), .A3(new_n521), .A4(KEYINPUT77), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n579), .B1(new_n529), .B2(new_n533), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n578), .A2(new_n580), .ZN(G303));
  AOI22_X1  g156(.A1(new_n535), .A2(G87), .B1(new_n550), .B2(G49), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(new_n535), .A2(G86), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n550), .A2(G48), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n526), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n530), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n530), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n527), .A2(new_n594), .B1(new_n540), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NOR2_X1   g174(.A1(G171), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT78), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OR3_X1    g177(.A1(new_n527), .A2(KEYINPUT79), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(KEYINPUT79), .B1(new_n527), .B2(new_n602), .ZN(new_n604));
  AOI21_X1  g179(.A(KEYINPUT10), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n526), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G54), .ZN(new_n607));
  OAI22_X1  g182(.A1(new_n606), .A2(new_n530), .B1(new_n607), .B2(new_n540), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n603), .A2(KEYINPUT10), .A3(new_n604), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT80), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n601), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n601), .B1(new_n612), .B2(G868), .ZN(G321));
  NAND2_X1  g189(.A1(G299), .A2(new_n599), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n599), .B2(G168), .ZN(G297));
  OAI21_X1  g191(.A(new_n615), .B1(new_n599), .B2(G168), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n612), .B1(new_n618), .B2(G860), .ZN(G148));
  NOR2_X1   g194(.A1(new_n555), .A2(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n612), .A2(new_n618), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT81), .Z(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n480), .A2(new_n471), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n489), .A2(G123), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n466), .A2(G111), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  AND3_X1   g206(.A1(new_n491), .A2(KEYINPUT82), .A3(G135), .ZN(new_n632));
  AOI21_X1  g207(.A(KEYINPUT82), .B1(new_n491), .B2(G135), .ZN(new_n633));
  OAI221_X1 g208(.A(new_n629), .B1(new_n630), .B2(new_n631), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  AOI22_X1  g209(.A1(new_n628), .A2(G2100), .B1(G2096), .B2(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(G2096), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n635), .B(new_n636), .C1(G2100), .C2(new_n628), .ZN(G156));
  INV_X1    g212(.A(KEYINPUT14), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n641), .B2(new_n640), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n643), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  AND3_X1   g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  NAND3_X1  g231(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT18), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT83), .B(KEYINPUT17), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n653), .B(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n656), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n660), .A2(new_n655), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n661), .B1(new_n654), .B2(new_n655), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n660), .B2(new_n655), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n658), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2096), .B(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT85), .Z(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n670), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT20), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n675), .A2(new_n671), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT84), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n676), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1991), .B(G1996), .Z(new_n684));
  XOR2_X1   g259(.A(new_n683), .B(new_n684), .Z(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G229));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n688), .A2(G33), .ZN(new_n689));
  AOI22_X1  g264(.A1(new_n480), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n690), .A2(new_n466), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT93), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n491), .A2(G139), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT92), .Z(new_n694));
  XOR2_X1   g269(.A(KEYINPUT91), .B(KEYINPUT25), .Z(new_n695));
  NAND3_X1  g270(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n692), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT94), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n689), .B1(new_n699), .B2(G29), .ZN(new_n700));
  INV_X1    g275(.A(G2072), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n489), .A2(G129), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n471), .A2(G105), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G141), .B2(new_n491), .ZN(new_n707));
  NAND3_X1  g282(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT96), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT26), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n712), .A2(new_n688), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n688), .B2(G32), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT27), .B(G1996), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT24), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G34), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n688), .B1(new_n716), .B2(G34), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT95), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n719), .B2(new_n718), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G160), .B2(G29), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n714), .A2(new_n715), .B1(G2084), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n702), .A2(new_n703), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT97), .ZN(new_n725));
  NOR2_X1   g300(.A1(G4), .A2(G16), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n612), .B2(G16), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT89), .B(G1348), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G20), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT23), .Z(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G299), .B2(G16), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1956), .ZN(new_n734));
  NOR2_X1   g309(.A1(G29), .A2(G35), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G162), .B2(G29), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G2090), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n734), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT100), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n738), .A2(new_n739), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n489), .A2(G128), .B1(G140), .B2(new_n491), .ZN(new_n743));
  NOR2_X1   g318(.A1(G104), .A2(G2105), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT90), .ZN(new_n745));
  OAI21_X1  g320(.A(G2104), .B1(new_n466), .B2(G116), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n743), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G29), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n688), .A2(G26), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT28), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G2067), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n714), .B2(new_n715), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n730), .A2(G21), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G168), .B2(new_n730), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n756), .A2(G1966), .ZN(new_n757));
  NOR2_X1   g332(.A1(G5), .A2(G16), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT98), .Z(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G171), .B2(G16), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G1961), .ZN(new_n761));
  INV_X1    g336(.A(new_n756), .ZN(new_n762));
  INV_X1    g337(.A(G1966), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT30), .B(G28), .ZN(new_n765));
  OR2_X1    g340(.A1(KEYINPUT31), .A2(G11), .ZN(new_n766));
  NAND2_X1  g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n765), .A2(new_n688), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI221_X1 g343(.A(new_n768), .B1(new_n688), .B2(new_n634), .C1(new_n760), .C2(G1961), .ZN(new_n769));
  NOR4_X1   g344(.A1(new_n754), .A2(new_n757), .A3(new_n764), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n730), .A2(G19), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n555), .B2(new_n730), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(G1341), .Z(new_n773));
  NAND2_X1  g348(.A1(G164), .A2(G29), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G27), .B2(G29), .ZN(new_n775));
  INV_X1    g350(.A(G2078), .ZN(new_n776));
  OAI22_X1  g351(.A1(new_n775), .A2(new_n776), .B1(G2084), .B2(new_n722), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n776), .B2(new_n775), .ZN(new_n778));
  AND4_X1   g353(.A1(new_n742), .A2(new_n770), .A3(new_n773), .A4(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n725), .A2(new_n729), .A3(new_n741), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT101), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n730), .A2(G23), .ZN(new_n782));
  INV_X1    g357(.A(G288), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n730), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT33), .B(G1976), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT87), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n784), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n730), .A2(G22), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G166), .B2(new_n730), .ZN(new_n789));
  INV_X1    g364(.A(G1971), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G6), .A2(G16), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n590), .B2(G16), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT32), .B(G1981), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n787), .A2(new_n791), .A3(new_n795), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n796), .A2(KEYINPUT34), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(KEYINPUT34), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n688), .A2(G25), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n489), .A2(G119), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n491), .A2(G131), .ZN(new_n801));
  OR2_X1    g376(.A1(G95), .A2(G2105), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n802), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n799), .B1(new_n805), .B2(new_n688), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT35), .B(G1991), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n730), .A2(G24), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT86), .Z(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G290), .B2(G16), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1986), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n797), .A2(new_n798), .A3(new_n808), .A4(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT88), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT36), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n813), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n781), .A2(new_n817), .ZN(G311));
  NAND2_X1  g393(.A1(new_n781), .A2(new_n817), .ZN(G150));
  AOI22_X1  g394(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n820), .A2(new_n530), .ZN(new_n821));
  INV_X1    g396(.A(G93), .ZN(new_n822));
  INV_X1    g397(.A(G55), .ZN(new_n823));
  OAI22_X1  g398(.A1(new_n527), .A2(new_n822), .B1(new_n540), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n555), .A2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n825), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n828), .A2(new_n553), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT38), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n612), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n835));
  AOI21_X1  g410(.A(G860), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n835), .B2(new_n834), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n828), .A2(G860), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(G145));
  INV_X1    g415(.A(new_n699), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n508), .A2(new_n509), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n747), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n711), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n698), .ZN(new_n846));
  OAI22_X1  g421(.A1(new_n845), .A2(KEYINPUT103), .B1(new_n846), .B2(new_n844), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n845), .A2(KEYINPUT103), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n489), .A2(G130), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n466), .A2(G118), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(G142), .B2(new_n491), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n626), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n805), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n849), .A2(new_n856), .ZN(new_n857));
  OR3_X1    g432(.A1(new_n847), .A2(new_n848), .A3(new_n856), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n857), .A2(KEYINPUT104), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(G160), .B(KEYINPUT102), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n495), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n634), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT104), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n849), .A2(new_n864), .A3(new_n856), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n859), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n863), .B1(new_n849), .B2(new_n856), .ZN(new_n867));
  AOI21_X1  g442(.A(G37), .B1(new_n867), .B2(new_n858), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g445(.A(new_n621), .B(new_n831), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n611), .B(G299), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT41), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n872), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT42), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n590), .B(G290), .ZN(new_n878));
  XNOR2_X1  g453(.A(G288), .B(G166), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT42), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n874), .A2(new_n882), .A3(new_n875), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n877), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n881), .B1(new_n877), .B2(new_n883), .ZN(new_n885));
  OAI21_X1  g460(.A(G868), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(G868), .B2(new_n825), .ZN(G295));
  OAI21_X1  g462(.A(new_n886), .B1(G868), .B2(new_n825), .ZN(G331));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n889));
  XNOR2_X1  g464(.A(G301), .B(G168), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n831), .A2(KEYINPUT105), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n872), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n827), .A2(new_n890), .A3(new_n830), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n891), .B1(new_n826), .B2(new_n829), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n892), .A2(new_n893), .A3(new_n894), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n894), .A2(new_n895), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n873), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(new_n900), .A3(new_n880), .ZN(new_n901));
  INV_X1    g476(.A(G37), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n898), .A2(new_n900), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n881), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n889), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n892), .A2(new_n894), .A3(new_n897), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n873), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n894), .A2(new_n893), .A3(new_n895), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n880), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n903), .A2(new_n911), .A3(KEYINPUT43), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT43), .B1(new_n904), .B2(new_n906), .ZN(new_n916));
  OR3_X1    g491(.A1(new_n903), .A2(new_n911), .A3(KEYINPUT106), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT106), .B1(new_n903), .B2(new_n911), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n916), .B1(new_n919), .B2(KEYINPUT43), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n915), .B1(new_n920), .B2(new_n914), .ZN(G397));
  XNOR2_X1  g496(.A(KEYINPUT107), .B(G40), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(G160), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(new_n842), .B2(G1384), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G1996), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n929), .B(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT46), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n931), .B(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n747), .B(G2067), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n927), .B1(new_n934), .B2(new_n711), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(KEYINPUT47), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n931), .A2(new_n712), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n934), .A2(new_n927), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n927), .A2(G1996), .A3(new_n711), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n940), .B(KEYINPUT110), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n805), .A2(new_n807), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n747), .A2(G2067), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n927), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  XOR2_X1   g521(.A(new_n804), .B(new_n807), .Z(new_n947));
  AOI21_X1  g522(.A(new_n942), .B1(new_n927), .B2(new_n947), .ZN(new_n948));
  NOR4_X1   g523(.A1(new_n924), .A2(G290), .A3(new_n926), .A4(G1986), .ZN(new_n949));
  XOR2_X1   g524(.A(new_n949), .B(KEYINPUT48), .Z(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n937), .A2(new_n946), .A3(new_n951), .ZN(new_n952));
  XOR2_X1   g527(.A(new_n952), .B(KEYINPUT127), .Z(new_n953));
  AOI211_X1 g528(.A(new_n473), .B(new_n922), .C1(new_n484), .C2(G2105), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n925), .A2(G1384), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n956), .B1(new_n510), .B2(new_n517), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT114), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n954), .B(new_n926), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  AOI211_X1 g534(.A(KEYINPUT114), .B(new_n956), .C1(new_n510), .C2(new_n517), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n763), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT115), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(G1384), .B1(new_n514), .B2(new_n516), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(G1384), .B1(new_n510), .B2(new_n517), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n954), .B(new_n966), .C1(new_n967), .C2(new_n965), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n968), .A2(G2084), .ZN(new_n969));
  OAI211_X1 g544(.A(KEYINPUT115), .B(new_n763), .C1(new_n959), .C2(new_n960), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n963), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G8), .ZN(new_n972));
  NOR2_X1   g547(.A1(G168), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  XOR2_X1   g549(.A(KEYINPUT122), .B(KEYINPUT51), .Z(new_n975));
  OAI211_X1 g550(.A(G8), .B(new_n975), .C1(new_n971), .C2(G286), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n973), .A2(KEYINPUT51), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n971), .B2(G8), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT123), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n976), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AOI211_X1 g556(.A(KEYINPUT123), .B(new_n978), .C1(new_n971), .C2(G8), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n974), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT62), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT62), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n985), .B(new_n974), .C1(new_n981), .C2(new_n982), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n578), .A2(new_n580), .A3(KEYINPUT55), .A4(G8), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n988));
  OR2_X1    g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n578), .A2(G8), .A3(new_n580), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n989), .A2(new_n990), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n955), .B1(new_n508), .B2(new_n509), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n954), .B(new_n995), .C1(new_n967), .C2(KEYINPUT45), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n790), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(G2090), .B2(new_n968), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n994), .A2(new_n998), .A3(G8), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n954), .B1(new_n965), .B2(new_n964), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  AOI211_X1 g577(.A(KEYINPUT50), .B(G1384), .C1(new_n510), .C2(new_n517), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n739), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n997), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n994), .B1(G8), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n972), .B1(new_n954), .B2(new_n964), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n783), .A2(G1976), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(new_n783), .B2(G1976), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n589), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT113), .B(G1981), .Z(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1014), .A2(new_n585), .A3(new_n586), .A4(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1981), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1017), .B1(new_n590), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT49), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1017), .B(KEYINPUT49), .C1(new_n590), .C2(new_n1018), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n1008), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1024), .B1(new_n1010), .B2(KEYINPUT52), .ZN(new_n1025));
  AOI211_X1 g600(.A(KEYINPUT112), .B(new_n1011), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1013), .B(new_n1023), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1000), .A2(new_n1007), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n518), .A2(new_n955), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT114), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n964), .A2(KEYINPUT45), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n924), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n957), .A2(new_n958), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(G2078), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .A4(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G1961), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n968), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1035), .B1(new_n996), .B2(G2078), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT124), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(G160), .A2(new_n923), .A3(new_n995), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1044), .B(new_n776), .C1(KEYINPUT45), .C2(new_n967), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(KEYINPUT124), .A3(new_n1035), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1040), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n1029), .A2(G301), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n984), .A2(new_n986), .A3(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1045), .A2(KEYINPUT124), .A3(new_n1035), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT124), .B1(new_n1045), .B2(new_n1035), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1050), .B(G301), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(G160), .A2(G40), .A3(new_n995), .A4(new_n1036), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(new_n1032), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n1038), .B2(new_n968), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1057), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1053), .B(KEYINPUT54), .C1(new_n1058), .C2(G301), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1028), .A2(new_n1059), .ZN(new_n1060));
  OAI211_X1 g635(.A(G301), .B(new_n1056), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n1047), .B2(G301), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT125), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT125), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1062), .A2(new_n1066), .A3(new_n1063), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1060), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n1069));
  INV_X1    g644(.A(G1348), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n967), .A2(new_n965), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n954), .A2(new_n966), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(G160), .A2(new_n752), .A3(new_n923), .A4(new_n964), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1073), .A2(KEYINPUT60), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(new_n1070), .B2(new_n968), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1082), .A2(KEYINPUT120), .A3(KEYINPUT60), .A4(new_n1076), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1080), .A2(new_n612), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1073), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT60), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n1080), .B2(new_n612), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1069), .B1(new_n1084), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT119), .B1(new_n996), .B2(G1996), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n967), .A2(KEYINPUT45), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1091), .A2(new_n1092), .A3(new_n928), .A4(new_n1044), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n954), .A2(new_n964), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT58), .B(G1341), .Z(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1090), .A2(new_n1093), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n555), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT59), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1097), .A2(new_n1100), .A3(new_n555), .ZN(new_n1101));
  INV_X1    g676(.A(G1956), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n568), .A2(new_n572), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1104), .B1(new_n568), .B2(new_n572), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(G2072), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1044), .B(new_n1109), .C1(KEYINPUT45), .C2(new_n967), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1103), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1107), .B1(new_n1103), .B2(new_n1110), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT61), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1103), .A2(new_n1110), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1107), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT61), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1117), .A2(new_n1118), .A3(new_n1111), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1099), .A2(new_n1101), .B1(new_n1114), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1080), .A2(new_n612), .A3(new_n1083), .ZN(new_n1121));
  XOR2_X1   g696(.A(new_n611), .B(KEYINPUT80), .Z(new_n1122));
  NAND3_X1  g697(.A1(new_n1122), .A2(new_n1079), .A3(new_n1078), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1121), .A2(new_n1123), .A3(KEYINPUT121), .A4(new_n1087), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1089), .A2(new_n1120), .A3(new_n1124), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n612), .A2(new_n1085), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1111), .B1(new_n1126), .B2(new_n1113), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1068), .A2(new_n1128), .A3(new_n983), .ZN(new_n1129));
  NOR2_X1   g704(.A1(G288), .A2(G1976), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1023), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1017), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1008), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1133), .B1(new_n999), .B2(new_n1027), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT63), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n971), .A2(G8), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(G168), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1135), .B1(new_n1029), .B2(new_n1137), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1000), .A2(new_n1027), .A3(new_n1135), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n998), .A2(G8), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n994), .B1(new_n1140), .B2(KEYINPUT116), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(KEYINPUT116), .B2(new_n1140), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1139), .A2(new_n1142), .A3(G168), .A4(new_n1136), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1134), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1049), .A2(new_n1129), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n1146));
  AND2_X1   g721(.A1(G290), .A2(G1986), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n949), .B1(new_n927), .B2(new_n1147), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n1148), .B(KEYINPUT108), .Z(new_n1149));
  AND2_X1   g724(.A1(new_n948), .A2(new_n1149), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1145), .A2(new_n1146), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1146), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n953), .B1(new_n1151), .B2(new_n1152), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g728(.A1(G401), .A2(new_n464), .A3(G227), .ZN(new_n1155));
  AOI211_X1 g729(.A(G229), .B(new_n1155), .C1(new_n866), .C2(new_n868), .ZN(new_n1156));
  NAND2_X1  g730(.A1(new_n1156), .A2(new_n913), .ZN(G225));
  INV_X1    g731(.A(G225), .ZN(G308));
endmodule


