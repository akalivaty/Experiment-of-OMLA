

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729;

  XNOR2_X1 U361 ( .A(n590), .B(KEYINPUT32), .ZN(n725) );
  NAND2_X1 U362 ( .A1(n589), .A2(n343), .ZN(n342) );
  INV_X1 U363 ( .A(n592), .ZN(n343) );
  XNOR2_X1 U364 ( .A(n384), .B(n385), .ZN(n383) );
  XNOR2_X1 U365 ( .A(n462), .B(G113), .ZN(n386) );
  XNOR2_X2 U366 ( .A(n341), .B(n441), .ZN(n704) );
  NAND2_X1 U367 ( .A1(n435), .A2(n436), .ZN(n341) );
  OR2_X1 U368 ( .A1(n596), .A2(n342), .ZN(n590) );
  NAND2_X1 U369 ( .A1(n587), .A2(n583), .ZN(n647) );
  XNOR2_X2 U370 ( .A(G119), .B(G116), .ZN(n384) );
  NAND2_X2 U371 ( .A1(n644), .A2(n600), .ZN(n391) );
  XNOR2_X2 U372 ( .A(KEYINPUT68), .B(KEYINPUT85), .ZN(n385) );
  XNOR2_X2 U373 ( .A(KEYINPUT3), .B(KEYINPUT69), .ZN(n462) );
  XNOR2_X2 U374 ( .A(n576), .B(n575), .ZN(n582) );
  XNOR2_X2 U375 ( .A(n405), .B(n373), .ZN(n592) );
  BUF_X2 U376 ( .A(n654), .Z(n405) );
  XNOR2_X1 U377 ( .A(n474), .B(n452), .ZN(n488) );
  XNOR2_X1 U378 ( .A(n579), .B(KEYINPUT94), .ZN(n625) );
  XNOR2_X1 U379 ( .A(n467), .B(n488), .ZN(n507) );
  XNOR2_X1 U380 ( .A(n696), .B(n466), .ZN(n467) );
  NAND2_X1 U381 ( .A1(n347), .A2(n344), .ZN(n346) );
  NOR2_X1 U382 ( .A1(n679), .A2(n551), .ZN(n542) );
  INV_X1 U383 ( .A(n582), .ZN(n594) );
  NOR2_X1 U384 ( .A1(n574), .A2(n573), .ZN(n576) );
  NOR2_X1 U385 ( .A1(n567), .A2(n662), .ZN(n550) );
  INV_X1 U386 ( .A(KEYINPUT93), .ZN(n505) );
  NAND2_X1 U387 ( .A1(n380), .A2(n378), .ZN(n429) );
  AND2_X1 U388 ( .A1(n381), .A2(n618), .ZN(n380) );
  NAND2_X1 U389 ( .A1(n379), .A2(n607), .ZN(n378) );
  NOR2_X1 U390 ( .A1(n704), .A2(n392), .ZN(n390) );
  AND2_X1 U391 ( .A1(n433), .A2(n438), .ZN(n432) );
  XNOR2_X1 U392 ( .A(n345), .B(KEYINPUT105), .ZN(n436) );
  NAND2_X1 U393 ( .A1(n348), .A2(n346), .ZN(n345) );
  XNOR2_X1 U394 ( .A(n363), .B(KEYINPUT96), .ZN(n347) );
  OR2_X1 U395 ( .A1(n541), .A2(n540), .ZN(n551) );
  XNOR2_X1 U396 ( .A(n366), .B(KEYINPUT41), .ZN(n679) );
  AND2_X1 U397 ( .A1(n667), .A2(n664), .ZN(n366) );
  XNOR2_X1 U398 ( .A(n580), .B(KEYINPUT95), .ZN(n657) );
  AND2_X1 U399 ( .A1(n591), .A2(n405), .ZN(n580) );
  INV_X1 U400 ( .A(n666), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n374), .B(G472), .ZN(n654) );
  NOR2_X1 U402 ( .A1(n609), .A2(G902), .ZN(n489) );
  XNOR2_X1 U403 ( .A(n406), .B(n488), .ZN(n609) );
  XNOR2_X1 U404 ( .A(n356), .B(n398), .ZN(n406) );
  XNOR2_X1 U405 ( .A(n399), .B(n487), .ZN(n398) );
  XNOR2_X1 U406 ( .A(n512), .B(KEYINPUT16), .ZN(n463) );
  XNOR2_X1 U407 ( .A(n404), .B(G146), .ZN(n492) );
  XOR2_X1 U408 ( .A(G140), .B(G107), .Z(n487) );
  INV_X1 U409 ( .A(n729), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n654), .B(n450), .ZN(n597) );
  XNOR2_X2 U411 ( .A(n422), .B(n509), .ZN(n567) );
  NOR2_X1 U412 ( .A1(n727), .A2(n445), .ZN(n552) );
  NAND2_X1 U413 ( .A1(n597), .A2(n560), .ZN(n395) );
  OR2_X1 U414 ( .A1(n614), .A2(G902), .ZN(n374) );
  XNOR2_X1 U415 ( .A(n421), .B(n419), .ZN(n548) );
  XNOR2_X1 U416 ( .A(n534), .B(n420), .ZN(n419) );
  OR2_X1 U417 ( .A1(n606), .A2(G902), .ZN(n421) );
  NOR2_X1 U418 ( .A1(n726), .A2(n728), .ZN(n543) );
  NOR2_X1 U419 ( .A1(G237), .A2(G902), .ZN(n471) );
  NAND2_X1 U420 ( .A1(n638), .A2(n439), .ZN(n438) );
  NOR2_X1 U421 ( .A1(n638), .A2(n439), .ZN(n437) );
  INV_X1 U422 ( .A(KEYINPUT44), .ZN(n401) );
  XNOR2_X1 U423 ( .A(G902), .B(KEYINPUT15), .ZN(n599) );
  XOR2_X1 U424 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n527) );
  XNOR2_X1 U425 ( .A(G113), .B(G122), .ZN(n523) );
  XOR2_X1 U426 ( .A(KEYINPUT97), .B(KEYINPUT12), .Z(n524) );
  XNOR2_X1 U427 ( .A(n530), .B(n417), .ZN(n416) );
  INV_X1 U428 ( .A(KEYINPUT11), .ZN(n417) );
  XNOR2_X1 U429 ( .A(G143), .B(G104), .ZN(n530) );
  INV_X1 U430 ( .A(KEYINPUT30), .ZN(n394) );
  XNOR2_X1 U431 ( .A(n428), .B(n479), .ZN(n614) );
  XOR2_X1 U432 ( .A(KEYINPUT65), .B(KEYINPUT10), .Z(n494) );
  XNOR2_X1 U433 ( .A(n492), .B(G140), .ZN(n493) );
  XNOR2_X1 U434 ( .A(n694), .B(KEYINPUT70), .ZN(n452) );
  XNOR2_X1 U435 ( .A(n449), .B(n448), .ZN(n541) );
  INV_X1 U436 ( .A(KEYINPUT28), .ZN(n448) );
  XNOR2_X1 U437 ( .A(n365), .B(KEYINPUT39), .ZN(n563) );
  NAND2_X1 U438 ( .A1(n545), .A2(n537), .ZN(n365) );
  INV_X1 U439 ( .A(KEYINPUT107), .ZN(n450) );
  INV_X1 U440 ( .A(KEYINPUT6), .ZN(n373) );
  XNOR2_X1 U441 ( .A(n402), .B(n585), .ZN(n596) );
  NAND2_X1 U442 ( .A1(n691), .A2(G472), .ZN(n616) );
  INV_X2 U443 ( .A(G953), .ZN(n715) );
  NAND2_X1 U444 ( .A1(n691), .A2(G217), .ZN(n456) );
  INV_X1 U445 ( .A(G210), .ZN(n360) );
  XNOR2_X1 U446 ( .A(n446), .B(KEYINPUT47), .ZN(n445) );
  NAND2_X1 U447 ( .A1(n444), .A2(n442), .ZN(n446) );
  NOR2_X1 U448 ( .A1(n666), .A2(n443), .ZN(n442) );
  INV_X1 U449 ( .A(n447), .ZN(n443) );
  INV_X1 U450 ( .A(KEYINPUT48), .ZN(n439) );
  NOR2_X1 U451 ( .A1(n410), .A2(G237), .ZN(n525) );
  NOR2_X1 U452 ( .A1(n555), .A2(n624), .ZN(n666) );
  XNOR2_X1 U453 ( .A(n472), .B(KEYINPUT87), .ZN(n662) );
  XOR2_X1 U454 ( .A(KEYINPUT5), .B(KEYINPUT74), .Z(n476) );
  INV_X1 U455 ( .A(G125), .ZN(n404) );
  XNOR2_X1 U456 ( .A(G122), .B(G107), .ZN(n512) );
  XNOR2_X1 U457 ( .A(n458), .B(G143), .ZN(n451) );
  INV_X1 U458 ( .A(G128), .ZN(n458) );
  XNOR2_X1 U459 ( .A(G137), .B(G134), .ZN(n473) );
  XNOR2_X1 U460 ( .A(n425), .B(n492), .ZN(n465) );
  XNOR2_X1 U461 ( .A(n427), .B(n426), .ZN(n425) );
  XNOR2_X1 U462 ( .A(KEYINPUT86), .B(KEYINPUT82), .ZN(n427) );
  XNOR2_X1 U463 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n426) );
  NAND2_X1 U464 ( .A1(G237), .A2(G234), .ZN(n480) );
  INV_X1 U465 ( .A(KEYINPUT2), .ZN(n392) );
  AND2_X1 U466 ( .A1(n556), .A2(n597), .ZN(n449) );
  XNOR2_X1 U467 ( .A(n550), .B(KEYINPUT19), .ZN(n574) );
  AND2_X2 U468 ( .A1(n440), .A2(n353), .ZN(n389) );
  NAND2_X1 U469 ( .A1(n432), .A2(n430), .ZN(n440) );
  INV_X1 U470 ( .A(KEYINPUT45), .ZN(n441) );
  XNOR2_X1 U471 ( .A(G110), .B(G104), .ZN(n461) );
  XNOR2_X1 U472 ( .A(G128), .B(G110), .ZN(n495) );
  XNOR2_X1 U473 ( .A(G116), .B(G134), .ZN(n510) );
  XNOR2_X1 U474 ( .A(n408), .B(n355), .ZN(n382) );
  NAND2_X1 U475 ( .A1(n358), .A2(n357), .ZN(n408) );
  NOR2_X1 U476 ( .A1(n643), .A2(n420), .ZN(n358) );
  XNOR2_X1 U477 ( .A(n533), .B(n713), .ZN(n606) );
  XNOR2_X1 U478 ( .A(n486), .B(n400), .ZN(n399) );
  XNOR2_X1 U479 ( .A(KEYINPUT76), .B(KEYINPUT89), .ZN(n400) );
  XNOR2_X1 U480 ( .A(n395), .B(n394), .ZN(n393) );
  BUF_X1 U481 ( .A(n567), .Z(n413) );
  INV_X1 U482 ( .A(n574), .ZN(n447) );
  INV_X1 U483 ( .A(n551), .ZN(n444) );
  BUF_X1 U484 ( .A(G953), .Z(n410) );
  XNOR2_X1 U485 ( .A(n542), .B(KEYINPUT42), .ZN(n728) );
  XNOR2_X1 U486 ( .A(n536), .B(n535), .ZN(n726) );
  AND2_X1 U487 ( .A1(n414), .A2(n598), .ZN(n638) );
  XNOR2_X1 U488 ( .A(n415), .B(KEYINPUT36), .ZN(n414) );
  NOR2_X1 U489 ( .A1(n564), .A2(n413), .ZN(n415) );
  INV_X1 U490 ( .A(KEYINPUT35), .ZN(n371) );
  NAND2_X1 U491 ( .A1(n444), .A2(n447), .ZN(n631) );
  OR2_X1 U492 ( .A1(n596), .A2(n369), .ZN(n368) );
  NAND2_X1 U493 ( .A1(n376), .A2(n370), .ZN(n369) );
  NOR2_X1 U494 ( .A1(n598), .A2(n377), .ZN(n376) );
  XNOR2_X1 U495 ( .A(n586), .B(KEYINPUT104), .ZN(n729) );
  NOR2_X1 U496 ( .A1(n596), .A2(n364), .ZN(n586) );
  NAND2_X1 U497 ( .A1(n411), .A2(n351), .ZN(n364) );
  INV_X1 U498 ( .A(KEYINPUT63), .ZN(n423) );
  AND2_X1 U499 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U500 ( .A1(n454), .A2(n618), .ZN(n453) );
  XNOR2_X1 U501 ( .A(n456), .B(n455), .ZN(n454) );
  NOR2_X1 U502 ( .A1(n612), .A2(n693), .ZN(n412) );
  OR2_X1 U503 ( .A1(n693), .A2(n603), .ZN(n605) );
  AND2_X1 U504 ( .A1(G221), .A2(n518), .ZN(n349) );
  XOR2_X1 U505 ( .A(G119), .B(G137), .Z(n350) );
  NOR2_X1 U506 ( .A1(n592), .A2(n650), .ZN(n351) );
  AND2_X1 U507 ( .A1(n548), .A2(n544), .ZN(n352) );
  AND2_X1 U508 ( .A1(n569), .A2(n642), .ZN(n353) );
  BUF_X1 U509 ( .A(n648), .Z(n411) );
  XNOR2_X1 U510 ( .A(KEYINPUT34), .B(KEYINPUT77), .ZN(n354) );
  XNOR2_X1 U511 ( .A(KEYINPUT59), .B(KEYINPUT83), .ZN(n355) );
  INV_X1 U512 ( .A(G475), .ZN(n420) );
  XNOR2_X1 U513 ( .A(n356), .B(n474), .ZN(n428) );
  XNOR2_X2 U514 ( .A(n709), .B(G146), .ZN(n356) );
  INV_X1 U515 ( .A(n391), .ZN(n357) );
  NOR2_X2 U516 ( .A1(n391), .A2(n643), .ZN(n691) );
  NAND2_X1 U517 ( .A1(n359), .A2(n357), .ZN(n601) );
  NOR2_X1 U518 ( .A1(n643), .A2(n360), .ZN(n359) );
  XNOR2_X1 U519 ( .A(n361), .B(n371), .ZN(n723) );
  AND2_X1 U520 ( .A1(n723), .A2(n368), .ZN(n375) );
  XNOR2_X1 U521 ( .A(n595), .B(n354), .ZN(n372) );
  NAND2_X1 U522 ( .A1(n372), .A2(n352), .ZN(n361) );
  NAND2_X1 U523 ( .A1(n594), .A2(n584), .ZN(n402) );
  XNOR2_X1 U524 ( .A(n397), .B(KEYINPUT75), .ZN(n396) );
  NAND2_X1 U525 ( .A1(n507), .A2(n599), .ZN(n422) );
  AND2_X2 U526 ( .A1(n387), .A2(n392), .ZN(n643) );
  AND2_X2 U527 ( .A1(n393), .A2(n396), .ZN(n545) );
  NOR2_X1 U528 ( .A1(n582), .A2(n405), .ZN(n577) );
  XNOR2_X1 U529 ( .A(n362), .B(n401), .ZN(n435) );
  NAND2_X1 U530 ( .A1(n375), .A2(n725), .ZN(n362) );
  NAND2_X1 U531 ( .A1(n594), .A2(n678), .ZN(n595) );
  XNOR2_X2 U532 ( .A(n593), .B(KEYINPUT33), .ZN(n678) );
  XNOR2_X1 U533 ( .A(n496), .B(n350), .ZN(n409) );
  NAND2_X1 U534 ( .A1(n625), .A2(n633), .ZN(n363) );
  XNOR2_X2 U535 ( .A(n478), .B(n463), .ZN(n696) );
  XNOR2_X2 U536 ( .A(n383), .B(n386), .ZN(n478) );
  INV_X1 U537 ( .A(n389), .ZN(n714) );
  NAND2_X1 U538 ( .A1(n388), .A2(n389), .ZN(n387) );
  NOR2_X2 U539 ( .A1(n407), .A2(n647), .ZN(n506) );
  NAND2_X1 U540 ( .A1(n563), .A2(n555), .ZN(n536) );
  NOR2_X2 U541 ( .A1(G902), .A2(n692), .ZN(n504) );
  XNOR2_X1 U542 ( .A(n497), .B(n409), .ZN(n499) );
  XNOR2_X2 U543 ( .A(n367), .B(n473), .ZN(n709) );
  XNOR2_X1 U544 ( .A(n367), .B(n416), .ZN(n531) );
  XNOR2_X2 U545 ( .A(n418), .B(KEYINPUT66), .ZN(n367) );
  INV_X1 U546 ( .A(n368), .ZN(n628) );
  INV_X1 U547 ( .A(n597), .ZN(n370) );
  INV_X1 U548 ( .A(n650), .ZN(n377) );
  INV_X1 U549 ( .A(n382), .ZN(n379) );
  NAND2_X1 U550 ( .A1(n382), .A2(n606), .ZN(n381) );
  INV_X1 U551 ( .A(n704), .ZN(n388) );
  NAND2_X1 U552 ( .A1(n390), .A2(n389), .ZN(n644) );
  NAND2_X1 U553 ( .A1(n578), .A2(n538), .ZN(n397) );
  XNOR2_X1 U554 ( .A(n407), .B(KEYINPUT1), .ZN(n648) );
  XNOR2_X2 U555 ( .A(n489), .B(G469), .ZN(n407) );
  XNOR2_X2 U556 ( .A(n504), .B(n503), .ZN(n587) );
  XNOR2_X1 U557 ( .A(n403), .B(n713), .ZN(n692) );
  XNOR2_X1 U558 ( .A(n499), .B(n349), .ZN(n403) );
  XNOR2_X1 U559 ( .A(n619), .B(n423), .ZN(G57) );
  XNOR2_X1 U560 ( .A(n506), .B(n505), .ZN(n578) );
  NAND2_X1 U561 ( .A1(n431), .A2(n437), .ZN(n430) );
  XNOR2_X1 U562 ( .A(n412), .B(KEYINPUT120), .ZN(G54) );
  XNOR2_X2 U563 ( .A(G131), .B(KEYINPUT67), .ZN(n418) );
  XNOR2_X1 U564 ( .A(n429), .B(n457), .ZN(G60) );
  INV_X1 U565 ( .A(n562), .ZN(n431) );
  NAND2_X1 U566 ( .A1(n562), .A2(n439), .ZN(n433) );
  XNOR2_X1 U567 ( .A(n451), .B(n459), .ZN(n460) );
  XNOR2_X1 U568 ( .A(n513), .B(n451), .ZN(n514) );
  XNOR2_X2 U569 ( .A(n711), .B(G101), .ZN(n474) );
  XNOR2_X1 U570 ( .A(n453), .B(KEYINPUT123), .ZN(G66) );
  INV_X1 U571 ( .A(n692), .ZN(n455) );
  XNOR2_X1 U572 ( .A(n611), .B(n610), .ZN(n612) );
  INV_X1 U573 ( .A(n460), .ZN(n711) );
  XNOR2_X1 U574 ( .A(KEYINPUT60), .B(KEYINPUT121), .ZN(n457) );
  INV_X1 U575 ( .A(n641), .ZN(n569) );
  XNOR2_X1 U576 ( .A(n614), .B(n613), .ZN(n615) );
  XNOR2_X1 U577 ( .A(n609), .B(n608), .ZN(n610) );
  XNOR2_X1 U578 ( .A(n616), .B(n615), .ZN(n617) );
  INV_X1 U579 ( .A(KEYINPUT40), .ZN(n535) );
  NOR2_X1 U580 ( .A1(G952), .A2(n715), .ZN(n693) );
  XNOR2_X1 U581 ( .A(n605), .B(n604), .ZN(G51) );
  XNOR2_X1 U582 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n459) );
  XNOR2_X1 U583 ( .A(n461), .B(KEYINPUT84), .ZN(n694) );
  NAND2_X1 U584 ( .A1(G224), .A2(n715), .ZN(n464) );
  XNOR2_X1 U585 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U586 ( .A(KEYINPUT55), .B(KEYINPUT54), .Z(n469) );
  XNOR2_X1 U587 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n468) );
  XNOR2_X1 U588 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U589 ( .A(n507), .B(n470), .ZN(n602) );
  XNOR2_X1 U590 ( .A(n471), .B(KEYINPUT73), .ZN(n508) );
  NAND2_X1 U591 ( .A1(n508), .A2(G214), .ZN(n472) );
  INV_X1 U592 ( .A(n662), .ZN(n560) );
  NAND2_X1 U593 ( .A1(n525), .A2(G210), .ZN(n475) );
  XNOR2_X1 U594 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U595 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U596 ( .A(n480), .B(KEYINPUT14), .ZN(n481) );
  NAND2_X1 U597 ( .A1(G952), .A2(n481), .ZN(n677) );
  NOR2_X1 U598 ( .A1(n410), .A2(n677), .ZN(n572) );
  NAND2_X1 U599 ( .A1(G902), .A2(n481), .ZN(n482) );
  XOR2_X1 U600 ( .A(KEYINPUT88), .B(n482), .Z(n483) );
  NAND2_X1 U601 ( .A1(n410), .A2(n483), .ZN(n570) );
  NOR2_X1 U602 ( .A1(G900), .A2(n570), .ZN(n484) );
  NOR2_X1 U603 ( .A1(n572), .A2(n484), .ZN(n485) );
  XOR2_X1 U604 ( .A(KEYINPUT78), .B(n485), .Z(n538) );
  NAND2_X1 U605 ( .A1(G227), .A2(n715), .ZN(n486) );
  NAND2_X1 U606 ( .A1(G234), .A2(n599), .ZN(n490) );
  XNOR2_X1 U607 ( .A(KEYINPUT20), .B(n490), .ZN(n500) );
  NAND2_X1 U608 ( .A1(n500), .A2(G221), .ZN(n491) );
  XNOR2_X1 U609 ( .A(KEYINPUT21), .B(n491), .ZN(n651) );
  XOR2_X1 U610 ( .A(KEYINPUT92), .B(n651), .Z(n583) );
  XNOR2_X1 U611 ( .A(n494), .B(n493), .ZN(n713) );
  XNOR2_X1 U612 ( .A(n495), .B(KEYINPUT90), .ZN(n497) );
  XOR2_X1 U613 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n496) );
  NAND2_X1 U614 ( .A1(G234), .A2(n715), .ZN(n498) );
  XOR2_X1 U615 ( .A(KEYINPUT8), .B(n498), .Z(n518) );
  XOR2_X1 U616 ( .A(KEYINPUT91), .B(KEYINPUT25), .Z(n502) );
  NAND2_X1 U617 ( .A1(n500), .A2(G217), .ZN(n501) );
  XNOR2_X1 U618 ( .A(n502), .B(n501), .ZN(n503) );
  NAND2_X1 U619 ( .A1(G210), .A2(n508), .ZN(n509) );
  XNOR2_X1 U620 ( .A(KEYINPUT38), .B(n567), .ZN(n537) );
  XNOR2_X1 U621 ( .A(KEYINPUT103), .B(G478), .ZN(n522) );
  XOR2_X1 U622 ( .A(KEYINPUT101), .B(KEYINPUT7), .Z(n511) );
  XNOR2_X1 U623 ( .A(n511), .B(n510), .ZN(n517) );
  XOR2_X1 U624 ( .A(KEYINPUT102), .B(KEYINPUT9), .Z(n515) );
  INV_X1 U625 ( .A(n512), .ZN(n513) );
  XNOR2_X1 U626 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U627 ( .A(n517), .B(n516), .Z(n520) );
  NAND2_X1 U628 ( .A1(G217), .A2(n518), .ZN(n519) );
  XNOR2_X1 U629 ( .A(n520), .B(n519), .ZN(n688) );
  NOR2_X1 U630 ( .A1(G902), .A2(n688), .ZN(n521) );
  XNOR2_X1 U631 ( .A(n522), .B(n521), .ZN(n544) );
  INV_X1 U632 ( .A(n544), .ZN(n549) );
  XNOR2_X1 U633 ( .A(n524), .B(n523), .ZN(n529) );
  NAND2_X1 U634 ( .A1(n525), .A2(G214), .ZN(n526) );
  XNOR2_X1 U635 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U636 ( .A(n529), .B(n528), .ZN(n532) );
  XNOR2_X1 U637 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U638 ( .A(KEYINPUT13), .B(KEYINPUT100), .ZN(n534) );
  NAND2_X1 U639 ( .A1(n549), .A2(n548), .ZN(n634) );
  INV_X1 U640 ( .A(n634), .ZN(n555) );
  INV_X1 U641 ( .A(n537), .ZN(n663) );
  NOR2_X1 U642 ( .A1(n662), .A2(n663), .ZN(n667) );
  NOR2_X1 U643 ( .A1(n544), .A2(n548), .ZN(n664) );
  INV_X1 U644 ( .A(n587), .ZN(n650) );
  NAND2_X1 U645 ( .A1(n650), .A2(n538), .ZN(n539) );
  NOR2_X1 U646 ( .A1(n651), .A2(n539), .ZN(n556) );
  XOR2_X1 U647 ( .A(n407), .B(KEYINPUT111), .Z(n540) );
  XNOR2_X1 U648 ( .A(n543), .B(KEYINPUT46), .ZN(n554) );
  NAND2_X1 U649 ( .A1(n545), .A2(n352), .ZN(n546) );
  NOR2_X1 U650 ( .A1(n546), .A2(n413), .ZN(n547) );
  XNOR2_X1 U651 ( .A(n547), .B(KEYINPUT110), .ZN(n727) );
  NOR2_X1 U652 ( .A1(n549), .A2(n548), .ZN(n624) );
  XNOR2_X1 U653 ( .A(n552), .B(KEYINPUT72), .ZN(n553) );
  NAND2_X1 U654 ( .A1(n554), .A2(n553), .ZN(n562) );
  INV_X1 U655 ( .A(n592), .ZN(n558) );
  NAND2_X1 U656 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U657 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U658 ( .A(KEYINPUT108), .B(n559), .ZN(n561) );
  NAND2_X1 U659 ( .A1(n561), .A2(n560), .ZN(n564) );
  AND2_X1 U660 ( .A1(n563), .A2(n624), .ZN(n641) );
  XOR2_X1 U661 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n566) );
  INV_X1 U662 ( .A(n411), .ZN(n598) );
  OR2_X1 U663 ( .A1(n564), .A2(n598), .ZN(n565) );
  XNOR2_X1 U664 ( .A(n566), .B(n565), .ZN(n568) );
  NAND2_X1 U665 ( .A1(n568), .A2(n413), .ZN(n642) );
  NOR2_X1 U666 ( .A1(G898), .A2(n570), .ZN(n571) );
  NOR2_X1 U667 ( .A1(n572), .A2(n571), .ZN(n573) );
  INV_X1 U668 ( .A(KEYINPUT0), .ZN(n575) );
  NAND2_X1 U669 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U670 ( .A1(n648), .A2(n647), .ZN(n591) );
  NOR2_X1 U671 ( .A1(n657), .A2(n582), .ZN(n581) );
  XNOR2_X1 U672 ( .A(n581), .B(KEYINPUT31), .ZN(n633) );
  XOR2_X1 U673 ( .A(KEYINPUT22), .B(KEYINPUT71), .Z(n585) );
  AND2_X1 U674 ( .A1(n664), .A2(n583), .ZN(n584) );
  NOR2_X1 U675 ( .A1(n411), .A2(n587), .ZN(n588) );
  XNOR2_X1 U676 ( .A(KEYINPUT106), .B(n588), .ZN(n589) );
  NAND2_X1 U677 ( .A1(n592), .A2(n591), .ZN(n593) );
  INV_X1 U678 ( .A(n599), .ZN(n600) );
  XNOR2_X1 U679 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U680 ( .A(KEYINPUT119), .B(KEYINPUT56), .ZN(n604) );
  INV_X1 U681 ( .A(n606), .ZN(n607) );
  INV_X1 U682 ( .A(n693), .ZN(n618) );
  NAND2_X1 U683 ( .A1(n691), .A2(G469), .ZN(n611) );
  XOR2_X1 U684 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n608) );
  XOR2_X1 U685 ( .A(KEYINPUT62), .B(KEYINPUT112), .Z(n613) );
  NOR2_X1 U686 ( .A1(n625), .A2(n634), .ZN(n621) );
  XNOR2_X1 U687 ( .A(G104), .B(KEYINPUT113), .ZN(n620) );
  XNOR2_X1 U688 ( .A(n621), .B(n620), .ZN(G6) );
  XOR2_X1 U689 ( .A(KEYINPUT26), .B(KEYINPUT114), .Z(n623) );
  XNOR2_X1 U690 ( .A(G107), .B(KEYINPUT27), .ZN(n622) );
  XNOR2_X1 U691 ( .A(n623), .B(n622), .ZN(n627) );
  INV_X1 U692 ( .A(n624), .ZN(n636) );
  NOR2_X1 U693 ( .A1(n625), .A2(n636), .ZN(n626) );
  XOR2_X1 U694 ( .A(n627), .B(n626), .Z(G9) );
  XOR2_X1 U695 ( .A(G110), .B(n628), .Z(G12) );
  NOR2_X1 U696 ( .A1(n636), .A2(n631), .ZN(n630) );
  XNOR2_X1 U697 ( .A(G128), .B(KEYINPUT29), .ZN(n629) );
  XNOR2_X1 U698 ( .A(n630), .B(n629), .ZN(G30) );
  NOR2_X1 U699 ( .A1(n634), .A2(n631), .ZN(n632) );
  XOR2_X1 U700 ( .A(G146), .B(n632), .Z(G48) );
  NOR2_X1 U701 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U702 ( .A(G113), .B(n635), .Z(G15) );
  NOR2_X1 U703 ( .A1(n636), .A2(n633), .ZN(n637) );
  XOR2_X1 U704 ( .A(G116), .B(n637), .Z(G18) );
  XOR2_X1 U705 ( .A(KEYINPUT115), .B(KEYINPUT37), .Z(n640) );
  XNOR2_X1 U706 ( .A(G125), .B(n638), .ZN(n639) );
  XNOR2_X1 U707 ( .A(n640), .B(n639), .ZN(G27) );
  XOR2_X1 U708 ( .A(G134), .B(n641), .Z(G36) );
  XNOR2_X1 U709 ( .A(G140), .B(n642), .ZN(G42) );
  XNOR2_X1 U710 ( .A(n643), .B(KEYINPUT79), .ZN(n646) );
  BUF_X1 U711 ( .A(n644), .Z(n645) );
  NAND2_X1 U712 ( .A1(n646), .A2(n645), .ZN(n684) );
  NAND2_X1 U713 ( .A1(n411), .A2(n647), .ZN(n649) );
  XNOR2_X1 U714 ( .A(n649), .B(KEYINPUT50), .ZN(n656) );
  AND2_X1 U715 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U716 ( .A(KEYINPUT49), .B(n652), .Z(n653) );
  NOR2_X1 U717 ( .A1(n405), .A2(n653), .ZN(n655) );
  NAND2_X1 U718 ( .A1(n656), .A2(n655), .ZN(n658) );
  NAND2_X1 U719 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U720 ( .A(KEYINPUT51), .B(n659), .ZN(n660) );
  NOR2_X1 U721 ( .A1(n679), .A2(n660), .ZN(n661) );
  XOR2_X1 U722 ( .A(KEYINPUT116), .B(n661), .Z(n674) );
  NAND2_X1 U723 ( .A1(n663), .A2(n662), .ZN(n665) );
  NAND2_X1 U724 ( .A1(n665), .A2(n664), .ZN(n670) );
  NAND2_X1 U725 ( .A1(n667), .A2(n344), .ZN(n668) );
  XOR2_X1 U726 ( .A(KEYINPUT117), .B(n668), .Z(n669) );
  NAND2_X1 U727 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U728 ( .A(KEYINPUT118), .B(n671), .ZN(n672) );
  NAND2_X1 U729 ( .A1(n672), .A2(n678), .ZN(n673) );
  NAND2_X1 U730 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U731 ( .A(KEYINPUT52), .B(n675), .Z(n676) );
  NOR2_X1 U732 ( .A1(n677), .A2(n676), .ZN(n682) );
  INV_X1 U733 ( .A(n678), .ZN(n680) );
  NOR2_X1 U734 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U735 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U736 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U737 ( .A1(n685), .A2(n410), .ZN(n686) );
  XNOR2_X1 U738 ( .A(n686), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U739 ( .A1(n691), .A2(G478), .ZN(n687) );
  XNOR2_X1 U740 ( .A(n687), .B(KEYINPUT122), .ZN(n689) );
  XNOR2_X1 U741 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U742 ( .A1(n693), .A2(n690), .ZN(G63) );
  XOR2_X1 U743 ( .A(n694), .B(KEYINPUT125), .Z(n695) );
  XNOR2_X1 U744 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U745 ( .A(n697), .B(G101), .ZN(n699) );
  NOR2_X1 U746 ( .A1(n715), .A2(G898), .ZN(n698) );
  NOR2_X1 U747 ( .A1(n699), .A2(n698), .ZN(n708) );
  XOR2_X1 U748 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n701) );
  NAND2_X1 U749 ( .A1(G224), .A2(n410), .ZN(n700) );
  XNOR2_X1 U750 ( .A(n701), .B(n700), .ZN(n703) );
  INV_X1 U751 ( .A(G898), .ZN(n702) );
  NOR2_X1 U752 ( .A1(n703), .A2(n702), .ZN(n706) );
  NOR2_X1 U753 ( .A1(n410), .A2(n704), .ZN(n705) );
  NOR2_X1 U754 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U755 ( .A(n708), .B(n707), .Z(G69) );
  XOR2_X1 U756 ( .A(n709), .B(KEYINPUT126), .Z(n710) );
  XNOR2_X1 U757 ( .A(n711), .B(n710), .ZN(n712) );
  XOR2_X1 U758 ( .A(n713), .B(n712), .Z(n717) );
  XOR2_X1 U759 ( .A(n717), .B(n714), .Z(n716) );
  NAND2_X1 U760 ( .A1(n716), .A2(n715), .ZN(n722) );
  XNOR2_X1 U761 ( .A(n717), .B(G227), .ZN(n718) );
  XNOR2_X1 U762 ( .A(n718), .B(KEYINPUT127), .ZN(n719) );
  NAND2_X1 U763 ( .A1(n719), .A2(G900), .ZN(n720) );
  NAND2_X1 U764 ( .A1(n410), .A2(n720), .ZN(n721) );
  NAND2_X1 U765 ( .A1(n722), .A2(n721), .ZN(G72) );
  BUF_X1 U766 ( .A(n723), .Z(n724) );
  XNOR2_X1 U767 ( .A(G122), .B(n724), .ZN(G24) );
  XNOR2_X1 U768 ( .A(G119), .B(n725), .ZN(G21) );
  XOR2_X1 U769 ( .A(n726), .B(G131), .Z(G33) );
  XOR2_X1 U770 ( .A(G143), .B(n727), .Z(G45) );
  XOR2_X1 U771 ( .A(n728), .B(G137), .Z(G39) );
  XOR2_X1 U772 ( .A(G101), .B(n729), .Z(G3) );
endmodule

