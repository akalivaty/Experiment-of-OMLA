//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 1 1 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT65), .Z(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  INV_X1    g0016(.A(new_n201), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(new_n213), .A2(new_n214), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n211), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n220), .B1(new_n214), .B2(new_n213), .C1(new_n227), .C2(KEYINPUT1), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  AND2_X1   g0044(.A1(KEYINPUT3), .A2(G33), .ZN(new_n245));
  NOR2_X1   g0045(.A1(KEYINPUT3), .A2(G33), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n247), .A2(G1698), .ZN(new_n248));
  AOI22_X1  g0048(.A1(new_n248), .A2(G222), .B1(G77), .B2(new_n247), .ZN(new_n249));
  INV_X1    g0049(.A(G223), .ZN(new_n250));
  OR2_X1    g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G1698), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n249), .B1(new_n250), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  INV_X1    g0058(.A(G45), .ZN(new_n259));
  AOI21_X1  g0059(.A(G1), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n260), .A2(G274), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n256), .A2(new_n260), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n261), .B1(new_n262), .B2(G226), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G190), .ZN(new_n265));
  AOI21_X1  g0065(.A(G200), .B1(new_n257), .B2(new_n263), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n215), .ZN(new_n269));
  XOR2_X1   g0069(.A(KEYINPUT8), .B(G58), .Z(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT66), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT8), .B(G58), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT66), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n271), .A2(new_n274), .A3(new_n209), .A4(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G150), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(KEYINPUT67), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n204), .A2(G20), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(KEYINPUT67), .B1(new_n275), .B2(new_n277), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n269), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(new_n269), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n209), .A2(G1), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(new_n202), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n285), .A2(new_n287), .B1(new_n202), .B2(new_n284), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n282), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT9), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT9), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n282), .A2(new_n291), .A3(new_n288), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n267), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT10), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT73), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n267), .A2(KEYINPUT10), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n282), .A2(new_n291), .A3(new_n288), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n291), .B1(new_n282), .B2(new_n288), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT72), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT72), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(new_n290), .B2(new_n292), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n296), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT73), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n297), .A2(new_n298), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n303), .B(KEYINPUT10), .C1(new_n304), .C2(new_n267), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n295), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n264), .A2(G169), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n307), .B1(new_n308), .B2(new_n264), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n289), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n248), .A2(G232), .B1(G107), .B2(new_n247), .ZN(new_n311));
  INV_X1    g0111(.A(G238), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n311), .B1(new_n312), .B2(new_n254), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n256), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n261), .B1(new_n262), .B2(G244), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G200), .ZN(new_n317));
  INV_X1    g0117(.A(new_n276), .ZN(new_n318));
  INV_X1    g0118(.A(G77), .ZN(new_n319));
  OAI22_X1  g0119(.A1(new_n272), .A2(new_n318), .B1(new_n209), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT68), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n209), .A2(G33), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT15), .B(G87), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n320), .A2(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n320), .A2(new_n321), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n269), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n284), .A2(KEYINPUT69), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT69), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n283), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(G77), .ZN(new_n331));
  INV_X1    g0131(.A(new_n330), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n332), .A2(new_n269), .A3(new_n286), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n331), .B1(new_n333), .B2(G77), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n317), .A2(KEYINPUT70), .A3(new_n326), .A4(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT70), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n326), .ZN(new_n337));
  INV_X1    g0137(.A(G200), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n338), .B1(new_n314), .B2(new_n315), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n336), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n316), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G190), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n335), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G169), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n316), .A2(new_n308), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n337), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT71), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n343), .A2(KEYINPUT71), .A3(new_n347), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n306), .A2(new_n310), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT74), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n306), .A2(KEYINPUT74), .A3(new_n310), .A4(new_n352), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n318), .A2(new_n202), .B1(new_n209), .B2(G68), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n322), .A2(new_n319), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n269), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XOR2_X1   g0159(.A(new_n359), .B(KEYINPUT11), .Z(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(G68), .B2(new_n333), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n283), .A2(KEYINPUT12), .A3(G68), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT12), .B1(new_n330), .B2(G68), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n362), .B1(new_n363), .B2(KEYINPUT77), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(KEYINPUT77), .B2(new_n363), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT13), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n261), .B1(new_n262), .B2(G238), .ZN(new_n368));
  INV_X1    g0168(.A(G1698), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n253), .A2(G226), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n253), .A2(G232), .A3(G1698), .ZN(new_n371));
  NAND2_X1  g0171(.A1(G33), .A2(G97), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT75), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT75), .A4(new_n372), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n256), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n367), .B(new_n368), .C1(new_n375), .C2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT76), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n373), .A2(new_n374), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n381), .A2(new_n256), .A3(new_n376), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n368), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT13), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n382), .A2(KEYINPUT76), .A3(new_n367), .A4(new_n368), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n380), .A2(new_n384), .A3(G190), .A4(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n378), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n367), .B1(new_n382), .B2(new_n368), .ZN(new_n388));
  OAI21_X1  g0188(.A(G200), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n366), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(KEYINPUT78), .A2(G169), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n387), .B2(new_n388), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT14), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n380), .A2(new_n384), .A3(G179), .A4(new_n385), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT14), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n395), .B(new_n391), .C1(new_n387), .C2(new_n388), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n393), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n366), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n390), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n271), .A2(new_n274), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n286), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n285), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n400), .A2(new_n284), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT79), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT7), .B1(new_n247), .B2(new_n209), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT7), .ZN(new_n408));
  NOR4_X1   g0208(.A1(new_n245), .A2(new_n246), .A3(new_n408), .A4(G20), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n406), .B(G68), .C1(new_n407), .C2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(G58), .ZN(new_n411));
  INV_X1    g0211(.A(G68), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(G20), .B1(new_n413), .B2(new_n201), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n276), .A2(G159), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n410), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n251), .A2(new_n209), .A3(new_n252), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n408), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n247), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n406), .B1(new_n422), .B2(G68), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT16), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n418), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n412), .B1(new_n420), .B2(new_n421), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n424), .B1(new_n426), .B2(new_n416), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n269), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n405), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(G223), .B(new_n369), .C1(new_n245), .C2(new_n246), .ZN(new_n430));
  OAI211_X1 g0230(.A(G226), .B(G1698), .C1(new_n245), .C2(new_n246), .ZN(new_n431));
  INV_X1    g0231(.A(G33), .ZN(new_n432));
  INV_X1    g0232(.A(G87), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n430), .B(new_n431), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n256), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n261), .B1(new_n262), .B2(G232), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n437), .A2(G179), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n438), .B1(new_n344), .B2(new_n437), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n429), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT18), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n440), .B(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n403), .A2(new_n404), .ZN(new_n443));
  INV_X1    g0243(.A(new_n269), .ZN(new_n444));
  OAI21_X1  g0244(.A(G68), .B1(new_n407), .B2(new_n409), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n417), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n444), .B1(new_n446), .B2(new_n424), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(KEYINPUT79), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n448), .A2(KEYINPUT16), .A3(new_n410), .A4(new_n417), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n443), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n437), .A2(new_n338), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(G190), .B2(new_n437), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n453), .B(KEYINPUT17), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n399), .A2(new_n442), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n355), .A2(new_n356), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(G250), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n459), .B1(new_n208), .B2(G45), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n208), .A2(G45), .A3(G274), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n256), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G116), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n432), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n253), .A2(G244), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n465), .B1(new_n466), .B2(G1698), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n253), .A2(new_n369), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT81), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n468), .A2(new_n469), .A3(new_n312), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT81), .B1(new_n248), .B2(G238), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n463), .B1(new_n472), .B2(new_n256), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n332), .A2(new_n323), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n253), .A2(new_n209), .A3(G68), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT19), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n209), .B1(new_n372), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G97), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n433), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(G107), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n476), .B1(new_n372), .B2(G20), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n475), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n269), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n474), .A2(new_n483), .ZN(new_n484));
  XOR2_X1   g0284(.A(new_n323), .B(KEYINPUT82), .Z(new_n485));
  NAND2_X1  g0285(.A1(new_n208), .A2(G33), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(new_n285), .A3(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n473), .A2(new_n308), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n463), .ZN(new_n489));
  INV_X1    g0289(.A(new_n465), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n253), .A2(G244), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n490), .B1(new_n491), .B2(new_n369), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n469), .B1(new_n468), .B2(new_n312), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n248), .A2(KEYINPUT81), .A3(G238), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n256), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n489), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n344), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n488), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n283), .A2(new_n486), .A3(new_n215), .A4(new_n268), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n474), .B(new_n483), .C1(new_n433), .C2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n501), .B1(new_n497), .B2(G200), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT83), .B1(new_n473), .B2(G190), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n493), .A2(new_n494), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n496), .B1(new_n504), .B2(new_n467), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT83), .ZN(new_n506));
  INV_X1    g0306(.A(G190), .ZN(new_n507));
  NOR4_X1   g0307(.A1(new_n505), .A2(new_n506), .A3(new_n507), .A4(new_n463), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n502), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n466), .A2(KEYINPUT4), .A3(new_n369), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT4), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n491), .A2(new_n511), .B1(G33), .B2(G283), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT4), .B1(new_n247), .B2(new_n459), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G1698), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n510), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n256), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT5), .ZN(new_n517));
  AOI211_X1 g0317(.A(G1), .B(new_n259), .C1(new_n517), .C2(G41), .ZN(new_n518));
  OR3_X1    g0318(.A1(new_n517), .A2(KEYINPUT80), .A3(G41), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT80), .B1(new_n517), .B2(G41), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(G257), .A3(new_n496), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n518), .A2(G274), .A3(new_n519), .A4(new_n520), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n516), .A2(new_n525), .A3(G179), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n344), .B1(new_n516), .B2(new_n525), .ZN(new_n527));
  INV_X1    g0327(.A(G107), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n528), .A2(KEYINPUT6), .A3(G97), .ZN(new_n529));
  XOR2_X1   g0329(.A(G97), .B(G107), .Z(new_n530));
  OAI21_X1  g0330(.A(new_n529), .B1(new_n530), .B2(KEYINPUT6), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n531), .A2(G20), .B1(G77), .B2(new_n276), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n422), .A2(G107), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n444), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n284), .A2(new_n478), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n500), .B2(new_n478), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n526), .A2(new_n527), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n534), .A2(new_n536), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n516), .A2(new_n525), .A3(new_n507), .ZN(new_n539));
  AOI21_X1  g0339(.A(G200), .B1(new_n516), .B2(new_n525), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND4_X1   g0341(.A1(new_n499), .A2(new_n509), .A3(new_n537), .A4(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n209), .A2(G107), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT23), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT23), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n209), .B2(G107), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n544), .A2(new_n546), .B1(new_n209), .B2(new_n465), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n253), .A2(new_n209), .A3(G87), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT22), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT22), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n253), .A2(new_n551), .A3(new_n209), .A4(G87), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n548), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n444), .B1(new_n553), .B2(KEYINPUT24), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n550), .A2(new_n552), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n547), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT24), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(G13), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n559), .A2(G1), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n543), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT25), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT25), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n560), .A2(new_n543), .A3(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n562), .B(new_n564), .C1(new_n528), .C2(new_n500), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT84), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OR2_X1    g0367(.A1(new_n565), .A2(new_n566), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n554), .A2(new_n558), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n253), .A2(G250), .A3(new_n369), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n253), .A2(G257), .A3(G1698), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G33), .A2(G294), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n256), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n521), .A2(G264), .A3(new_n496), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n574), .A2(new_n507), .A3(new_n575), .A4(new_n523), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n523), .A3(new_n575), .ZN(new_n577));
  AOI22_X1  g0377(.A1(KEYINPUT86), .A2(new_n576), .B1(new_n577), .B2(new_n338), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n577), .A2(KEYINPUT86), .A3(new_n338), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n569), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n568), .A2(new_n567), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n269), .B1(new_n556), .B2(new_n557), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n553), .A2(KEYINPUT24), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT85), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n574), .A2(G179), .A3(new_n575), .A4(new_n523), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n585), .A2(new_n586), .B1(new_n577), .B2(G169), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n577), .A2(new_n585), .A3(G169), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n584), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n580), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n253), .A2(G264), .A3(G1698), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n253), .A2(G257), .A3(new_n369), .ZN(new_n592));
  INV_X1    g0392(.A(G303), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n591), .B(new_n592), .C1(new_n593), .C2(new_n253), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n594), .A2(new_n256), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n521), .A2(G270), .A3(new_n496), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n523), .ZN(new_n597));
  OAI211_X1 g0397(.A(KEYINPUT21), .B(G169), .C1(new_n595), .C2(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n596), .A2(new_n523), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n594), .A2(new_n256), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(G179), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n330), .A2(G116), .A3(new_n444), .A4(new_n486), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(G116), .B2(new_n330), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n432), .A2(G97), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G33), .A2(G283), .ZN(new_n606));
  AOI21_X1  g0406(.A(G20), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n209), .A2(new_n464), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n269), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g0409(.A(new_n609), .B(KEYINPUT20), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n602), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n600), .A2(new_n523), .A3(new_n596), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n614), .B(G169), .C1(new_n610), .C2(new_n604), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT21), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(G200), .B1(new_n599), .B2(new_n600), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n595), .A2(new_n597), .A3(G190), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n611), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n613), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n590), .A2(new_n621), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n458), .A2(new_n542), .A3(new_n622), .ZN(G372));
  NAND2_X1  g0423(.A1(new_n516), .A2(new_n525), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(G169), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n524), .B1(new_n256), .B2(new_n515), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(G179), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n538), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  AND4_X1   g0428(.A1(KEYINPUT26), .A2(new_n509), .A3(new_n499), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT87), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT87), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n509), .A2(new_n628), .A3(new_n499), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n630), .B1(new_n629), .B2(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n537), .A2(new_n541), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n602), .A2(new_n612), .B1(new_n615), .B2(new_n616), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n589), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n506), .B1(new_n497), .B2(new_n507), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n473), .A2(KEYINPUT83), .A3(G190), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n641), .A2(new_n502), .B1(new_n498), .B2(new_n488), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n636), .A2(new_n638), .A3(new_n642), .A4(new_n580), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n643), .A2(new_n499), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n635), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n458), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT17), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n453), .B(new_n647), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n390), .A2(new_n347), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n397), .A2(new_n398), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n440), .B(KEYINPUT18), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n306), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n310), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n646), .A2(new_n655), .ZN(G369));
  NAND2_X1  g0456(.A1(new_n560), .A2(new_n209), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n659), .A3(G213), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n611), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(new_n637), .B2(new_n620), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n665), .B1(new_n637), .B2(new_n664), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n589), .A2(new_n663), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n580), .B(new_n589), .C1(new_n569), .C2(new_n663), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n637), .A2(new_n662), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(new_n669), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n589), .B2(new_n662), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n671), .A2(new_n674), .ZN(G399));
  INV_X1    g0475(.A(new_n212), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(G41), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n479), .A2(G107), .A3(G116), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G1), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n218), .B2(new_n678), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT28), .ZN(new_n682));
  AOI21_X1  g0482(.A(KEYINPUT26), .B1(new_n642), .B2(new_n628), .ZN(new_n683));
  OAI211_X1 g0483(.A(new_n643), .B(new_n499), .C1(new_n683), .C2(new_n629), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n684), .A2(KEYINPUT29), .A3(new_n663), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n645), .A2(new_n663), .ZN(new_n686));
  XOR2_X1   g0486(.A(KEYINPUT88), .B(KEYINPUT29), .Z(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n685), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G330), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT31), .ZN(new_n691));
  AOI21_X1  g0491(.A(G179), .B1(new_n599), .B2(new_n600), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n692), .A2(new_n624), .A3(new_n497), .A4(new_n577), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n614), .A2(new_n308), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n574), .A2(new_n575), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n694), .A2(new_n473), .A3(new_n626), .A4(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n693), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n624), .A2(new_n601), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n473), .A2(new_n695), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT30), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n691), .B(new_n662), .C1(new_n698), .C2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n542), .A2(new_n622), .A3(new_n663), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n696), .A2(new_n697), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n699), .A2(new_n700), .A3(KEYINPUT30), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(new_n706), .A3(new_n693), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n691), .B1(new_n707), .B2(new_n662), .ZN(new_n708));
  AOI211_X1 g0508(.A(new_n690), .B(new_n703), .C1(new_n704), .C2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n689), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n682), .B1(new_n710), .B2(G1), .ZN(G364));
  NOR2_X1   g0511(.A1(new_n559), .A2(G20), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G45), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n678), .A2(G1), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n676), .A2(new_n247), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n715), .A2(G355), .B1(new_n464), .B2(new_n676), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n212), .A2(new_n247), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT90), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n219), .A2(G45), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n719), .B1(new_n240), .B2(G45), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n716), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G13), .A2(G33), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G20), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n215), .B1(G20), .B2(new_n344), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n714), .B1(new_n721), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n725), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n308), .A2(new_n338), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n209), .A2(new_n507), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n507), .A2(G179), .A3(G200), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n209), .ZN(new_n733));
  OAI221_X1 g0533(.A(new_n253), .B1(new_n731), .B2(new_n202), .C1(new_n733), .C2(new_n478), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n338), .A2(G179), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n209), .A2(G190), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n308), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI22_X1  g0541(.A1(G87), .A2(new_n737), .B1(new_n741), .B2(G77), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n729), .A2(new_n738), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n738), .A2(new_n735), .ZN(new_n744));
  OAI221_X1 g0544(.A(new_n742), .B1(new_n412), .B2(new_n743), .C1(new_n528), .C2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n730), .A2(new_n739), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT91), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n746), .A2(new_n747), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n734), .B(new_n745), .C1(G58), .C2(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n738), .A2(new_n308), .A3(new_n338), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n754), .A2(KEYINPUT92), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(KEYINPUT92), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(KEYINPUT93), .B(G159), .Z(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT32), .ZN(new_n760));
  INV_X1    g0560(.A(new_n731), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n253), .B1(new_n761), .B2(G326), .ZN(new_n762));
  INV_X1    g0562(.A(G294), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n762), .B1(new_n763), .B2(new_n733), .ZN(new_n764));
  XOR2_X1   g0564(.A(KEYINPUT33), .B(G317), .Z(new_n765));
  INV_X1    g0565(.A(G311), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n765), .A2(new_n743), .B1(new_n740), .B2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G283), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n736), .A2(new_n593), .B1(new_n744), .B2(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n764), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n757), .ZN(new_n771));
  AOI22_X1  g0571(.A1(G322), .A2(new_n752), .B1(new_n771), .B2(G329), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n753), .A2(new_n760), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n724), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n727), .B1(new_n728), .B2(new_n773), .C1(new_n666), .C2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n714), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n666), .A2(G330), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n776), .B1(new_n777), .B2(KEYINPUT89), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n777), .B1(KEYINPUT89), .B2(new_n667), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n775), .B1(new_n779), .B2(new_n780), .ZN(G396));
  AOI21_X1  g0581(.A(new_n247), .B1(new_n737), .B2(G50), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n782), .B1(new_n411), .B2(new_n733), .C1(new_n412), .C2(new_n744), .ZN(new_n783));
  INV_X1    g0583(.A(new_n758), .ZN(new_n784));
  AOI22_X1  g0584(.A1(G137), .A2(new_n761), .B1(new_n784), .B2(new_n741), .ZN(new_n785));
  INV_X1    g0585(.A(G150), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n785), .B1(new_n786), .B2(new_n743), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(G143), .B2(new_n752), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT34), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n783), .B(new_n789), .C1(G132), .C2(new_n771), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n247), .B1(new_n736), .B2(new_n528), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT94), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n792), .B1(new_n763), .B2(new_n751), .C1(new_n766), .C2(new_n757), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n733), .A2(new_n478), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n731), .A2(new_n593), .B1(new_n740), .B2(new_n464), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n743), .A2(new_n768), .B1(new_n744), .B2(new_n433), .ZN(new_n796));
  NOR4_X1   g0596(.A1(new_n793), .A2(new_n794), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n725), .B1(new_n790), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n725), .A2(new_n722), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n714), .B1(new_n319), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n337), .A2(new_n662), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n343), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n347), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n347), .A2(new_n662), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n798), .B(new_n800), .C1(new_n807), .C2(new_n723), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT95), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n686), .A2(new_n806), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n662), .B1(new_n635), .B2(new_n644), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n807), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n703), .B1(new_n704), .B2(new_n708), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G330), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n714), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n813), .A2(new_n815), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n809), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G384));
  OAI211_X1 g0620(.A(G116), .B(new_n216), .C1(new_n531), .C2(KEYINPUT35), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(KEYINPUT35), .B2(new_n531), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT36), .ZN(new_n823));
  OR3_X1    g0623(.A1(new_n218), .A2(new_n319), .A3(new_n413), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n412), .A2(G50), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT96), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n208), .B(G13), .C1(new_n824), .C2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n390), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT97), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n650), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n366), .A2(new_n663), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n832), .B1(new_n399), .B2(new_n830), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n662), .B(new_n806), .C1(new_n635), .C2(new_n644), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n836), .B1(new_n837), .B2(new_n804), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT38), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n440), .A2(new_n453), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT37), .ZN(new_n841));
  INV_X1    g0641(.A(new_n660), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n429), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n840), .A2(KEYINPUT100), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n440), .A2(new_n843), .A3(new_n841), .A4(new_n453), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT100), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT99), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n448), .A2(new_n410), .A3(new_n417), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n424), .A2(KEYINPUT98), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n444), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n448), .A2(new_n410), .A3(new_n417), .A4(new_n850), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n443), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n848), .B1(new_n854), .B2(new_n660), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n851), .B1(new_n418), .B2(new_n423), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n856), .A2(new_n269), .A3(new_n853), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n405), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n858), .A2(new_n439), .B1(new_n450), .B2(new_n452), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(KEYINPUT99), .A3(new_n842), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n855), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n844), .A2(new_n847), .B1(new_n861), .B2(KEYINPUT37), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT99), .B1(new_n858), .B2(new_n842), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n848), .B(new_n660), .C1(new_n857), .C2(new_n405), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n442), .B2(new_n454), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n839), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n652), .A2(new_n648), .B1(new_n863), .B2(new_n864), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n845), .B(KEYINPUT100), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n841), .B1(new_n865), .B2(new_n859), .ZN(new_n870));
  OAI211_X1 g0670(.A(KEYINPUT38), .B(new_n868), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n838), .A2(new_n872), .B1(new_n442), .B2(new_n842), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n841), .B1(new_n840), .B2(new_n843), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n847), .B2(new_n844), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n843), .B1(new_n442), .B2(new_n454), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n839), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n877), .A2(new_n871), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT102), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT102), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n877), .A2(new_n871), .A3(new_n881), .A4(new_n878), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n867), .A2(new_n871), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT101), .B1(new_n883), .B2(KEYINPUT39), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT101), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n885), .B(new_n878), .C1(new_n867), .C2(new_n871), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n880), .B(new_n882), .C1(new_n884), .C2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n650), .A2(new_n662), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n873), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n455), .B1(new_n353), .B2(new_n354), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n689), .A2(KEYINPUT103), .A3(new_n356), .A4(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT103), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n684), .A2(KEYINPUT29), .A3(new_n663), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n811), .B2(new_n687), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n892), .B1(new_n457), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n891), .A2(new_n895), .A3(new_n655), .ZN(new_n896));
  XOR2_X1   g0696(.A(new_n889), .B(new_n896), .Z(new_n897));
  INV_X1    g0697(.A(KEYINPUT40), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n877), .B2(new_n871), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n831), .A2(new_n833), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n399), .A2(new_n830), .A3(new_n832), .ZN(new_n901));
  AND4_X1   g0701(.A1(new_n814), .A2(new_n900), .A3(new_n807), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n814), .A2(new_n900), .A3(new_n901), .A4(new_n807), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n872), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n903), .B(G330), .C1(new_n905), .C2(KEYINPUT40), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n355), .A2(new_n356), .A3(new_n456), .A4(new_n709), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n902), .A2(new_n883), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n909), .A2(new_n898), .B1(new_n902), .B2(new_n899), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(new_n458), .A3(new_n814), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n897), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n208), .B2(new_n712), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n897), .A2(new_n912), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n828), .B1(new_n914), .B2(new_n915), .ZN(G367));
  INV_X1    g0716(.A(new_n642), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n501), .A2(new_n662), .ZN(new_n918));
  MUX2_X1   g0718(.A(new_n499), .B(new_n917), .S(new_n918), .Z(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n724), .ZN(new_n920));
  OAI221_X1 g0720(.A(new_n726), .B1(new_n212), .B2(new_n323), .C1(new_n718), .C2(new_n236), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n921), .A2(new_n776), .ZN(new_n922));
  INV_X1    g0722(.A(new_n743), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n923), .A2(G294), .B1(new_n741), .B2(G283), .ZN(new_n924));
  INV_X1    g0724(.A(G317), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n924), .B1(new_n766), .B2(new_n731), .C1(new_n757), .C2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(G303), .B2(new_n752), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT46), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n736), .B2(new_n464), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT105), .Z(new_n930));
  OAI21_X1  g0730(.A(new_n247), .B1(new_n744), .B2(new_n478), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n736), .A2(new_n928), .A3(new_n464), .ZN(new_n932));
  INV_X1    g0732(.A(new_n733), .ZN(new_n933));
  AOI211_X1 g0733(.A(new_n931), .B(new_n932), .C1(G107), .C2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n927), .A2(new_n930), .A3(new_n934), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT106), .Z(new_n936));
  XOR2_X1   g0736(.A(KEYINPUT107), .B(G137), .Z(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n771), .A2(new_n938), .B1(G58), .B2(new_n737), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n940), .A2(KEYINPUT108), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(KEYINPUT108), .ZN(new_n942));
  OAI221_X1 g0742(.A(new_n253), .B1(new_n740), .B2(new_n202), .C1(new_n733), .C2(new_n412), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n923), .A2(new_n784), .B1(new_n761), .B2(G143), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n319), .B2(new_n744), .ZN(new_n945));
  AOI211_X1 g0745(.A(new_n943), .B(new_n945), .C1(G150), .C2(new_n752), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n941), .A2(new_n942), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n936), .A2(KEYINPUT47), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n725), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT47), .B1(new_n936), .B2(new_n947), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n920), .B(new_n922), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n713), .A2(G1), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n636), .B1(new_n538), .B2(new_n663), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n628), .A2(new_n662), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n674), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT44), .Z(new_n957));
  NOR2_X1   g0757(.A1(new_n674), .A2(new_n955), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT45), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(new_n671), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n667), .A2(KEYINPUT104), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n670), .A2(new_n672), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n673), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n962), .B(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n710), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n710), .B1(new_n961), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n677), .B(KEYINPUT41), .Z(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n952), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n955), .A2(new_n673), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT42), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n537), .B1(new_n953), .B2(new_n589), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n663), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n971), .A2(new_n972), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT43), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n976), .A2(new_n977), .B1(new_n978), .B2(new_n919), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n919), .A2(new_n978), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n671), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n982), .A2(new_n955), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n981), .B(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n951), .B1(new_n970), .B2(new_n984), .ZN(G387));
  AOI22_X1  g0785(.A1(new_n761), .A2(G322), .B1(new_n741), .B2(G303), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n766), .B2(new_n743), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G317), .B2(new_n752), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n988), .A2(KEYINPUT48), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(KEYINPUT48), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n933), .A2(G283), .B1(new_n737), .B2(G294), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT49), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n992), .A2(new_n993), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n247), .B1(new_n744), .B2(new_n464), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n771), .B2(G326), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n994), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n737), .A2(G77), .ZN(new_n999));
  INV_X1    g0799(.A(G159), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n999), .B1(new_n740), .B2(new_n412), .C1(new_n1000), .C2(new_n731), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n744), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n247), .B(new_n1001), .C1(G97), .C2(new_n1002), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n752), .A2(G50), .B1(new_n401), .B2(new_n923), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n771), .A2(G150), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n485), .A2(new_n933), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n728), .B1(new_n998), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n270), .A2(new_n202), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT50), .Z(new_n1010));
  INV_X1    g0810(.A(new_n679), .ZN(new_n1011));
  AOI211_X1 g0811(.A(G45), .B(new_n1011), .C1(G68), .C2(G77), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n718), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n233), .B2(new_n259), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n715), .A2(new_n1011), .B1(new_n528), .B2(new_n676), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n714), .B(new_n1008), .C1(new_n726), .C2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT109), .Z(new_n1018));
  NAND2_X1  g0818(.A1(new_n670), .A2(new_n724), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n1018), .A2(new_n1019), .B1(new_n965), .B2(new_n952), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n966), .A2(new_n677), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n710), .A2(new_n965), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(G393));
  NAND2_X1  g0823(.A1(new_n955), .A2(new_n724), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n751), .A2(new_n1000), .B1(new_n786), .B2(new_n731), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT51), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n253), .B1(new_n744), .B2(new_n433), .C1(new_n733), .C2(new_n319), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n923), .A2(G50), .B1(new_n741), .B2(new_n270), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n412), .B2(new_n736), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1027), .B(new_n1029), .C1(G143), .C2(new_n771), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n751), .A2(new_n766), .B1(new_n925), .B2(new_n731), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT52), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n247), .B1(new_n744), .B2(new_n528), .C1(new_n733), .C2(new_n464), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n923), .A2(G303), .B1(new_n741), .B2(G294), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n768), .B2(new_n736), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1033), .B(new_n1035), .C1(G322), .C2(new_n771), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n1026), .A2(new_n1030), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1037), .A2(KEYINPUT110), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n728), .B1(new_n1037), .B2(KEYINPUT110), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n726), .B1(new_n478), .B2(new_n212), .C1(new_n718), .C2(new_n243), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1024), .A2(new_n776), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n952), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n961), .A2(new_n966), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n677), .B1(new_n961), .B2(new_n966), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1042), .B1(new_n961), .B2(new_n1043), .C1(new_n1045), .C2(new_n1046), .ZN(G390));
  AOI21_X1  g0847(.A(new_n888), .B1(new_n877), .B2(new_n871), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n684), .A2(new_n663), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n804), .B1(new_n1049), .B2(new_n803), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n900), .A2(new_n901), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n836), .A2(new_n709), .A3(new_n807), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n812), .A2(new_n805), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n888), .B1(new_n1054), .B2(new_n836), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1052), .B(new_n1053), .C1(new_n887), .C2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT112), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n885), .B1(new_n872), .B2(new_n878), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n883), .A2(KEYINPUT101), .A3(KEYINPUT39), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n880), .A2(new_n882), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n888), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n838), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1065), .A2(KEYINPUT112), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1058), .A2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n836), .A2(KEYINPUT111), .A3(new_n709), .A4(new_n807), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT111), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n900), .A2(new_n901), .A3(new_n807), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1069), .B1(new_n1070), .B2(new_n815), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n1065), .B2(new_n1052), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1067), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1051), .B1(new_n815), .B2(new_n806), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1053), .A2(new_n1050), .A3(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n709), .A2(new_n807), .B1(new_n900), .B2(new_n901), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1054), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1077), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT113), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n907), .B(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n457), .A2(new_n894), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n654), .B1(new_n1084), .B2(KEYINPUT103), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1081), .A2(new_n1083), .A3(new_n1085), .A4(new_n895), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1075), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1086), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1067), .A2(new_n1074), .A3(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1087), .A2(new_n677), .A3(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1067), .A2(new_n952), .A3(new_n1074), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(KEYINPUT114), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1073), .B1(new_n1058), .B2(new_n1066), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT114), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n1094), .A3(new_n952), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n714), .B1(new_n400), .B2(new_n799), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n752), .A2(G132), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n771), .A2(G125), .ZN(new_n1099));
  INV_X1    g0899(.A(G128), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n253), .B1(new_n744), .B2(new_n202), .C1(new_n1100), .C2(new_n731), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n737), .A2(G150), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT53), .ZN(new_n1103));
  NOR4_X1   g0903(.A1(new_n1098), .A2(new_n1099), .A3(new_n1101), .A4(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT54), .B(G143), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n923), .A2(new_n938), .B1(new_n741), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n1000), .B2(new_n733), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT115), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n247), .B1(new_n736), .B2(new_n433), .C1(new_n733), .C2(new_n319), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n412), .A2(new_n744), .B1(new_n740), .B2(new_n478), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n731), .A2(new_n768), .B1(new_n743), .B2(new_n528), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G116), .A2(new_n752), .B1(new_n771), .B2(G294), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1104), .A2(new_n1109), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1097), .B1(new_n728), .B2(new_n1115), .C1(new_n887), .C2(new_n723), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1090), .A2(new_n1096), .A3(new_n1116), .ZN(G378));
  INV_X1    g0917(.A(KEYINPUT57), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n907), .B(KEYINPUT113), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n896), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1089), .A2(new_n1120), .ZN(new_n1121));
  XOR2_X1   g0921(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1122));
  NAND3_X1  g0922(.A1(new_n306), .A2(new_n310), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1122), .B1(new_n306), .B2(new_n310), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n289), .A2(new_n842), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT116), .Z(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n1124), .A2(new_n1125), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n306), .A2(new_n310), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1122), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1127), .B1(new_n1132), .B2(new_n1123), .ZN(new_n1133));
  OAI21_X1  g0933(.A(KEYINPUT117), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1128), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1132), .A2(new_n1127), .A3(new_n1123), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT117), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n910), .A2(new_n1134), .A3(G330), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n906), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n889), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1063), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1141), .B(new_n1139), .C1(new_n1144), .C2(new_n873), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1118), .B1(new_n1121), .B2(new_n1147), .ZN(new_n1148));
  AOI211_X1 g0948(.A(KEYINPUT57), .B(new_n1146), .C1(new_n1089), .C2(new_n1120), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n677), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n722), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n714), .B1(new_n202), .B2(new_n799), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G132), .A2(new_n923), .B1(new_n737), .B2(new_n1106), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n761), .A2(G125), .B1(new_n741), .B2(G137), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1156), .B1(new_n786), .B2(new_n733), .C1(new_n1100), .C2(new_n751), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n771), .A2(G124), .ZN(new_n1160));
  AOI211_X1 g0960(.A(G33), .B(G41), .C1(new_n784), .C2(new_n1002), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n752), .A2(G107), .B1(new_n485), .B2(new_n741), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n768), .B2(new_n757), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n253), .A2(G41), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n411), .B2(new_n744), .C1(new_n464), .C2(new_n731), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n999), .B1(new_n743), .B2(new_n478), .C1(new_n733), .C2(new_n412), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n1164), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1168), .A2(KEYINPUT58), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(KEYINPUT58), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1165), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1171), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1172));
  AND4_X1   g0972(.A1(new_n1162), .A2(new_n1169), .A3(new_n1170), .A4(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1152), .B(new_n1153), .C1(new_n728), .C2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n1146), .B2(new_n1043), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1150), .A2(new_n1176), .ZN(G375));
  NAND3_X1  g0977(.A1(new_n1083), .A2(new_n1085), .A3(new_n895), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1081), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1180), .A2(new_n969), .A3(new_n1086), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n714), .B1(new_n412), .B2(new_n799), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n761), .A2(G294), .B1(new_n741), .B2(G107), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(new_n478), .B2(new_n736), .C1(new_n464), .C2(new_n743), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n253), .B(new_n1184), .C1(G77), .C2(new_n1002), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1006), .B1(new_n593), .B2(new_n757), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G283), .B2(new_n752), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n757), .A2(new_n1100), .B1(new_n1000), .B2(new_n736), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT118), .Z(new_n1189));
  OAI221_X1 g0989(.A(new_n253), .B1(new_n744), .B2(new_n411), .C1(new_n733), .C2(new_n202), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G132), .A2(new_n761), .B1(new_n923), .B2(new_n1106), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n786), .B2(new_n740), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1190), .B(new_n1192), .C1(new_n752), .C2(new_n938), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1185), .A2(new_n1187), .B1(new_n1189), .B2(new_n1193), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1182), .B1(new_n728), .B2(new_n1194), .C1(new_n836), .C2(new_n723), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n1179), .B2(new_n1043), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1181), .A2(new_n1197), .ZN(G381));
  AND4_X1   g0998(.A1(new_n1094), .A2(new_n1067), .A3(new_n952), .A4(new_n1074), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1094), .B1(new_n1093), .B2(new_n952), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1116), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1089), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n677), .B1(new_n1093), .B2(new_n1088), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1201), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1150), .A2(new_n1205), .A3(new_n1176), .ZN(new_n1206));
  OR2_X1    g1006(.A1(G387), .A2(G390), .ZN(new_n1207));
  OR3_X1    g1007(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1208));
  OR4_X1    g1008(.A1(G381), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(G407));
  OAI211_X1 g1009(.A(G407), .B(G213), .C1(G343), .C2(new_n1206), .ZN(G409));
  NAND2_X1  g1010(.A1(new_n661), .A2(G213), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1146), .B1(new_n1089), .B2(new_n1120), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1118), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1178), .B1(new_n1093), .B2(new_n1088), .ZN(new_n1214));
  OAI21_X1  g1014(.A(KEYINPUT57), .B1(new_n1214), .B2(new_n1146), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n678), .B1(new_n1213), .B2(new_n1215), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1216), .A2(new_n1205), .A3(new_n1175), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1175), .B1(new_n1212), .B2(new_n969), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(G378), .A2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1211), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT121), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1086), .A2(new_n677), .ZN(new_n1222));
  OAI21_X1  g1022(.A(KEYINPUT60), .B1(new_n1120), .B2(new_n1081), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT60), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1178), .A2(new_n1179), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1222), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n1226), .A2(new_n819), .A3(new_n1196), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n678), .B1(new_n1120), .B2(new_n1081), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1120), .A2(KEYINPUT60), .A3(new_n1081), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1224), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1228), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(G384), .B1(new_n1231), .B2(new_n1197), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1221), .B1(new_n1227), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1211), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n819), .B1(new_n1226), .B2(new_n1196), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1231), .A2(G384), .A3(new_n1197), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n1236), .A3(KEYINPUT121), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1233), .A2(G2897), .A3(new_n1234), .A4(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1234), .A2(G2897), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1235), .A2(new_n1236), .A3(KEYINPUT121), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT121), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1239), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1238), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(KEYINPUT61), .B1(new_n1220), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1150), .A2(G378), .A3(new_n1176), .ZN(new_n1246));
  OR2_X1    g1046(.A1(G378), .A2(new_n1218), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1227), .A2(new_n1232), .ZN(new_n1249));
  AND4_X1   g1049(.A1(KEYINPUT62), .A2(new_n1248), .A3(new_n1211), .A4(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1234), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT62), .B1(new_n1251), .B2(new_n1249), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1245), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G387), .A2(G390), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1207), .A2(new_n1254), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(G393), .B(G396), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1207), .A2(new_n1256), .A3(new_n1254), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  XOR2_X1   g1060(.A(new_n1260), .B(KEYINPUT124), .Z(new_n1261));
  NAND2_X1  g1061(.A1(new_n1253), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT61), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1258), .A2(new_n1263), .A3(new_n1259), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1243), .B1(new_n1248), .B2(new_n1211), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT122), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1264), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(KEYINPUT122), .B1(new_n1251), .B2(new_n1243), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT120), .ZN(new_n1269));
  XOR2_X1   g1069(.A(KEYINPUT119), .B(KEYINPUT63), .Z(new_n1270));
  AOI211_X1 g1070(.A(new_n1269), .B(new_n1270), .C1(new_n1251), .C2(new_n1249), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1211), .B(new_n1249), .C1(new_n1217), .C2(new_n1219), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1270), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT120), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1267), .B(new_n1268), .C1(new_n1271), .C2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1251), .A2(KEYINPUT63), .A3(new_n1249), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT123), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1276), .B(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1262), .B1(new_n1275), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT125), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1262), .B(KEYINPUT125), .C1(new_n1275), .C2(new_n1278), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(G405));
  NAND2_X1  g1083(.A1(G375), .A2(G378), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1206), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1249), .A2(KEYINPUT126), .ZN(new_n1286));
  OR2_X1    g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(new_n1260), .A3(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1260), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1289), .B1(new_n1290), .B2(KEYINPUT127), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1291), .B1(KEYINPUT127), .B2(new_n1290), .ZN(G402));
endmodule


