//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1294, new_n1295, new_n1296;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  INV_X1    g0006(.A(G244), .ZN(new_n207));
  INV_X1    g0007(.A(G116), .ZN(new_n208));
  INV_X1    g0008(.A(G270), .ZN(new_n209));
  OAI22_X1  g0009(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n211), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n210), .B(new_n215), .C1(G68), .C2(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(KEYINPUT65), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n218), .A2(KEYINPUT65), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n202), .B2(new_n217), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT66), .Z(new_n224));
  INV_X1    g0024(.A(KEYINPUT1), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT67), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(KEYINPUT64), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g0030(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(G20), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(G50), .B1(G58), .B2(G68), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n222), .A2(G13), .ZN(new_n238));
  OAI211_X1 g0038(.A(new_n238), .B(G250), .C1(G257), .C2(G264), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n239), .B(KEYINPUT0), .Z(new_n240));
  AOI21_X1  g0040(.A(new_n240), .B1(new_n224), .B2(new_n225), .ZN(new_n241));
  NAND3_X1  g0041(.A1(new_n227), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT68), .ZN(G361));
  XNOR2_X1  g0043(.A(G238), .B(G244), .ZN(new_n244));
  INV_X1    g0044(.A(G232), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT2), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n217), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G250), .B(G257), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G264), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(new_n209), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G358));
  XNOR2_X1  g0052(.A(G87), .B(G97), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(G107), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(new_n208), .ZN(new_n255));
  XOR2_X1   g0055(.A(new_n255), .B(KEYINPUT70), .Z(new_n256));
  XNOR2_X1  g0056(.A(G68), .B(G77), .ZN(new_n257));
  INV_X1    g0057(.A(G58), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n259), .B(KEYINPUT69), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(new_n202), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n256), .B(new_n261), .ZN(G351));
  INV_X1    g0062(.A(KEYINPUT72), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n263), .B1(new_n232), .B2(new_n265), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n230), .A2(KEYINPUT72), .A3(new_n231), .A4(new_n264), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G232), .A3(G1698), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT75), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n276), .B1(new_n217), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G97), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n280), .B1(new_n274), .B2(new_n275), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n268), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G1), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(G41), .B2(G45), .ZN(new_n284));
  INV_X1    g0084(.A(G274), .ZN(new_n285));
  OR2_X1    g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G238), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n264), .A2(G1), .A3(G13), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n284), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n287), .B1(new_n290), .B2(KEYINPUT76), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(KEYINPUT76), .B2(new_n290), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n282), .A2(new_n286), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT13), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n293), .B(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  OR3_X1    g0096(.A1(new_n295), .A2(KEYINPUT14), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(G179), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT14), .B1(new_n295), .B2(new_n296), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n301));
  AND3_X1   g0101(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n302));
  AOI21_X1  g0102(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT73), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n232), .A2(KEYINPUT73), .A3(new_n301), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(G1), .B2(new_n233), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT12), .ZN(new_n312));
  INV_X1    g0112(.A(G13), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(G1), .ZN(new_n314));
  INV_X1    g0114(.A(G68), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(G20), .A3(new_n315), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n311), .A2(G68), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n312), .B2(new_n316), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(G20), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n233), .A2(G33), .ZN(new_n320));
  NOR2_X1   g0120(.A1(G20), .A2(G33), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  OAI221_X1 g0122(.A(new_n319), .B1(new_n320), .B2(new_n206), .C1(new_n322), .C2(new_n202), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n308), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT77), .B(KEYINPUT11), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n324), .B(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n318), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n300), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G200), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n295), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n295), .A2(G190), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(new_n327), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n273), .A2(G223), .A3(G1698), .ZN(new_n335));
  INV_X1    g0135(.A(G222), .ZN(new_n336));
  OAI221_X1 g0136(.A(new_n335), .B1(new_n206), .B2(new_n273), .C1(new_n278), .C2(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT71), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n268), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n290), .A2(G226), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n339), .A2(new_n286), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G200), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n283), .A2(G13), .A3(G20), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n202), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT8), .B(G58), .ZN(new_n346));
  INV_X1    g0146(.A(G150), .ZN(new_n347));
  OAI22_X1  g0147(.A1(new_n346), .A2(new_n320), .B1(new_n347), .B2(new_n322), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(G20), .B2(new_n203), .ZN(new_n349));
  OAI221_X1 g0149(.A(new_n345), .B1(new_n309), .B2(new_n349), .C1(new_n310), .C2(new_n202), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT9), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n339), .A2(G190), .A3(new_n286), .A4(new_n340), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n350), .A2(new_n351), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n342), .A2(new_n352), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT10), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n341), .A2(new_n296), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n350), .B1(new_n341), .B2(G179), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(KEYINPUT78), .A2(G33), .ZN(new_n362));
  NOR2_X1   g0162(.A1(KEYINPUT78), .A2(G33), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n362), .A2(new_n363), .A3(new_n269), .ZN(new_n364));
  NOR2_X1   g0164(.A1(KEYINPUT3), .A2(G33), .ZN(new_n365));
  OAI211_X1 g0165(.A(G223), .B(new_n277), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT80), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n270), .A2(new_n211), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT78), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n270), .ZN(new_n370));
  NAND2_X1  g0170(.A1(KEYINPUT78), .A2(G33), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(KEYINPUT3), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n277), .B1(new_n372), .B2(new_n271), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n368), .B1(new_n373), .B2(G226), .ZN(new_n374));
  AOI21_X1  g0174(.A(G1698), .B1(new_n372), .B2(new_n271), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT80), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(new_n376), .A3(G223), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n367), .A2(new_n374), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n268), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n286), .B1(new_n289), .B2(new_n245), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(G179), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n380), .B1(new_n378), .B2(new_n268), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n296), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n372), .A2(new_n271), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT79), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n372), .A2(KEYINPUT79), .A3(new_n271), .ZN(new_n388));
  NOR2_X1   g0188(.A1(KEYINPUT7), .A2(G20), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n372), .A2(new_n233), .A3(new_n271), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n315), .B1(new_n391), .B2(KEYINPUT7), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g0193(.A(G58), .B(G68), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(G20), .B1(G159), .B2(new_n321), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(KEYINPUT16), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT16), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n269), .B1(new_n362), .B2(new_n363), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n398), .A2(KEYINPUT7), .A3(new_n233), .A4(new_n272), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT7), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(new_n273), .B2(G20), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n315), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n395), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n397), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n396), .A2(new_n404), .A3(new_n308), .ZN(new_n405));
  INV_X1    g0205(.A(new_n346), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(new_n344), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(new_n310), .B2(new_n406), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n384), .A2(new_n410), .A3(KEYINPUT18), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT18), .B1(new_n384), .B2(new_n410), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT82), .ZN(new_n414));
  INV_X1    g0214(.A(G190), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n379), .A2(new_n415), .A3(new_n381), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(G200), .B2(new_n383), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n403), .B1(new_n390), .B2(new_n392), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n309), .B1(new_n418), .B2(KEYINPUT16), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n408), .B1(new_n419), .B2(new_n404), .ZN(new_n420));
  XOR2_X1   g0220(.A(KEYINPUT81), .B(KEYINPUT17), .Z(new_n421));
  AND3_X1   g0221(.A1(new_n417), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(KEYINPUT81), .A2(KEYINPUT17), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n417), .B2(new_n420), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n414), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(G200), .B1(new_n379), .B2(new_n381), .ZN(new_n427));
  AOI211_X1 g0227(.A(G190), .B(new_n380), .C1(new_n378), .C2(new_n268), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n423), .B1(new_n429), .B2(new_n410), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n417), .A2(new_n420), .A3(new_n421), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(KEYINPUT82), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n413), .B1(new_n426), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n344), .A2(new_n206), .ZN(new_n434));
  XNOR2_X1  g0234(.A(KEYINPUT15), .B(G87), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(new_n320), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n346), .A2(new_n322), .B1(new_n233), .B2(new_n206), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n308), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n434), .B(new_n438), .C1(new_n310), .C2(new_n206), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n286), .B1(new_n289), .B2(new_n207), .ZN(new_n440));
  XOR2_X1   g0240(.A(new_n440), .B(KEYINPUT74), .Z(new_n441));
  NAND2_X1  g0241(.A1(G238), .A2(G1698), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n273), .B(new_n442), .C1(new_n245), .C2(G1698), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n268), .B(new_n443), .C1(G107), .C2(new_n273), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n439), .B1(G200), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n415), .B2(new_n445), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n433), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(new_n296), .ZN(new_n449));
  INV_X1    g0249(.A(G179), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n441), .A2(new_n444), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n439), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g0253(.A1(new_n334), .A2(new_n361), .A3(new_n448), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n283), .A2(G33), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n306), .A2(new_n307), .A3(new_n343), .A4(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(new_n213), .ZN(new_n457));
  AND2_X1   g0257(.A1(KEYINPUT83), .A2(G97), .ZN(new_n458));
  NOR2_X1   g0258(.A1(KEYINPUT83), .A2(G97), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G107), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(KEYINPUT6), .A3(new_n461), .ZN(new_n462));
  XOR2_X1   g0262(.A(G97), .B(G107), .Z(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(KEYINPUT6), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G20), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n399), .A2(new_n401), .ZN(new_n466));
  OAI221_X1 g0266(.A(new_n465), .B1(new_n206), .B2(new_n322), .C1(new_n466), .C2(new_n461), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n457), .B1(new_n467), .B2(new_n308), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n343), .A2(G97), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT85), .ZN(new_n471));
  INV_X1    g0271(.A(new_n288), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT5), .B(G41), .ZN(new_n473));
  INV_X1    g0273(.A(G45), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(G1), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n472), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n473), .A2(new_n475), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n476), .A2(G257), .B1(new_n478), .B2(G274), .ZN(new_n479));
  AND2_X1   g0279(.A1(KEYINPUT4), .A2(G244), .ZN(new_n480));
  AND2_X1   g0280(.A1(KEYINPUT3), .A2(G33), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n277), .B(new_n480), .C1(new_n481), .C2(new_n365), .ZN(new_n482));
  OAI211_X1 g0282(.A(G250), .B(G1698), .C1(new_n481), .C2(new_n365), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G283), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(G244), .B(new_n277), .C1(new_n364), .C2(new_n365), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT4), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n266), .A2(new_n267), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n479), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n471), .B1(new_n490), .B2(G179), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT4), .B1(new_n375), .B2(G244), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n268), .B1(new_n492), .B2(new_n485), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n493), .A2(KEYINPUT85), .A3(new_n450), .A4(new_n479), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n468), .A2(new_n470), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT84), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n479), .B(new_n496), .C1(new_n488), .C2(new_n489), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n496), .B1(new_n493), .B2(new_n479), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n296), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n490), .A2(KEYINPUT84), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n497), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G190), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n490), .A2(G200), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n505), .A2(new_n470), .A3(new_n468), .A4(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n208), .A2(G20), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n509), .A2(G1), .A3(new_n313), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n232), .A2(new_n301), .B1(G20), .B2(new_n208), .ZN(new_n512));
  XNOR2_X1  g0312(.A(KEYINPUT83), .B(G97), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n233), .B(new_n484), .C1(new_n513), .C2(G33), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n512), .A2(KEYINPUT20), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT20), .B1(new_n512), .B2(new_n514), .ZN(new_n516));
  OAI221_X1 g0316(.A(new_n511), .B1(new_n456), .B2(new_n208), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(G264), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G1698), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n214), .A2(new_n277), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n385), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n273), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G303), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n521), .A2(new_n523), .B1(new_n266), .B2(new_n267), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n478), .A2(G274), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n477), .A2(new_n288), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n527), .A2(new_n209), .ZN(new_n528));
  NOR3_X1   g0328(.A1(new_n524), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n517), .A2(new_n529), .A3(G179), .ZN(new_n530));
  OAI22_X1  g0330(.A1(new_n515), .A2(new_n516), .B1(new_n456), .B2(new_n208), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(new_n510), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n476), .A2(G270), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n372), .A2(new_n271), .B1(new_n214), .B2(new_n277), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n534), .A2(new_n519), .B1(G303), .B2(new_n522), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n525), .B(new_n533), .C1(new_n535), .C2(new_n489), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G169), .ZN(new_n537));
  OAI21_X1  g0337(.A(KEYINPUT21), .B1(new_n532), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n521), .A2(new_n523), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n528), .B1(new_n539), .B2(new_n268), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n296), .B1(new_n540), .B2(new_n525), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT21), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n542), .A3(new_n517), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n530), .B1(new_n538), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n536), .A2(G200), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n415), .B2(new_n536), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n544), .B1(new_n517), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n214), .A2(G1698), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n212), .A2(new_n277), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n385), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n362), .A2(new_n363), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G294), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n268), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n476), .A2(G264), .B1(new_n478), .B2(G274), .ZN(new_n556));
  AOI21_X1  g0356(.A(G200), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n525), .B1(new_n518), .B2(new_n527), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT87), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n372), .A2(new_n271), .B1(new_n212), .B2(new_n277), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n560), .A2(new_n549), .B1(G294), .B2(new_n552), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n559), .B1(new_n561), .B2(new_n489), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n554), .A2(KEYINPUT87), .A3(new_n268), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n558), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n557), .B1(new_n564), .B2(new_n415), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n211), .A2(G20), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n385), .A2(KEYINPUT22), .A3(new_n566), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n362), .A2(new_n363), .A3(new_n208), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n566), .B1(new_n481), .B2(new_n365), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT22), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n233), .A2(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n233), .A2(G107), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n572), .B(KEYINPUT23), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n567), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT24), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n567), .A2(new_n571), .A3(KEYINPUT24), .A4(new_n573), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(new_n308), .A3(new_n577), .ZN(new_n578));
  OR2_X1    g0378(.A1(new_n456), .A2(new_n461), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n314), .A2(new_n572), .ZN(new_n580));
  XOR2_X1   g0380(.A(new_n580), .B(KEYINPUT25), .Z(new_n581));
  NAND3_X1  g0381(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  OR2_X1    g0382(.A1(new_n565), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n555), .A2(G179), .A3(new_n556), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n564), .B2(new_n296), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n582), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g0387(.A(KEYINPUT86), .B(G87), .Z(new_n588));
  NAND3_X1  g0388(.A1(new_n588), .A2(new_n461), .A3(new_n513), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT19), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n233), .B1(new_n280), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n385), .A2(new_n233), .A3(G68), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n590), .B1(new_n513), .B2(new_n320), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n595), .A2(new_n308), .B1(new_n344), .B2(new_n435), .ZN(new_n596));
  OR2_X1    g0396(.A1(new_n456), .A2(new_n435), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n475), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(G250), .A3(new_n288), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n285), .B2(new_n599), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n372), .A2(new_n271), .B1(new_n207), .B2(G1698), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n287), .A2(new_n277), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n568), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n601), .B1(new_n606), .B2(new_n268), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n450), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n598), .B(new_n608), .C1(G169), .C2(new_n607), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(G190), .ZN(new_n610));
  INV_X1    g0410(.A(new_n601), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n568), .B1(new_n602), .B2(new_n603), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n611), .B1(new_n612), .B2(new_n489), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(G200), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n456), .A2(new_n211), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n610), .A2(new_n596), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n609), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n587), .A2(new_n617), .ZN(new_n618));
  AND4_X1   g0418(.A1(new_n454), .A2(new_n508), .A3(new_n548), .A4(new_n618), .ZN(G372));
  INV_X1    g0419(.A(new_n360), .ZN(new_n620));
  INV_X1    g0420(.A(new_n333), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n329), .B2(new_n452), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n422), .A2(new_n425), .A3(new_n414), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT82), .B1(new_n430), .B2(new_n431), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n411), .A2(new_n412), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n620), .B1(new_n627), .B2(new_n356), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n495), .A2(new_n501), .A3(new_n609), .A4(new_n616), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n598), .A2(new_n608), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n606), .A2(KEYINPUT88), .A3(new_n268), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT88), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n612), .B2(new_n489), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n631), .A2(new_n633), .A3(new_n611), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n296), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT89), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT89), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n630), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n629), .A2(KEYINPUT26), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n502), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n565), .A2(new_n582), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n544), .B2(new_n586), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n641), .B1(new_n643), .B2(new_n507), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n634), .A2(G200), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n645), .A2(new_n596), .A3(new_n610), .A4(new_n615), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n636), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n640), .B1(new_n644), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n454), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n628), .A2(new_n650), .ZN(G369));
  NAND2_X1  g0451(.A1(new_n314), .A2(new_n233), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT90), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n653), .A2(KEYINPUT90), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n654), .A2(G213), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n517), .ZN(new_n660));
  XOR2_X1   g0460(.A(new_n660), .B(KEYINPUT91), .Z(new_n661));
  NOR2_X1   g0461(.A1(new_n548), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n661), .A2(new_n544), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n665));
  INV_X1    g0465(.A(new_n659), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n583), .B(new_n586), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n584), .ZN(new_n668));
  AOI221_X4 g0468(.A(new_n559), .B1(new_n266), .B2(new_n267), .C1(new_n551), .C2(new_n553), .ZN(new_n669));
  AOI21_X1  g0469(.A(KEYINPUT87), .B1(new_n554), .B2(new_n268), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n556), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n668), .B1(new_n671), .B2(G169), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(new_n665), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n659), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n664), .A2(G330), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n643), .A2(new_n666), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(G399));
  OR2_X1    g0478(.A1(new_n589), .A2(G116), .ZN(new_n679));
  INV_X1    g0479(.A(new_n238), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G41), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G1), .ZN(new_n683));
  OAI22_X1  g0483(.A1(new_n679), .A2(new_n683), .B1(new_n235), .B2(new_n682), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT29), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n649), .A2(new_n686), .A3(new_n666), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n636), .A2(new_n646), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT95), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n502), .A2(new_n507), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n690), .B1(new_n502), .B2(new_n507), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n643), .B(new_n689), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n689), .A2(new_n641), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n694), .A2(KEYINPUT26), .B1(new_n637), .B2(new_n639), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n693), .B(new_n695), .C1(KEYINPUT26), .C2(new_n629), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n686), .B1(new_n696), .B2(new_n666), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT92), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n558), .B1(new_n268), .B2(new_n554), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n699), .A2(new_n607), .A3(G179), .A4(new_n540), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n698), .B1(new_n500), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n613), .A2(new_n524), .A3(new_n528), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n504), .A2(KEYINPUT92), .A3(new_n668), .A4(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT93), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n500), .A2(new_n702), .A3(new_n700), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n699), .A2(G179), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n709), .A2(new_n490), .A3(new_n634), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n708), .B1(new_n536), .B2(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n701), .A2(KEYINPUT93), .A3(new_n704), .A4(new_n702), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n707), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n659), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT94), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n711), .A2(new_n705), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT31), .B1(new_n713), .B2(new_n659), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT94), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n618), .A2(new_n508), .A3(new_n548), .A4(new_n666), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n718), .A2(new_n720), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  AOI211_X1 g0524(.A(new_n688), .B(new_n697), .C1(new_n724), .C2(G330), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n685), .B1(new_n725), .B2(G1), .ZN(G364));
  NAND2_X1  g0526(.A1(new_n664), .A2(G330), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n313), .A2(G20), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n283), .B1(new_n728), .B2(G45), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n681), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(G330), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(new_n662), .B2(new_n663), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n727), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n387), .A2(new_n388), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n680), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n236), .A2(new_n474), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n737), .B(new_n738), .C1(new_n261), .C2(new_n474), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n273), .A2(G355), .A3(new_n238), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n739), .B(new_n740), .C1(G116), .C2(new_n238), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n232), .B1(G20), .B2(new_n296), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G303), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n415), .A2(new_n330), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(G20), .A3(new_n450), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n233), .A2(new_n450), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(new_n415), .A3(new_n330), .ZN(new_n751));
  INV_X1    g0551(.A(G311), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n747), .A2(new_n749), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n415), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n756), .A2(G322), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n233), .A2(G190), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n758), .A2(G179), .A3(G200), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(KEYINPUT33), .B(G317), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n753), .B(new_n757), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n233), .B1(new_n754), .B2(new_n450), .ZN(new_n763));
  INV_X1    g0563(.A(G294), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n758), .A2(new_n450), .A3(G200), .ZN(new_n766));
  INV_X1    g0566(.A(G283), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n522), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n758), .A2(new_n450), .A3(new_n330), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n765), .B(new_n768), .C1(G329), .C2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G326), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n748), .A2(G20), .A3(G179), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n762), .B(new_n771), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n763), .A2(KEYINPUT98), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n763), .A2(KEYINPUT98), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G97), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n751), .B(KEYINPUT96), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G77), .ZN(new_n781));
  XNOR2_X1  g0581(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n770), .A2(G159), .A3(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n782), .ZN(new_n784));
  INV_X1    g0584(.A(G159), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n769), .B2(new_n785), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n779), .A2(new_n781), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n773), .A2(new_n202), .B1(new_n755), .B2(new_n258), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(G68), .B2(new_n760), .ZN(new_n789));
  INV_X1    g0589(.A(new_n766), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G107), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n749), .A2(new_n588), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n789), .A2(new_n273), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n774), .B1(new_n787), .B2(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n741), .A2(new_n746), .B1(new_n742), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n745), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n731), .B(new_n795), .C1(new_n664), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n735), .A2(new_n797), .ZN(G396));
  NAND2_X1  g0598(.A1(new_n724), .A2(G330), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n439), .A2(new_n659), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n453), .B1(new_n447), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n452), .A2(new_n659), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(new_n649), .B2(new_n666), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n517), .A2(new_n529), .A3(G179), .ZN(new_n805));
  AND4_X1   g0605(.A1(new_n542), .A2(new_n517), .A3(G169), .A4(new_n536), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n542), .B1(new_n541), .B2(new_n517), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n507), .B(new_n583), .C1(new_n808), .C2(new_n673), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n648), .B1(new_n809), .B2(new_n502), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n637), .A2(new_n639), .ZN(new_n811));
  INV_X1    g0611(.A(new_n629), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n812), .B2(new_n647), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n666), .B(new_n803), .C1(new_n810), .C2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT99), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n649), .A2(KEYINPUT99), .A3(new_n666), .A4(new_n803), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n804), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n799), .B(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n732), .ZN(new_n820));
  INV_X1    g0620(.A(new_n773), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G137), .A2(new_n821), .B1(new_n760), .B2(G150), .ZN(new_n822));
  INV_X1    g0622(.A(new_n780), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n823), .B2(new_n785), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G143), .B2(new_n756), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT34), .Z(new_n826));
  OAI22_X1  g0626(.A1(new_n749), .A2(new_n202), .B1(new_n766), .B2(new_n315), .ZN(new_n827));
  INV_X1    g0627(.A(new_n736), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n827), .B(new_n828), .C1(G132), .C2(new_n770), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n826), .B(new_n829), .C1(new_n258), .C2(new_n763), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n755), .A2(new_n764), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n790), .A2(G87), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n752), .B2(new_n769), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n273), .B(new_n833), .C1(G283), .C2(new_n760), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n749), .A2(new_n461), .B1(new_n773), .B2(new_n747), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(new_n780), .B2(G116), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n834), .A2(new_n779), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n830), .B1(new_n831), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n742), .A2(new_n743), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n838), .A2(new_n742), .B1(new_n206), .B2(new_n839), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n840), .B(new_n731), .C1(new_n744), .C2(new_n803), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n820), .A2(new_n841), .ZN(G384));
  AOI21_X1  g0642(.A(new_n208), .B1(new_n464), .B2(KEYINPUT35), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n843), .B(new_n234), .C1(KEYINPUT35), .C2(new_n464), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT36), .ZN(new_n845));
  OAI21_X1  g0645(.A(G77), .B1(new_n258), .B2(new_n315), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n846), .A2(new_n235), .B1(G50), .B2(new_n315), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n847), .A2(G1), .A3(new_n313), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n329), .B(new_n333), .C1(new_n327), .C2(new_n666), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n328), .B(new_n659), .C1(new_n621), .C2(new_n300), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AND3_X1   g0651(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n852), .A2(new_n721), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT102), .B1(new_n853), .B2(new_n723), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n716), .A2(KEYINPUT102), .A3(new_n723), .A4(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n803), .B(new_n851), .C1(new_n854), .C2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT38), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n417), .A2(new_n420), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n384), .A2(new_n410), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n860), .B(new_n861), .C1(new_n420), .C2(new_n657), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(KEYINPUT37), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n419), .B1(KEYINPUT16), .B2(new_n418), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n409), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n384), .ZN(new_n866));
  INV_X1    g0666(.A(new_n657), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n866), .A2(new_n868), .A3(new_n860), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n863), .B1(KEYINPUT37), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT100), .B1(new_n433), .B2(new_n868), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n626), .B1(new_n623), .B2(new_n624), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT100), .ZN(new_n873));
  INV_X1    g0673(.A(new_n868), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n859), .B(new_n870), .C1(new_n871), .C2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n626), .A2(new_n430), .A3(new_n431), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(new_n410), .A3(new_n867), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n862), .B(KEYINPUT37), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT38), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT40), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n858), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT101), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n871), .A2(new_n875), .ZN(new_n884));
  INV_X1    g0684(.A(new_n870), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT38), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n883), .B1(new_n886), .B2(new_n876), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n873), .B1(new_n872), .B2(new_n874), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n433), .A2(KEYINPUT100), .A3(new_n868), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n885), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n859), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n884), .A2(KEYINPUT38), .A3(new_n885), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(KEYINPUT101), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n803), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n716), .A2(new_n723), .A3(new_n855), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT102), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n894), .B1(new_n897), .B2(new_n856), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n887), .A2(new_n893), .A3(new_n851), .A4(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT40), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n882), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n897), .A2(new_n856), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n902), .A2(new_n454), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n901), .B(new_n903), .Z(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(G330), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT39), .B1(new_n886), .B2(new_n876), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  INV_X1    g0707(.A(new_n880), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n892), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n300), .A2(new_n328), .A3(new_n666), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n413), .A2(new_n657), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n802), .B1(new_n816), .B2(new_n817), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n887), .A2(new_n893), .A3(new_n851), .A4(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n913), .A2(new_n914), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n454), .B1(new_n697), .B2(new_n688), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n628), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n918), .B(new_n920), .ZN(new_n921));
  OAI22_X1  g0721(.A1(new_n905), .A2(new_n921), .B1(new_n283), .B2(new_n728), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT103), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n905), .A2(new_n921), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n845), .B(new_n848), .C1(new_n923), .C2(new_n924), .ZN(G367));
  NAND2_X1  g0725(.A1(new_n596), .A2(new_n615), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n659), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n689), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n811), .B2(new_n927), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n691), .A2(new_n692), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n468), .A2(new_n470), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n659), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n667), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n544), .A2(new_n659), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n939), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n935), .A2(new_n936), .A3(new_n937), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n935), .A2(new_n673), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n659), .B1(new_n944), .B2(new_n502), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n930), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(KEYINPUT104), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT104), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n949), .B(new_n930), .C1(new_n943), .C2(new_n945), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n947), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n948), .B1(new_n947), .B2(new_n950), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT106), .ZN(new_n953));
  INV_X1    g0753(.A(new_n676), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n934), .B1(new_n502), .B2(new_n666), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n951), .A2(new_n952), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n953), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n681), .B(KEYINPUT41), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n955), .A2(new_n677), .ZN(new_n963));
  XNOR2_X1  g0763(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n964), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT108), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT44), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n931), .A2(new_n677), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n965), .A2(new_n966), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n954), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n965), .A2(new_n676), .A3(new_n966), .A4(new_n971), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n937), .A2(new_n587), .ZN(new_n976));
  INV_X1    g0776(.A(new_n675), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n976), .B1(new_n977), .B2(new_n937), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n727), .B(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n725), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT109), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n725), .A2(KEYINPUT109), .A3(new_n979), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n975), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n962), .B1(new_n984), .B2(new_n725), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n959), .B(new_n960), .C1(new_n730), .C2(new_n985), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n828), .B1(new_n461), .B2(new_n763), .C1(new_n513), .C2(new_n766), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n773), .A2(new_n752), .B1(new_n755), .B2(new_n747), .ZN(new_n988));
  INV_X1    g0788(.A(new_n749), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(G116), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT46), .Z(new_n991));
  AOI211_X1 g0791(.A(new_n988), .B(new_n991), .C1(G283), .C2(new_n780), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n764), .B2(new_n759), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n987), .B(new_n993), .C1(G317), .C2(new_n770), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT110), .Z(new_n995));
  NOR2_X1   g0795(.A1(new_n755), .A2(new_n347), .ZN(new_n996));
  INV_X1    g0796(.A(G137), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n206), .A2(new_n766), .B1(new_n769), .B2(new_n997), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n522), .B(new_n998), .C1(G143), .C2(new_n821), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n778), .A2(G68), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n749), .A2(new_n258), .B1(new_n759), .B2(new_n785), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n780), .B2(G50), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n995), .B1(new_n996), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT47), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n732), .B1(new_n1005), .B2(new_n742), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n737), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n746), .B1(new_n238), .B2(new_n435), .C1(new_n1007), .C2(new_n251), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1006), .B(new_n1008), .C1(new_n796), .C2(new_n929), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n986), .A2(new_n1009), .ZN(G387));
  NAND2_X1  g0810(.A1(new_n982), .A2(new_n983), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n681), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT115), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n725), .A2(new_n979), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G322), .A2(new_n821), .B1(new_n760), .B2(G311), .ZN(new_n1016));
  INV_X1    g0816(.A(G317), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1016), .B1(new_n1017), .B2(new_n755), .C1(new_n823), .C2(new_n747), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT48), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n1018), .A2(new_n1019), .B1(new_n764), .B2(new_n749), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n763), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1020), .B1(G283), .B2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT113), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT49), .Z(new_n1026));
  OAI221_X1 g0826(.A(new_n828), .B1(new_n208), .B2(new_n766), .C1(new_n772), .C2(new_n769), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT114), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n773), .A2(new_n785), .B1(new_n769), .B2(new_n347), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n989), .A2(G77), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n202), .B2(new_n755), .C1(new_n315), .C2(new_n751), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1030), .B(new_n1032), .C1(G97), .C2(new_n790), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n777), .A2(new_n435), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n736), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n406), .B2(new_n760), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n742), .B1(new_n1029), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n977), .A2(new_n745), .ZN(new_n1038));
  XOR2_X1   g0838(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n346), .B2(G50), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n406), .A2(new_n1039), .A3(new_n202), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1041), .A2(new_n474), .A3(new_n1042), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n679), .B(new_n1043), .C1(G68), .C2(G77), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n737), .B1(new_n248), .B2(new_n474), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n679), .A2(new_n238), .A3(new_n273), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n238), .A2(G107), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n746), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AND3_X1   g0849(.A1(new_n1037), .A2(new_n1038), .A3(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1014), .A2(new_n1015), .B1(new_n731), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n979), .A2(new_n730), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT111), .Z(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1053), .ZN(G393));
  NAND3_X1  g0854(.A1(new_n973), .A2(new_n730), .A3(new_n974), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n746), .B1(new_n238), .B2(new_n513), .C1(new_n1007), .C2(new_n255), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n522), .B1(new_n759), .B2(new_n747), .C1(new_n767), .C2(new_n749), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n751), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1057), .B1(G294), .B2(new_n1058), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n773), .A2(new_n1017), .B1(new_n755), .B2(new_n752), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT52), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n770), .A2(G322), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G116), .A2(new_n1021), .B1(new_n790), .B2(G107), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n832), .B1(new_n315), .B2(new_n749), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G143), .B2(new_n770), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1066), .B(new_n736), .C1(new_n202), .C2(new_n759), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n778), .A2(G77), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n773), .A2(new_n347), .B1(new_n755), .B2(new_n785), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT51), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1068), .B(new_n1070), .C1(new_n346), .C2(new_n823), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1064), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n732), .B1(new_n1072), .B2(new_n742), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1056), .B(new_n1073), .C1(new_n955), .C2(new_n796), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1055), .A2(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT116), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n973), .A2(new_n974), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n682), .B1(new_n1011), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n984), .ZN(new_n1079));
  AOI21_X1  g0879(.A(KEYINPUT117), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1076), .A2(KEYINPUT117), .A3(new_n1079), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(G390));
  INV_X1    g0883(.A(new_n851), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n911), .B1(new_n915), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n906), .A2(new_n1085), .A3(new_n909), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n892), .A2(new_n908), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n696), .A2(new_n666), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n801), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n802), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1087), .B(new_n911), .C1(new_n1090), .C2(new_n1084), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n724), .A2(new_n851), .A3(G330), .A4(new_n803), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n1086), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n858), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1086), .A2(new_n1091), .B1(new_n1095), .B2(G330), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n902), .A2(G330), .A3(new_n454), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1098), .A2(new_n628), .A3(new_n919), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n851), .B1(new_n898), .B2(G330), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1092), .A2(new_n1090), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n902), .A2(G330), .A3(new_n803), .A4(new_n851), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n724), .A2(G330), .A3(new_n803), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n1084), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n915), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1100), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(KEYINPUT118), .B1(new_n1097), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1086), .A2(new_n1091), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n1104), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1086), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n916), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n733), .B(new_n894), .C1(new_n897), .C2(new_n856), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1090), .B(new_n1092), .C1(new_n1116), .C2(new_n851), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1099), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1113), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1109), .A2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1121), .B(new_n681), .C1(new_n1113), .C2(new_n1118), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1113), .A2(new_n730), .ZN(new_n1123));
  INV_X1    g0923(.A(G125), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n769), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n989), .A2(G150), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT53), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1125), .B(new_n1127), .C1(G50), .C2(new_n790), .ZN(new_n1128));
  INV_X1    g0928(.A(G132), .ZN(new_n1129));
  INV_X1    g0929(.A(G128), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n273), .B1(new_n755), .B2(new_n1129), .C1(new_n1130), .C2(new_n773), .ZN(new_n1131));
  XOR2_X1   g0931(.A(KEYINPUT54), .B(G143), .Z(new_n1132));
  AOI21_X1  g0932(.A(new_n1131), .B1(new_n780), .B2(new_n1132), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1128), .B(new_n1133), .C1(new_n785), .C2(new_n777), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G137), .B2(new_n760), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n315), .A2(new_n766), .B1(new_n769), .B2(new_n764), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n273), .B(new_n1136), .C1(G107), .C2(new_n760), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n749), .A2(new_n211), .B1(new_n755), .B2(new_n208), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n780), .B2(new_n460), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(new_n1068), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(G283), .B2(new_n821), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n742), .B1(new_n1135), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n839), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n731), .B1(new_n1143), .B2(new_n406), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT119), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1142), .B(new_n1145), .C1(new_n910), .C2(new_n744), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1122), .A2(new_n1123), .A3(new_n1146), .ZN(G378));
  INV_X1    g0947(.A(new_n918), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n899), .A2(new_n900), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n361), .B1(new_n350), .B2(new_n867), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n350), .A2(new_n867), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n356), .B2(new_n360), .ZN(new_n1152));
  OR3_X1    g0952(.A1(new_n1150), .A2(KEYINPUT55), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(KEYINPUT55), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1153), .A2(KEYINPUT56), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT56), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n882), .ZN(new_n1158));
  AND4_X1   g0958(.A1(G330), .A2(new_n1149), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1157), .B1(new_n901), .B2(G330), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1148), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1149), .A2(G330), .A3(new_n1158), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1157), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n901), .A2(G330), .A3(new_n1157), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1164), .A2(new_n918), .A3(new_n1165), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1121), .A2(new_n1100), .B1(new_n1161), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n681), .B1(new_n1167), .B2(KEYINPUT57), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1161), .A2(KEYINPUT120), .A3(new_n1166), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1097), .A2(new_n1108), .A3(KEYINPUT118), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1119), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1100), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT120), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1173), .B(new_n1148), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1174));
  AND4_X1   g0974(.A1(KEYINPUT57), .A2(new_n1169), .A3(new_n1172), .A4(new_n1174), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1168), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1157), .A2(new_n743), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n839), .A2(new_n202), .ZN(new_n1178));
  INV_X1    g0978(.A(G41), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n770), .A2(G283), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1000), .A2(new_n1179), .A3(new_n1031), .A4(new_n1180), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n821), .A2(G116), .B1(new_n756), .B2(G107), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1182), .B1(new_n213), .B2(new_n759), .C1(new_n435), .C2(new_n751), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n766), .A2(new_n258), .ZN(new_n1184));
  NOR4_X1   g0984(.A1(new_n1181), .A2(new_n1183), .A3(new_n736), .A4(new_n1184), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT58), .Z(new_n1186));
  OAI22_X1  g0986(.A1(new_n1124), .A2(new_n773), .B1(new_n751), .B2(new_n997), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n1129), .A2(new_n759), .B1(new_n755), .B2(new_n1130), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1187), .B(new_n1188), .C1(new_n778), .C2(G150), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1132), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1189), .B1(new_n749), .B2(new_n1190), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1193));
  AOI21_X1  g0993(.A(G33), .B1(new_n790), .B2(G159), .ZN(new_n1194));
  AOI21_X1  g0994(.A(G41), .B1(new_n770), .B2(G124), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G41), .B1(new_n736), .B2(G33), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1186), .B(new_n1196), .C1(G50), .C2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n732), .B1(new_n1198), .B2(new_n742), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1177), .A2(new_n1178), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1161), .A2(new_n1166), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1201), .B1(new_n1202), .B2(new_n730), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1176), .A2(new_n1203), .ZN(G375));
  AOI21_X1  g1004(.A(new_n729), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n206), .A2(new_n766), .B1(new_n769), .B2(new_n747), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n273), .B(new_n1206), .C1(G294), .C2(new_n821), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n989), .A2(G97), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n208), .A2(new_n759), .B1(new_n755), .B2(new_n767), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n780), .B2(G107), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1207), .A2(new_n1034), .A3(new_n1208), .A4(new_n1210), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n778), .A2(G50), .B1(G150), .B2(new_n1058), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1213), .A2(KEYINPUT121), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(KEYINPUT121), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G159), .A2(new_n989), .B1(new_n760), .B2(new_n1132), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n997), .B2(new_n755), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1184), .B(new_n1217), .C1(G128), .C2(new_n770), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1214), .A2(new_n736), .A3(new_n1215), .A4(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n773), .A2(new_n1129), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1211), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n742), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(G68), .B2(new_n1143), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n1084), .B2(new_n743), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1205), .B1(new_n731), .B2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1115), .A2(new_n1099), .A3(new_n1117), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1108), .A2(new_n1226), .A3(new_n961), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1227), .ZN(G381));
  INV_X1    g1028(.A(G375), .ZN(new_n1229));
  INV_X1    g1029(.A(G378), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1081), .A2(new_n986), .A3(new_n1009), .A4(new_n1082), .ZN(new_n1231));
  INV_X1    g1031(.A(G396), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1051), .A2(new_n1232), .A3(new_n1053), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(G381), .A2(G384), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1229), .A2(new_n1230), .A3(new_n1234), .A4(new_n1235), .ZN(G407));
  NAND3_X1  g1036(.A1(new_n1229), .A2(new_n658), .A3(new_n1230), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(G407), .A2(G213), .A3(new_n1237), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1238), .B(KEYINPUT122), .Z(G409));
  NAND2_X1  g1039(.A1(G390), .A2(G387), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1231), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1232), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1241), .A2(new_n1233), .A3(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1233), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1240), .B(new_n1231), .C1(new_n1245), .C2(new_n1242), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT61), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1244), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT126), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G378), .B(new_n1203), .C1(new_n1168), .C2(new_n1175), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1169), .A2(new_n730), .A3(new_n1174), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1172), .A2(new_n961), .A3(new_n1202), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1251), .A2(new_n1252), .A3(new_n1200), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1230), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1250), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT123), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n658), .A2(G213), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT124), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT60), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n682), .B1(new_n1226), .B2(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1261), .B(new_n1108), .C1(new_n1260), .C2(new_n1226), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1225), .ZN(new_n1263));
  INV_X1    g1063(.A(G384), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1259), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  AOI211_X1 g1065(.A(KEYINPUT124), .B(G384), .C1(new_n1262), .C2(new_n1225), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1250), .A2(KEYINPUT123), .A3(new_n1254), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1257), .A2(new_n1258), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n1271));
  OR2_X1    g1071(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1257), .A2(new_n1258), .A3(new_n1269), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n658), .A2(G213), .A3(G2897), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1268), .B(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1250), .A2(new_n1254), .B1(G213), .B2(new_n658), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1268), .A2(KEYINPUT63), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n1274), .A2(new_n1277), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1249), .A2(new_n1273), .A3(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1247), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1255), .A2(KEYINPUT62), .A3(new_n1258), .A4(new_n1268), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT127), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1278), .A2(KEYINPUT127), .A3(KEYINPUT62), .A4(new_n1268), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT62), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1270), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1282), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1281), .B1(new_n1290), .B2(new_n1292), .ZN(G405));
  XNOR2_X1  g1093(.A(new_n1291), .B(new_n1268), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G375), .A2(new_n1230), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1250), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(new_n1294), .B(new_n1296), .ZN(G402));
endmodule


