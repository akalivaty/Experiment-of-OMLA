//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  INV_X1    g000(.A(KEYINPUT6), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT87), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n189), .A2(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT4), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G101), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT80), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n195), .A2(KEYINPUT80), .A3(new_n196), .A4(G101), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n190), .A2(new_n193), .A3(new_n201), .A4(new_n194), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT79), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n195), .A2(G101), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT4), .B1(new_n205), .B2(KEYINPUT79), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n199), .B(new_n200), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n209));
  INV_X1    g023(.A(G116), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G119), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(G119), .ZN(new_n212));
  INV_X1    g026(.A(G119), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT66), .A3(G116), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT2), .B(G113), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n211), .A2(new_n214), .A3(KEYINPUT67), .A4(new_n212), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n217), .B1(new_n221), .B2(new_n216), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n188), .B1(new_n208), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n207), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n204), .A2(new_n205), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n199), .A2(new_n200), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n221), .A2(new_n216), .ZN(new_n229));
  INV_X1    g043(.A(new_n217), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n226), .A2(new_n228), .A3(new_n231), .A4(KEYINPUT87), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n219), .A2(KEYINPUT5), .A3(new_n220), .ZN(new_n233));
  NOR3_X1   g047(.A1(new_n210), .A2(KEYINPUT5), .A3(G119), .ZN(new_n234));
  INV_X1    g048(.A(G113), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n233), .A2(KEYINPUT88), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT88), .B1(new_n233), .B2(new_n236), .ZN(new_n238));
  NOR3_X1   g052(.A1(new_n237), .A2(new_n238), .A3(new_n217), .ZN(new_n239));
  XNOR2_X1  g053(.A(G104), .B(G107), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT81), .B1(new_n240), .B2(new_n201), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT81), .ZN(new_n242));
  INV_X1    g056(.A(new_n194), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n189), .A2(G107), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n242), .B(G101), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n241), .A2(new_n245), .A3(new_n202), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT83), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT83), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n241), .A2(new_n245), .A3(new_n248), .A4(new_n202), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n223), .A2(new_n232), .B1(new_n239), .B2(new_n250), .ZN(new_n251));
  XOR2_X1   g065(.A(G110), .B(G122), .Z(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n187), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n223), .A2(new_n232), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n239), .A2(new_n250), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n252), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n257), .A2(new_n187), .A3(new_n252), .ZN(new_n260));
  INV_X1    g074(.A(G146), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G143), .ZN(new_n262));
  INV_X1    g076(.A(G143), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G146), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT1), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n262), .A2(new_n264), .A3(new_n265), .A4(G128), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n263), .A2(G146), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT64), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n268), .B1(new_n261), .B2(G143), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n263), .A2(KEYINPUT64), .A3(G146), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n267), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G128), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n272), .B1(new_n262), .B2(KEYINPUT1), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n266), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  OR2_X1    g088(.A1(new_n274), .A2(G125), .ZN(new_n275));
  INV_X1    g089(.A(G125), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n263), .A2(KEYINPUT64), .A3(G146), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT64), .B1(new_n263), .B2(G146), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n262), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  XOR2_X1   g093(.A(KEYINPUT0), .B(G128), .Z(new_n280));
  AND3_X1   g094(.A1(new_n262), .A2(new_n264), .A3(G128), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n279), .A2(new_n280), .B1(new_n281), .B2(KEYINPUT0), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n275), .B1(new_n276), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G224), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(G953), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n283), .B(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n259), .A2(new_n260), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT7), .B1(new_n284), .B2(G953), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n283), .B(new_n288), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n211), .A2(new_n214), .A3(KEYINPUT5), .A4(new_n212), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n217), .B1(new_n290), .B2(new_n236), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n250), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n246), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n292), .B1(new_n239), .B2(new_n293), .ZN(new_n294));
  XOR2_X1   g108(.A(new_n252), .B(KEYINPUT8), .Z(new_n295));
  AOI21_X1  g109(.A(new_n289), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n251), .A2(new_n253), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n287), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G210), .B1(G237), .B2(G902), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g116(.A1(new_n302), .A2(KEYINPUT89), .ZN(new_n303));
  OAI21_X1  g117(.A(G214), .B1(G237), .B2(G902), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n287), .A2(new_n298), .A3(new_n300), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n302), .A2(KEYINPUT89), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n303), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT90), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT71), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n311), .B(G101), .ZN(new_n312));
  NOR2_X1   g126(.A1(G237), .A2(G953), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G210), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n312), .B(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT11), .ZN(new_n316));
  INV_X1    g130(.A(G134), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(G137), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(G137), .ZN(new_n319));
  INV_X1    g133(.A(G137), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(KEYINPUT11), .A3(G134), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n318), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G131), .ZN(new_n323));
  INV_X1    g137(.A(G131), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n318), .A2(new_n321), .A3(new_n324), .A4(new_n319), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n282), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT65), .B1(new_n317), .B2(G137), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT65), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n320), .A3(G134), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n330), .A3(new_n319), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G131), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n274), .A2(new_n325), .A3(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n222), .A2(new_n327), .A3(new_n333), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n332), .A2(new_n325), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n335), .A2(new_n274), .B1(new_n282), .B2(new_n326), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n336), .A2(KEYINPUT69), .A3(new_n222), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT69), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n327), .A2(new_n333), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(new_n231), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n334), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  XOR2_X1   g155(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT70), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT28), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n334), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n344), .B1(new_n334), .B2(new_n345), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n315), .B1(new_n343), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT30), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n327), .A2(new_n350), .A3(new_n333), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n350), .B1(new_n327), .B2(new_n333), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n231), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(new_n334), .A3(new_n315), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT31), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT31), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n353), .A2(new_n356), .A3(new_n334), .A4(new_n315), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n310), .B1(new_n349), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n315), .ZN(new_n360));
  INV_X1    g174(.A(new_n342), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT69), .B1(new_n336), .B2(new_n222), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n339), .A2(new_n231), .A3(new_n338), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n361), .B1(new_n364), .B2(new_n334), .ZN(new_n365));
  INV_X1    g179(.A(new_n347), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n334), .A2(new_n344), .A3(new_n345), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n360), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n369), .A2(KEYINPUT71), .A3(new_n357), .A4(new_n355), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n359), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(G472), .A2(G902), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT73), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n372), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n378), .B1(new_n359), .B2(new_n370), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT74), .B(G902), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n339), .A2(new_n231), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n334), .ZN(new_n383));
  AOI211_X1 g197(.A(new_n347), .B(new_n346), .C1(KEYINPUT28), .C2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT29), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n362), .A2(new_n363), .B1(new_n222), .B2(new_n336), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n348), .B(new_n385), .C1(new_n361), .C2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n387), .A3(new_n315), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n353), .A2(new_n334), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(new_n315), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(new_n387), .B2(new_n315), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n381), .B(new_n388), .C1(new_n391), .C2(KEYINPUT29), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n379), .A2(KEYINPUT32), .B1(new_n392), .B2(G472), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT73), .B1(new_n379), .B2(new_n375), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n377), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n276), .A2(KEYINPUT16), .A3(G140), .ZN(new_n396));
  OR2_X1    g210(.A1(G125), .A2(G140), .ZN(new_n397));
  NAND2_X1  g211(.A1(G125), .A2(G140), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n396), .B1(new_n399), .B2(KEYINPUT16), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G146), .ZN(new_n401));
  AOI21_X1  g215(.A(G146), .B1(new_n397), .B2(new_n398), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n402), .B(KEYINPUT77), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n272), .A2(G119), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n213), .A2(G128), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  XOR2_X1   g220(.A(new_n406), .B(KEYINPUT75), .Z(new_n407));
  XOR2_X1   g221(.A(KEYINPUT24), .B(G110), .Z(new_n408));
  NOR2_X1   g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(KEYINPUT76), .B1(new_n405), .B2(KEYINPUT23), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(new_n404), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(G110), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n401), .B(new_n403), .C1(new_n409), .C2(new_n412), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n407), .A2(new_n408), .B1(new_n411), .B2(G110), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n400), .B(new_n261), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G953), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(G221), .A3(G234), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(KEYINPUT22), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(G137), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n413), .A2(new_n417), .A3(new_n422), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n381), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT25), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n428), .A2(KEYINPUT78), .ZN(new_n429));
  INV_X1    g243(.A(G217), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n430), .B1(new_n381), .B2(G234), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n424), .A2(new_n425), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(KEYINPUT25), .A3(new_n381), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(new_n428), .A3(KEYINPUT78), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n431), .A2(G902), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n433), .A2(new_n436), .B1(new_n437), .B2(new_n434), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n395), .A2(new_n438), .ZN(new_n439));
  XOR2_X1   g253(.A(KEYINPUT9), .B(G234), .Z(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G221), .B1(new_n441), .B2(G902), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G902), .ZN(new_n444));
  XNOR2_X1  g258(.A(G110), .B(G140), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n419), .A2(G227), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n445), .B(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n227), .B1(new_n225), .B2(new_n224), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT10), .ZN(new_n450));
  OAI21_X1  g264(.A(G128), .B1(new_n267), .B2(new_n265), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n262), .A2(new_n264), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n265), .A2(new_n281), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n450), .B1(new_n246), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT82), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g270(.A(KEYINPUT82), .B(new_n450), .C1(new_n246), .C2(new_n453), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n449), .A2(new_n282), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n326), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n274), .A2(KEYINPUT10), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n247), .A3(new_n249), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT84), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT84), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n460), .A2(new_n247), .A3(new_n463), .A4(new_n249), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n458), .A2(new_n459), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n274), .B1(new_n247), .B2(new_n249), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n246), .A2(new_n453), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n326), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT12), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT12), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n471), .B(new_n326), .C1(new_n467), .C2(new_n468), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n448), .B1(new_n466), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT85), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n462), .A2(new_n464), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n456), .A2(new_n457), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n226), .A2(new_n228), .A3(new_n282), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n326), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n458), .A2(new_n465), .A3(new_n459), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n481), .A3(new_n447), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n474), .A2(new_n475), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n475), .B1(new_n474), .B2(new_n482), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n444), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G469), .ZN(new_n486));
  INV_X1    g300(.A(G469), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n481), .A2(new_n470), .A3(new_n472), .A4(new_n447), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n447), .B1(new_n480), .B2(new_n481), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n487), .B(new_n381), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT86), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n459), .B1(new_n458), .B2(new_n465), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n448), .B1(new_n466), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n380), .B1(new_n494), .B2(new_n488), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT86), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n496), .A3(new_n487), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n443), .B1(new_n486), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT97), .ZN(new_n501));
  INV_X1    g315(.A(G478), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(KEYINPUT15), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G122), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G116), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n210), .A2(G122), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n508), .A2(new_n192), .ZN(new_n509));
  XNOR2_X1  g323(.A(G128), .B(G143), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(G134), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n505), .A2(G116), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT14), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n506), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT95), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n512), .A2(new_n513), .ZN(new_n517));
  OAI211_X1 g331(.A(KEYINPUT95), .B(new_n506), .C1(new_n512), .C2(new_n513), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  AOI211_X1 g333(.A(new_n509), .B(new_n511), .C1(G107), .C2(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n508), .B(new_n192), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n510), .A2(KEYINPUT13), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n263), .A2(G128), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n522), .B(G134), .C1(KEYINPUT13), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n510), .A2(new_n317), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n521), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT96), .B1(new_n520), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n509), .B1(new_n519), .B2(G107), .ZN(new_n529));
  INV_X1    g343(.A(new_n511), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT96), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(new_n526), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n441), .A2(new_n430), .A3(G953), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n528), .A2(new_n535), .A3(new_n533), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n504), .B1(new_n539), .B2(new_n381), .ZN(new_n540));
  AOI211_X1 g354(.A(new_n380), .B(new_n503), .C1(new_n537), .C2(new_n538), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n501), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n538), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n535), .B1(new_n528), .B2(new_n533), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n381), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n503), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n539), .A2(new_n381), .A3(new_n504), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(KEYINPUT97), .A3(new_n547), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n542), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(G475), .ZN(new_n550));
  INV_X1    g364(.A(G237), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(new_n419), .A3(G214), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(KEYINPUT91), .A3(new_n263), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n263), .A2(KEYINPUT91), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(G214), .A3(new_n313), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT18), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n553), .B(new_n555), .C1(new_n556), .C2(new_n324), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(KEYINPUT92), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n397), .A2(G146), .A3(new_n398), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n403), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n553), .A2(new_n555), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G131), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n558), .B(new_n560), .C1(new_n556), .C2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(KEYINPUT17), .A3(G131), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n561), .B(G131), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n415), .B(new_n564), .C1(new_n565), .C2(KEYINPUT17), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(G113), .B(G122), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(new_n189), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n563), .A2(new_n569), .A3(new_n566), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n550), .B1(new_n573), .B2(new_n444), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT19), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n399), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n397), .A2(KEYINPUT19), .A3(new_n398), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n261), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT93), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n578), .A2(new_n579), .B1(G146), .B2(new_n400), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n565), .B(new_n580), .C1(new_n579), .C2(new_n578), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n560), .B1(new_n556), .B2(new_n562), .ZN(new_n582));
  XOR2_X1   g396(.A(new_n557), .B(KEYINPUT92), .Z(new_n583));
  OAI21_X1  g397(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n570), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n572), .ZN(new_n586));
  NOR2_X1   g400(.A1(G475), .A2(G902), .ZN(new_n587));
  XOR2_X1   g401(.A(new_n587), .B(KEYINPUT94), .Z(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT20), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT20), .ZN(new_n591));
  AOI211_X1 g405(.A(new_n591), .B(new_n588), .C1(new_n585), .C2(new_n572), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n574), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n419), .A2(G952), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n594), .B1(G234), .B2(G237), .ZN(new_n595));
  AOI211_X1 g409(.A(new_n419), .B(new_n381), .C1(G234), .C2(G237), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT21), .B(G898), .Z(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n595), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n549), .A2(new_n593), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n500), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n309), .A2(new_n439), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT98), .B(G101), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G3));
  NAND2_X1  g419(.A1(new_n371), .A2(new_n381), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(G472), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n373), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(new_n438), .A3(new_n499), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n539), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n537), .A2(KEYINPUT33), .A3(new_n538), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n612), .A2(G478), .A3(new_n381), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n545), .A2(new_n502), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n593), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n304), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n302), .B2(new_n305), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n600), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n610), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT99), .B(KEYINPUT34), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G104), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n622), .B(new_n624), .ZN(G6));
  NOR4_X1   g439(.A1(new_n610), .A2(new_n617), .A3(new_n549), .A4(new_n621), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT35), .B(G107), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  NAND2_X1  g442(.A1(new_n433), .A2(new_n436), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n423), .A2(KEYINPUT36), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n418), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n437), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n309), .A2(new_n602), .A3(new_n609), .A4(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n634), .B(KEYINPUT37), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G110), .ZN(G12));
  AOI22_X1  g450(.A1(new_n485), .A2(G469), .B1(new_n492), .B2(new_n497), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n287), .A2(new_n300), .A3(new_n298), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n300), .B1(new_n287), .B2(new_n298), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n304), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n637), .A2(new_n640), .A3(new_n443), .ZN(new_n641));
  INV_X1    g455(.A(G900), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n595), .B1(new_n596), .B2(new_n642), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n549), .A2(new_n617), .A3(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n641), .A2(new_n395), .A3(new_n633), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G128), .ZN(G30));
  XNOR2_X1  g460(.A(new_n643), .B(KEYINPUT39), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n499), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT100), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n649), .A2(KEYINPUT100), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n593), .B1(new_n542), .B2(new_n548), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n303), .A2(new_n306), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT38), .ZN(new_n659));
  OR2_X1    g473(.A1(new_n651), .A2(new_n652), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n659), .B1(new_n660), .B2(KEYINPUT40), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n379), .A2(KEYINPUT32), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n389), .A2(new_n315), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n444), .B1(new_n383), .B2(new_n315), .ZN(new_n665));
  OAI21_X1  g479(.A(G472), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n377), .A2(new_n394), .A3(new_n662), .A4(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n633), .A2(new_n619), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n657), .A2(new_n661), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G143), .ZN(G45));
  INV_X1    g484(.A(new_n643), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n616), .A2(new_n617), .A3(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n641), .A2(new_n395), .A3(new_n633), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G146), .ZN(G48));
  NOR2_X1   g489(.A1(new_n621), .A2(new_n618), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n495), .A2(new_n487), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n492), .B2(new_n497), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(new_n443), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n439), .A2(new_n676), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  NOR3_X1   g497(.A1(new_n621), .A2(new_n617), .A3(new_n549), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(new_n439), .A3(new_n680), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  AND2_X1   g500(.A1(new_n395), .A2(new_n633), .ZN(new_n687));
  INV_X1    g501(.A(new_n601), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n620), .A2(new_n442), .A3(new_n678), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n687), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G119), .ZN(G21));
  INV_X1    g506(.A(KEYINPUT101), .ZN(new_n693));
  INV_X1    g507(.A(new_n656), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n693), .B1(new_n640), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n620), .A2(KEYINPUT101), .A3(new_n656), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n384), .A2(new_n315), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n372), .B1(new_n698), .B2(new_n358), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n607), .A2(new_n438), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n697), .A2(new_n600), .A3(new_n680), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G122), .ZN(G24));
  NAND3_X1  g517(.A1(new_n607), .A2(new_n633), .A3(new_n699), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n689), .A2(new_n672), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n276), .ZN(G27));
  NOR2_X1   g520(.A1(new_n443), .A2(new_n619), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n658), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n474), .A2(KEYINPUT102), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT102), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n711), .B(new_n448), .C1(new_n466), .C2(new_n473), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n710), .A2(new_n482), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n444), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(G469), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n498), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n709), .A2(KEYINPUT42), .A3(new_n673), .A4(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n438), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n379), .A2(KEYINPUT32), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n718), .B1(new_n720), .B2(new_n393), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(KEYINPUT103), .B1(new_n717), .B2(new_n722), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n714), .A2(G469), .B1(new_n492), .B2(new_n497), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n708), .A2(new_n672), .A3(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT103), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n725), .A2(new_n726), .A3(KEYINPUT42), .A4(new_n721), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n708), .A2(new_n724), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n439), .A3(new_n673), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G131), .ZN(G33));
  NAND3_X1  g548(.A1(new_n729), .A2(new_n439), .A3(new_n644), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G134), .ZN(G36));
  NAND2_X1  g550(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n616), .A2(new_n593), .ZN(new_n739));
  MUX2_X1   g553(.A(new_n737), .B(new_n738), .S(new_n739), .Z(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n608), .A3(new_n633), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n658), .A2(new_n304), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n741), .B2(new_n742), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n746), .B1(new_n483), .B2(new_n484), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n747), .B(G469), .C1(new_n746), .C2(new_n713), .ZN(new_n748));
  NAND2_X1  g562(.A1(G469), .A2(G902), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT46), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n497), .B2(new_n492), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n748), .A2(KEYINPUT46), .A3(new_n749), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n443), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n743), .A2(new_n745), .A3(new_n648), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G137), .ZN(G39));
  AND2_X1   g569(.A1(new_n753), .A2(KEYINPUT47), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n753), .A2(KEYINPUT47), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n744), .A2(new_n395), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n758), .A2(new_n718), .A3(new_n673), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G140), .ZN(G42));
  XNOR2_X1  g575(.A(new_n678), .B(KEYINPUT49), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n659), .A2(new_n438), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n667), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n763), .A2(new_n764), .A3(new_n707), .A4(new_n739), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n740), .A2(new_n595), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n766), .A2(new_n701), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n767), .A2(new_n619), .A3(new_n659), .A4(new_n680), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n709), .A2(new_n678), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n764), .A2(new_n595), .ZN(new_n772));
  NOR4_X1   g586(.A1(new_n771), .A2(new_n772), .A3(new_n718), .A4(new_n616), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n766), .A2(new_n678), .A3(new_n709), .ZN(new_n774));
  INV_X1    g588(.A(new_n704), .ZN(new_n775));
  AOI22_X1  g589(.A1(new_n593), .A2(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AOI211_X1 g590(.A(new_n757), .B(new_n756), .C1(new_n443), .C2(new_n678), .ZN(new_n777));
  INV_X1    g591(.A(new_n744), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n767), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n770), .B(new_n776), .C1(new_n777), .C2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT108), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n780), .A2(new_n781), .A3(KEYINPUT51), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n594), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n610), .A2(new_n599), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n593), .A2(new_n546), .A3(new_n547), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n616), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n789), .B1(new_n790), .B2(new_n617), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n309), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n634), .A2(new_n603), .A3(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n685), .A2(new_n681), .A3(new_n691), .A4(new_n702), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n788), .A2(new_n643), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n500), .B1(new_n796), .B2(KEYINPUT105), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n796), .A2(KEYINPUT105), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n797), .A2(new_n687), .A3(new_n778), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n704), .A2(new_n672), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n729), .A2(new_n800), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n799), .A2(new_n735), .A3(new_n801), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n795), .A2(new_n733), .A3(new_n802), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n724), .A2(new_n443), .A3(new_n633), .A4(new_n643), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n697), .A2(new_n804), .A3(new_n667), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n690), .A2(new_n800), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(new_n645), .A3(new_n674), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT52), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT106), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n633), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n716), .A2(new_n442), .A3(new_n812), .A4(new_n671), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n764), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n705), .B1(new_n814), .B2(new_n697), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n687), .B(new_n641), .C1(new_n644), .C2(new_n673), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT106), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n809), .B1(new_n811), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n803), .A2(KEYINPUT53), .A3(new_n808), .A4(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n795), .A2(new_n733), .A3(new_n802), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT107), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n695), .A2(new_n696), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n633), .B1(new_n715), .B2(new_n498), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n667), .A2(new_n823), .A3(new_n442), .A4(new_n671), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n806), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n395), .A2(new_n499), .A3(new_n620), .A4(new_n633), .ZN(new_n826));
  INV_X1    g640(.A(new_n644), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n826), .B1(new_n827), .B2(new_n672), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n810), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n816), .A2(KEYINPUT106), .A3(new_n806), .A4(new_n805), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n829), .A2(KEYINPUT52), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT52), .B1(new_n829), .B2(new_n830), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n821), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n829), .A2(KEYINPUT52), .A3(new_n830), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n818), .A2(KEYINPUT107), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n820), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n819), .B1(new_n836), .B2(KEYINPUT53), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n837), .A2(KEYINPUT54), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n767), .A2(new_n690), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n836), .A2(KEYINPUT53), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n820), .A2(new_n832), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT53), .B1(new_n841), .B2(new_n808), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT54), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n786), .A2(new_n838), .A3(new_n839), .A4(new_n843), .ZN(new_n844));
  NOR4_X1   g658(.A1(new_n771), .A2(new_n772), .A3(new_n718), .A4(new_n618), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n774), .A2(new_n721), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n846), .B(KEYINPUT48), .Z(new_n847));
  NOR3_X1   g661(.A1(new_n844), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(G952), .A2(G953), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n765), .B1(new_n848), .B2(new_n849), .ZN(G75));
  NAND2_X1  g664(.A1(new_n833), .A2(new_n835), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT53), .B1(new_n851), .B2(new_n803), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  INV_X1    g667(.A(new_n808), .ZN(new_n854));
  NOR4_X1   g668(.A1(new_n820), .A2(new_n853), .A3(new_n854), .A4(new_n832), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n380), .B(new_n301), .C1(new_n852), .C2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT56), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n259), .A2(new_n260), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT109), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n286), .B(KEYINPUT55), .Z(new_n860));
  XOR2_X1   g674(.A(new_n859), .B(new_n860), .Z(new_n861));
  NAND3_X1  g675(.A1(new_n856), .A2(new_n857), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT112), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT112), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n856), .A2(new_n864), .A3(new_n857), .A4(new_n861), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n419), .A2(G952), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT110), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n856), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n837), .A2(KEYINPUT110), .A3(new_n380), .A4(new_n301), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n857), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT111), .ZN(new_n874));
  INV_X1    g688(.A(new_n861), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n873), .A2(new_n875), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT111), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n869), .B1(new_n876), .B2(new_n878), .ZN(G51));
  NAND2_X1  g693(.A1(new_n494), .A2(new_n488), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT113), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n837), .B(KEYINPUT54), .Z(new_n882));
  XNOR2_X1  g696(.A(new_n749), .B(KEYINPUT57), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n837), .A2(new_n380), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n748), .B(KEYINPUT114), .Z(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n867), .B1(new_n884), .B2(new_n887), .ZN(G54));
  NAND3_X1  g702(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT115), .ZN(new_n890));
  INV_X1    g704(.A(new_n586), .ZN(new_n891));
  OR3_X1    g705(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n867), .B1(new_n889), .B2(new_n891), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n890), .B1(new_n889), .B2(new_n891), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(G60));
  XOR2_X1   g709(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n896));
  NOR2_X1   g710(.A1(new_n502), .A2(new_n444), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n896), .B(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n838), .B2(new_n843), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n613), .B2(new_n612), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n612), .A2(new_n613), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n882), .A2(new_n902), .A3(new_n899), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n901), .A2(new_n903), .A3(new_n867), .ZN(G63));
  NAND2_X1  g718(.A1(G217), .A2(G902), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT60), .Z(new_n906));
  NAND3_X1  g720(.A1(new_n837), .A2(new_n631), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT117), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n908), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n434), .B1(new_n837), .B2(new_n906), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n912), .A2(KEYINPUT118), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n912), .B2(KEYINPUT118), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n911), .A2(new_n868), .A3(new_n913), .A4(new_n915), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n912), .A2(new_n867), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n917), .B1(new_n910), .B2(new_n909), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n916), .B1(KEYINPUT61), .B2(new_n918), .ZN(G66));
  NOR2_X1   g733(.A1(new_n795), .A2(G953), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT119), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n419), .B1(new_n597), .B2(G224), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n923), .B1(new_n921), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n859), .B1(G898), .B2(new_n419), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT120), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n924), .B(new_n926), .ZN(G69));
  OR2_X1    g741(.A1(new_n351), .A2(new_n352), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n576), .A2(new_n577), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n928), .B(new_n929), .Z(new_n930));
  AOI21_X1  g744(.A(new_n419), .B1(G227), .B2(G900), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n828), .A2(new_n705), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(new_n669), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT122), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n669), .A2(new_n933), .A3(new_n934), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT121), .ZN(new_n938));
  INV_X1    g752(.A(new_n760), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n653), .A2(new_n439), .A3(new_n791), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n754), .B1(new_n744), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT123), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n939), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n936), .A2(new_n938), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n932), .B1(new_n946), .B2(G953), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n760), .A2(new_n733), .A3(new_n735), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n753), .A2(new_n648), .A3(new_n697), .A4(new_n721), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n754), .A2(new_n934), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT124), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(KEYINPUT125), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n948), .A2(new_n954), .A3(new_n949), .A4(new_n951), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n953), .A2(new_n955), .A3(new_n419), .ZN(new_n956));
  OAI21_X1  g770(.A(G953), .B1(new_n642), .B2(G227), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n956), .A2(new_n930), .A3(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT126), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n947), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n959), .B1(new_n947), .B2(new_n958), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n960), .A2(new_n961), .ZN(G72));
  NAND3_X1  g776(.A1(new_n953), .A2(new_n955), .A3(new_n795), .ZN(new_n963));
  NAND2_X1  g777(.A1(G472), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT63), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n390), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n664), .A2(new_n390), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n965), .B(new_n968), .C1(new_n840), .C2(new_n842), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n967), .A2(new_n868), .A3(new_n969), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n936), .A2(new_n938), .A3(new_n795), .A4(new_n945), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n971), .A2(KEYINPUT127), .A3(new_n965), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT127), .B1(new_n971), .B2(new_n965), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n972), .A2(new_n973), .A3(new_n663), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n970), .A2(new_n974), .ZN(G57));
endmodule


