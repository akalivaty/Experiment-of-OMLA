//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n569, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n619, new_n620, new_n622, new_n623, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n464), .A3(G125), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n465), .A2(new_n466), .B1(G113), .B2(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n462), .A2(new_n464), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(KEYINPUT67), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n472), .A2(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT68), .B1(new_n463), .B2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(new_n461), .A3(KEYINPUT3), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n473), .A2(new_n474), .A3(new_n476), .A4(new_n464), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT69), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n461), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G101), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n471), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT70), .Z(G160));
  NAND3_X1  g057(.A1(new_n474), .A2(new_n476), .A3(new_n464), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n483), .B(new_n484), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n485), .A2(new_n472), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n485), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT72), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n487), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  NOR3_X1   g069(.A1(new_n463), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AND2_X1   g072(.A1(G126), .A2(G2105), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n497), .A2(KEYINPUT73), .A3(new_n474), .A4(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n474), .A2(new_n476), .A3(new_n464), .A4(new_n498), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT73), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G138), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(G2105), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n474), .A2(new_n476), .A3(new_n464), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n468), .A2(new_n508), .A3(new_n505), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT74), .B(G114), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(G2105), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n503), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT75), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n526), .B1(new_n522), .B2(new_n523), .ZN(new_n527));
  OAI21_X1  g102(.A(G651), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n520), .A2(new_n521), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  AND2_X1   g105(.A1(KEYINPUT6), .A2(G651), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G88), .ZN(new_n533));
  INV_X1    g108(.A(G50), .ZN(new_n534));
  OAI21_X1  g109(.A(G543), .B1(new_n531), .B2(new_n530), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n532), .A2(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n528), .A2(new_n537), .ZN(G303));
  INV_X1    g113(.A(G303), .ZN(G166));
  NAND3_X1  g114(.A1(new_n529), .A2(G63), .A3(G651), .ZN(new_n540));
  INV_X1    g115(.A(new_n535), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G51), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  INV_X1    g119(.A(G89), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n532), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n540), .B(new_n542), .C1(new_n546), .C2(KEYINPUT76), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n546), .A2(KEYINPUT76), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(G168));
  INV_X1    g124(.A(new_n532), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n550), .A2(G90), .B1(new_n541), .B2(G52), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n529), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G651), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AND2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(G171));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(new_n529), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n553), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n561), .B1(new_n560), .B2(new_n559), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n550), .A2(G81), .B1(new_n541), .B2(G43), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT78), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g143(.A(KEYINPUT79), .B(KEYINPUT8), .Z(new_n569));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  NAND2_X1  g147(.A1(new_n541), .A2(G53), .ZN(new_n573));
  XOR2_X1   g148(.A(new_n573), .B(KEYINPUT9), .Z(new_n574));
  AOI22_X1  g149(.A1(new_n529), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G91), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n575), .A2(new_n553), .B1(new_n532), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G299));
  XNOR2_X1  g154(.A(G171), .B(KEYINPUT80), .ZN(G301));
  INV_X1    g155(.A(G168), .ZN(G286));
  NAND2_X1  g156(.A1(new_n550), .A2(G87), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n541), .A2(G49), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n529), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT81), .ZN(G288));
  NAND2_X1  g161(.A1(new_n529), .A2(G61), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n553), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(KEYINPUT82), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(KEYINPUT82), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n550), .A2(G86), .B1(new_n541), .B2(G48), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(G305));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  INV_X1    g170(.A(G47), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n532), .A2(new_n595), .B1(new_n596), .B2(new_n535), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n529), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n553), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G290));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OR3_X1    g177(.A1(new_n532), .A2(KEYINPUT83), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(KEYINPUT83), .B1(new_n532), .B2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n603), .A2(KEYINPUT10), .A3(new_n604), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  XOR2_X1   g184(.A(KEYINPUT84), .B(G66), .Z(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n557), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n611), .A2(G651), .B1(G54), .B2(new_n541), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n607), .A2(new_n608), .A3(new_n612), .ZN(new_n613));
  MUX2_X1   g188(.A(new_n613), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g189(.A(new_n613), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n578), .ZN(G297));
  OAI21_X1  g192(.A(new_n616), .B1(G868), .B2(new_n578), .ZN(G280));
  AND3_X1   g193(.A1(new_n607), .A2(new_n608), .A3(new_n612), .ZN(new_n619));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n565), .ZN(G323));
  XNOR2_X1  g199(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n625));
  XNOR2_X1  g200(.A(G323), .B(new_n625), .ZN(G282));
  NAND2_X1  g201(.A1(new_n468), .A2(new_n479), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n486), .A2(G135), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n488), .A2(G123), .ZN(new_n632));
  OR2_X1    g207(.A1(G99), .A2(G2105), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n633), .B(G2104), .C1(G111), .C2(new_n472), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n635), .A2(G2096), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(G2096), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n630), .A2(new_n636), .A3(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n644), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT86), .ZN(new_n652));
  OAI21_X1  g227(.A(G14), .B1(new_n649), .B2(new_n650), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(G401));
  INV_X1    g229(.A(KEYINPUT18), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT17), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2100), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n658), .B2(KEYINPUT18), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2096), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(G227));
  XOR2_X1   g241(.A(G1971), .B(G1976), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1961), .B(G1966), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT20), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n668), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n668), .B2(new_n674), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(G1981), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G1986), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT87), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G229));
  NAND2_X1  g260(.A1(G166), .A2(G16), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(G16), .B2(G22), .ZN(new_n687));
  INV_X1    g262(.A(G1971), .ZN(new_n688));
  OR2_X1    g263(.A1(G6), .A2(G16), .ZN(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(G305), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT32), .B(G1981), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  AOI22_X1  g268(.A1(new_n687), .A2(new_n688), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(new_n688), .B2(new_n687), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n690), .A2(G23), .ZN(new_n696));
  INV_X1    g271(.A(new_n585), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n690), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT33), .B(G1976), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n691), .A2(new_n693), .ZN(new_n701));
  NOR3_X1   g276(.A1(new_n695), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT34), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  NOR2_X1   g280(.A1(G25), .A2(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n488), .A2(G119), .ZN(new_n707));
  OR2_X1    g282(.A1(G95), .A2(G2105), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n708), .B(G2104), .C1(G107), .C2(new_n472), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G131), .B2(new_n486), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n706), .B1(new_n711), .B2(G29), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT35), .B(G1991), .Z(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n690), .A2(G24), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n600), .B2(new_n690), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1986), .ZN(new_n718));
  INV_X1    g293(.A(new_n712), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(new_n713), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n704), .A2(new_n705), .A3(new_n715), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT36), .ZN(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G26), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT28), .Z(new_n725));
  NAND2_X1  g300(.A1(new_n486), .A2(G140), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT88), .ZN(new_n727));
  OAI21_X1  g302(.A(G2104), .B1(new_n472), .B2(G116), .ZN(new_n728));
  OR3_X1    g303(.A1(KEYINPUT89), .A2(G104), .A3(G2105), .ZN(new_n729));
  OAI21_X1  g304(.A(KEYINPUT89), .B1(G104), .B2(G2105), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n488), .B2(G128), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n725), .B1(new_n733), .B2(G29), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G2067), .ZN(new_n735));
  NOR2_X1   g310(.A1(G4), .A2(G16), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n619), .B2(G16), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G1348), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(G1348), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n690), .A2(G19), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n565), .B2(new_n690), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(G1341), .Z(new_n742));
  NAND4_X1  g317(.A1(new_n735), .A2(new_n738), .A3(new_n739), .A4(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT90), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n723), .A2(G35), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G162), .B2(new_n723), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT29), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G2090), .ZN(new_n748));
  NAND2_X1  g323(.A1(G168), .A2(G16), .ZN(new_n749));
  NOR2_X1   g324(.A1(G16), .A2(G21), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(KEYINPUT92), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(KEYINPUT92), .B2(new_n749), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1966), .ZN(new_n753));
  NOR2_X1   g328(.A1(G164), .A2(new_n723), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G27), .B2(new_n723), .ZN(new_n755));
  INV_X1    g330(.A(G2078), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n690), .A2(G5), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G171), .B2(new_n690), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(G1961), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n690), .A2(G20), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT23), .Z(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G299), .B2(G16), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1956), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n753), .A2(new_n757), .A3(new_n760), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n723), .A2(G32), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n486), .A2(G141), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n488), .A2(G129), .ZN(new_n768));
  NAND3_X1  g343(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT26), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n771), .A2(new_n772), .B1(G105), .B2(new_n479), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n767), .A2(new_n768), .A3(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n766), .B1(new_n775), .B2(new_n723), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT27), .B(G1996), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT30), .B(G28), .ZN(new_n779));
  OR2_X1    g354(.A1(KEYINPUT31), .A2(G11), .ZN(new_n780));
  NAND2_X1  g355(.A1(KEYINPUT31), .A2(G11), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n779), .A2(new_n723), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n635), .B2(new_n723), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT93), .Z(new_n784));
  AND2_X1   g359(.A1(new_n723), .A2(G33), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n486), .A2(G139), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n468), .A2(G127), .ZN(new_n787));
  INV_X1    g362(.A(G115), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n461), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT25), .ZN(new_n790));
  NAND2_X1  g365(.A1(G103), .A2(G2104), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(G2105), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n472), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n789), .A2(G2105), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n786), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n785), .B1(new_n795), .B2(G29), .ZN(new_n796));
  INV_X1    g371(.A(G2072), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n755), .A2(new_n756), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n784), .A2(new_n798), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NOR4_X1   g376(.A1(new_n748), .A2(new_n765), .A3(new_n778), .A4(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G34), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n803), .A2(KEYINPUT24), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(KEYINPUT24), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n723), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G160), .B2(new_n723), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT91), .ZN(new_n808));
  INV_X1    g383(.A(G2084), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n722), .A2(new_n744), .A3(new_n802), .A4(new_n810), .ZN(G150));
  INV_X1    g386(.A(G150), .ZN(G311));
  NOR2_X1   g387(.A1(new_n613), .A2(new_n620), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(G93), .ZN(new_n816));
  INV_X1    g391(.A(G55), .ZN(new_n817));
  OAI22_X1  g392(.A1(new_n532), .A2(new_n816), .B1(new_n817), .B2(new_n535), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n529), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(new_n553), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n564), .B(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n815), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT39), .ZN(new_n824));
  AOI21_X1  g399(.A(G860), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n824), .B2(new_n823), .ZN(new_n826));
  OAI21_X1  g401(.A(G860), .B1(new_n818), .B2(new_n820), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT37), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT95), .ZN(G145));
  AND2_X1   g405(.A1(new_n727), .A2(new_n732), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G164), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n733), .A2(new_n515), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n795), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n832), .A2(new_n795), .A3(new_n833), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n835), .A2(new_n775), .A3(new_n836), .ZN(new_n837));
  AND3_X1   g412(.A1(new_n832), .A2(new_n795), .A3(new_n833), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n774), .B1(new_n838), .B2(new_n834), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n486), .A2(G142), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n488), .A2(G130), .ZN(new_n842));
  OR3_X1    g417(.A1(new_n472), .A2(KEYINPUT96), .A3(G118), .ZN(new_n843));
  OAI21_X1  g418(.A(KEYINPUT96), .B1(new_n472), .B2(G118), .ZN(new_n844));
  OR2_X1    g419(.A1(G106), .A2(G2105), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n843), .A2(G2104), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n841), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n628), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n848), .A2(new_n711), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n711), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT97), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n849), .A2(KEYINPUT97), .A3(new_n850), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n840), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n837), .A2(new_n839), .A3(new_n850), .A4(new_n849), .ZN(new_n858));
  XNOR2_X1  g433(.A(G160), .B(new_n493), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n635), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n857), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n857), .A2(KEYINPUT99), .A3(new_n858), .A4(new_n860), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G37), .ZN(new_n866));
  INV_X1    g441(.A(new_n860), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n855), .A2(new_n837), .A3(new_n839), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n855), .B1(new_n837), .B2(new_n839), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT98), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n840), .A2(new_n856), .A3(new_n870), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n867), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n865), .A2(new_n866), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n865), .A2(new_n866), .A3(new_n874), .A4(new_n876), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(G395));
  XNOR2_X1  g455(.A(G305), .B(new_n600), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n697), .B(G303), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n883), .A2(KEYINPUT42), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(KEYINPUT103), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(new_n888), .B2(new_n887), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n822), .B(new_n622), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT101), .B1(new_n619), .B2(G299), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n619), .A2(G299), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n613), .A2(new_n578), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n892), .B1(new_n895), .B2(KEYINPUT101), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(KEYINPUT41), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT102), .ZN(new_n899));
  INV_X1    g474(.A(new_n895), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n899), .B1(new_n900), .B2(KEYINPUT41), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(KEYINPUT102), .B2(new_n898), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n897), .B1(new_n903), .B2(new_n891), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n890), .B(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(G868), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(G868), .B2(new_n821), .ZN(G295));
  OAI21_X1  g482(.A(new_n906), .B1(G868), .B2(new_n821), .ZN(G331));
  NAND2_X1  g483(.A1(G301), .A2(G168), .ZN(new_n909));
  NAND2_X1  g484(.A1(G286), .A2(G171), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(G286), .A2(KEYINPUT105), .A3(G171), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n909), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n822), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT106), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n914), .A2(new_n822), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n916), .B(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n896), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n917), .A2(new_n915), .ZN(new_n920));
  AOI22_X1  g495(.A1(new_n918), .A2(new_n903), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n885), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(G37), .B1(new_n921), .B2(new_n922), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT43), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n918), .A2(new_n896), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n896), .A2(KEYINPUT41), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n929));
  AOI22_X1  g504(.A1(new_n928), .A2(new_n929), .B1(KEYINPUT41), .B2(new_n900), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT107), .B1(new_n896), .B2(KEYINPUT41), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n920), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n885), .B1(new_n927), .B2(new_n932), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n925), .A2(KEYINPUT43), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT44), .B1(new_n926), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n925), .A2(new_n933), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n936), .B1(new_n924), .B2(new_n925), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n935), .B1(new_n940), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g516(.A(G1384), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n515), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT45), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n471), .A2(new_n478), .A3(G40), .A4(new_n480), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G2067), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n831), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n733), .A2(G2067), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n947), .B1(new_n951), .B2(new_n774), .ZN(new_n952));
  INV_X1    g527(.A(new_n947), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n953), .A2(G1996), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT46), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT127), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n952), .B(new_n956), .C1(KEYINPUT46), .C2(new_n954), .ZN(new_n957));
  XOR2_X1   g532(.A(new_n957), .B(KEYINPUT47), .Z(new_n958));
  XNOR2_X1  g533(.A(new_n733), .B(new_n948), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT108), .B1(new_n959), .B2(new_n953), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n951), .A2(new_n961), .A3(new_n947), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n774), .B(G1996), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n960), .A2(new_n962), .B1(new_n947), .B2(new_n963), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n711), .A2(new_n713), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n953), .B1(new_n966), .B2(new_n949), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n711), .A2(new_n713), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n947), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n963), .A2(new_n947), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n959), .A2(KEYINPUT108), .A3(new_n953), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n961), .B1(new_n951), .B2(new_n947), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n969), .B(new_n970), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n953), .A2(G1986), .A3(G290), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT48), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n958), .A2(new_n967), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n600), .B(G1986), .Z(new_n979));
  NAND2_X1  g554(.A1(new_n947), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n978), .B1(new_n973), .B2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n964), .A2(KEYINPUT109), .A3(new_n980), .A4(new_n969), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n578), .B(KEYINPUT57), .ZN(new_n985));
  INV_X1    g560(.A(G1956), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n943), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n513), .B1(new_n499), .B2(new_n502), .ZN(new_n990));
  AOI21_X1  g565(.A(G1384), .B1(new_n990), .B2(new_n510), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT110), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n987), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n946), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(KEYINPUT50), .B2(new_n943), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n986), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n946), .B1(new_n943), .B2(new_n944), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n991), .A2(KEYINPUT45), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT56), .B(G2072), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n985), .B1(new_n996), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n989), .A2(new_n992), .A3(new_n994), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n989), .A2(new_n992), .A3(KEYINPUT118), .A4(new_n994), .ZN(new_n1005));
  AOI21_X1  g580(.A(G2067), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT119), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n989), .A2(new_n992), .A3(KEYINPUT111), .A4(new_n987), .ZN(new_n1008));
  AOI211_X1 g583(.A(new_n988), .B(G1384), .C1(new_n990), .C2(new_n510), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT110), .B1(new_n515), .B2(new_n942), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n1009), .A2(new_n1010), .A3(KEYINPUT50), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT111), .B1(new_n991), .B2(new_n987), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1008), .B(new_n994), .C1(new_n1011), .C2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT120), .ZN(new_n1015));
  INV_X1    g590(.A(G1348), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n989), .A2(new_n987), .A3(new_n992), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n1012), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT120), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1018), .A2(new_n1019), .A3(new_n1008), .A4(new_n994), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1015), .A2(new_n1016), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1007), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT50), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n946), .B1(new_n987), .B2(new_n991), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1956), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n578), .B(new_n1026), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1028));
  NOR3_X1   g603(.A1(new_n1025), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(new_n613), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1001), .B1(new_n1022), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT60), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1021), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n948), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT119), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT119), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1006), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1032), .B1(new_n1033), .B2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1021), .A2(new_n1036), .A3(KEYINPUT60), .A4(new_n1038), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1040), .A2(new_n619), .A3(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1007), .A2(KEYINPUT60), .A3(new_n613), .A4(new_n1021), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT61), .B1(new_n1029), .B2(new_n1001), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n996), .A2(new_n985), .A3(new_n1000), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1027), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT61), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1049));
  XOR2_X1   g624(.A(KEYINPUT58), .B(G1341), .Z(new_n1050));
  NAND3_X1  g625(.A1(new_n1004), .A2(new_n1005), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT121), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G1996), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n997), .A2(new_n1054), .A3(new_n998), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1004), .A2(KEYINPUT121), .A3(new_n1005), .A4(new_n1050), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1057), .A2(new_n1058), .A3(new_n565), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1058), .B1(new_n1057), .B2(new_n565), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1043), .B(new_n1049), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1031), .B1(new_n1042), .B2(new_n1061), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT122), .B(G1961), .Z(new_n1063));
  NAND3_X1  g638(.A1(new_n1015), .A2(new_n1020), .A3(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n945), .A2(new_n998), .A3(new_n756), .A4(new_n994), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT123), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1067), .B(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n998), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(new_n1066), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n944), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1071), .A2(new_n1072), .A3(new_n756), .A4(new_n994), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1064), .A2(new_n1069), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G301), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n997), .B(KEYINPUT124), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT125), .B(G2078), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1071), .A3(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1064), .A2(new_n1079), .A3(G301), .A4(new_n1069), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT54), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1018), .A2(new_n809), .A3(new_n1008), .A4(new_n994), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1072), .A2(new_n994), .A3(new_n998), .ZN(new_n1083));
  INV_X1    g658(.A(G1966), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1082), .A2(new_n1085), .A3(G168), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(G8), .ZN(new_n1087));
  AOI21_X1  g662(.A(G168), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT51), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1086), .A2(new_n1090), .A3(G8), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G8), .ZN(new_n1093));
  INV_X1    g668(.A(new_n997), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n688), .B1(new_n1094), .B2(new_n1070), .ZN(new_n1095));
  INV_X1    g670(.A(G2090), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1023), .A2(new_n1096), .A3(new_n1024), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1093), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1099));
  INV_X1    g674(.A(new_n527), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n553), .B1(new_n1100), .B2(new_n524), .ZN(new_n1101));
  OAI211_X1 g676(.A(KEYINPUT55), .B(G8), .C1(new_n1101), .C2(new_n536), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT112), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT112), .ZN(new_n1104));
  NAND4_X1  g679(.A1(G303), .A2(new_n1104), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1099), .B1(new_n1106), .B2(KEYINPUT113), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT113), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1103), .A2(new_n1105), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1098), .A2(new_n1110), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1107), .A2(KEYINPUT114), .A3(new_n1109), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT114), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1018), .A2(new_n1096), .A3(new_n1008), .A4(new_n994), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1093), .B1(new_n1115), .B2(new_n1095), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1111), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT116), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT115), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1009), .A2(new_n1010), .A3(new_n946), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1119), .B1(new_n1120), .B2(new_n1093), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1002), .A2(KEYINPUT115), .A3(G8), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1121), .A2(new_n1122), .B1(G1976), .B2(new_n697), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT52), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1118), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n697), .A2(G1976), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1002), .A2(KEYINPUT115), .A3(G8), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT115), .B1(new_n1002), .B2(G8), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1129), .A2(KEYINPUT116), .A3(KEYINPUT52), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n593), .A2(new_n592), .ZN(new_n1132));
  OAI21_X1  g707(.A(G1981), .B1(new_n1132), .B2(new_n590), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT49), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n591), .A2(new_n678), .A3(new_n593), .A4(new_n592), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1134), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1138), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1139));
  INV_X1    g714(.A(G1976), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT52), .B1(G288), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1139), .B1(new_n1123), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1117), .A2(new_n1131), .A3(new_n1142), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1081), .A2(new_n1092), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1064), .A2(new_n1079), .A3(new_n1069), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(G171), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1146), .B(KEYINPUT54), .C1(new_n1075), .C2(new_n1074), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1062), .A2(new_n1144), .A3(new_n1147), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1123), .A2(new_n1118), .A3(new_n1124), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT116), .B1(new_n1129), .B2(KEYINPUT52), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1142), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1152));
  NOR2_X1   g727(.A1(G286), .A2(new_n1093), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1152), .B(new_n1153), .C1(new_n1116), .C2(new_n1110), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT63), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1113), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1107), .A2(KEYINPUT114), .A3(new_n1109), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1116), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT63), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1160), .B1(new_n1098), .B2(new_n1110), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1158), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1162), .A2(new_n1131), .A3(new_n1142), .ZN(new_n1163));
  NOR2_X1   g738(.A1(G288), .A2(G1976), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1135), .B1(new_n1139), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT117), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1166), .A2(new_n1167), .B1(new_n1122), .B2(new_n1121), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1168), .B1(new_n1167), .B2(new_n1166), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1155), .A2(new_n1163), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1171), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1172), .A2(new_n1143), .A3(new_n1076), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1092), .A2(new_n1171), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1170), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  AOI211_X1 g750(.A(KEYINPUT126), .B(new_n984), .C1(new_n1148), .C2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT126), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1143), .A2(new_n1076), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1172), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1174), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1170), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1031), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1049), .B1(new_n1041), .B2(new_n619), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1040), .A2(new_n619), .A3(new_n1041), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1182), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1076), .A2(new_n1080), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT54), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1143), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1190), .A2(new_n1191), .A3(new_n1147), .A4(new_n1192), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1180), .B(new_n1181), .C1(new_n1187), .C2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n984), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1177), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n977), .B1(new_n1176), .B2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g772(.A(new_n925), .ZN(new_n1199));
  OAI21_X1  g773(.A(KEYINPUT43), .B1(new_n1199), .B2(new_n923), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n1200), .A2(new_n937), .ZN(new_n1201));
  NOR4_X1   g775(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1202));
  AND3_X1   g776(.A1(new_n1201), .A2(new_n875), .A3(new_n1202), .ZN(G308));
  NAND3_X1  g777(.A1(new_n1201), .A2(new_n875), .A3(new_n1202), .ZN(G225));
endmodule


