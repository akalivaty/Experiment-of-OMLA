//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n789, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988;
  XNOR2_X1  g000(.A(KEYINPUT98), .B(KEYINPUT13), .ZN(new_n202));
  NAND2_X1  g001(.A1(G229gat), .A2(G233gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT97), .ZN(new_n206));
  INV_X1    g005(.A(G1gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT16), .ZN(new_n208));
  INV_X1    g007(.A(G22gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G15gat), .ZN(new_n210));
  INV_X1    g009(.A(G15gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G22gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT96), .ZN(new_n213));
  AND3_X1   g012(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n213), .B1(new_n210), .B2(new_n212), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n208), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n210), .A2(new_n212), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT96), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(new_n207), .ZN(new_n220));
  INV_X1    g019(.A(G8gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n216), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n221), .B1(new_n216), .B2(new_n220), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n206), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G29gat), .ZN(new_n226));
  INV_X1    g025(.A(G36gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT14), .ZN(new_n228));
  NAND2_X1  g027(.A1(G29gat), .A2(G36gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT91), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT14), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G29gat), .B2(G36gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(KEYINPUT91), .A2(G29gat), .A3(G36gat), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n228), .A2(new_n231), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G50gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G43gat), .ZN(new_n237));
  INV_X1    g036(.A(G43gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G50gat), .ZN(new_n239));
  AND3_X1   g038(.A1(new_n237), .A2(new_n239), .A3(KEYINPUT15), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n235), .A2(new_n240), .A3(KEYINPUT92), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n235), .A2(new_n240), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT92), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n231), .A2(new_n234), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n245), .B1(new_n240), .B2(KEYINPUT93), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT15), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT94), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(new_n236), .B2(G43gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n237), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n239), .A2(new_n248), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n247), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n228), .A2(new_n233), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT95), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT95), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n228), .A2(new_n233), .A3(new_n256), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n255), .B(new_n257), .C1(new_n240), .C2(KEYINPUT93), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n241), .B(new_n244), .C1(new_n253), .C2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n216), .A2(new_n220), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G8gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(new_n222), .A3(KEYINPUT97), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n225), .A2(new_n260), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n260), .B1(new_n225), .B2(new_n263), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n205), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n262), .A2(new_n222), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n259), .A2(KEYINPUT17), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT17), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n244), .A2(new_n241), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n255), .A2(new_n257), .ZN(new_n273));
  OR2_X1    g072(.A1(new_n240), .A2(KEYINPUT93), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n273), .A2(new_n274), .A3(new_n246), .A4(new_n252), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n271), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n269), .B1(new_n270), .B2(new_n276), .ZN(new_n277));
  NOR3_X1   g076(.A1(new_n223), .A2(new_n224), .A3(new_n206), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT97), .B1(new_n262), .B2(new_n222), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n259), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n277), .A2(new_n280), .A3(KEYINPUT18), .A4(new_n203), .ZN(new_n281));
  XNOR2_X1  g080(.A(G113gat), .B(G141gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(G197gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT11), .B(G169gat), .ZN(new_n284));
  XOR2_X1   g083(.A(new_n283), .B(new_n284), .Z(new_n285));
  XNOR2_X1  g084(.A(new_n285), .B(KEYINPUT12), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n267), .A2(new_n281), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n277), .A2(new_n280), .A3(new_n203), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT18), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT99), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n288), .A2(KEYINPUT99), .A3(new_n289), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n287), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n290), .A2(new_n267), .A3(new_n281), .ZN(new_n295));
  INV_X1    g094(.A(new_n286), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT100), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  AND2_X1   g099(.A1(G127gat), .A2(G134gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(G127gat), .A2(G134gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT1), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n305), .B1(G113gat), .B2(G120gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(G113gat), .A2(G120gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n303), .B(new_n304), .C1(new_n306), .C2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n306), .A2(new_n308), .ZN(new_n310));
  INV_X1    g109(.A(G127gat), .ZN(new_n311));
  INV_X1    g110(.A(G134gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G127gat), .A2(G134gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT70), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT72), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(new_n301), .B2(new_n302), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n313), .A2(KEYINPUT72), .A3(new_n314), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(KEYINPUT71), .A2(G113gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(KEYINPUT71), .A2(G113gat), .ZN(new_n322));
  OAI21_X1  g121(.A(G120gat), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G113gat), .ZN(new_n324));
  INV_X1    g123(.A(G120gat), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT1), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n309), .B(new_n316), .C1(new_n320), .C2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT77), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT71), .B(G113gat), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n306), .B1(new_n331), .B2(G120gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n318), .A2(new_n319), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n334), .A2(KEYINPUT77), .A3(new_n309), .A4(new_n316), .ZN(new_n335));
  NAND2_X1  g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT2), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT76), .ZN(new_n338));
  XNOR2_X1  g137(.A(G155gat), .B(G162gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(G141gat), .B(G148gat), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n336), .A2(KEYINPUT2), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n338), .B(new_n339), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(G141gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G148gat), .ZN(new_n344));
  INV_X1    g143(.A(G148gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G141gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AND2_X1   g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n337), .B(new_n347), .C1(new_n350), .C2(KEYINPUT76), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n342), .A2(new_n351), .A3(KEYINPUT3), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n342), .A2(new_n351), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n330), .A2(new_n335), .A3(new_n352), .A4(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT5), .ZN(new_n357));
  NAND2_X1  g156(.A1(G225gat), .A2(G233gat), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n358), .B(KEYINPUT78), .Z(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n356), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n342), .A2(new_n351), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT4), .B1(new_n328), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT81), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT80), .ZN(new_n365));
  INV_X1    g164(.A(new_n328), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(new_n367), .A3(new_n353), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n353), .A2(new_n309), .A3(new_n334), .A4(new_n316), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT4), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n364), .A2(new_n365), .A3(new_n368), .A4(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n365), .B1(new_n369), .B2(KEYINPUT4), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT4), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n370), .B1(new_n369), .B2(KEYINPUT4), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n372), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT82), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n361), .A2(new_n376), .A3(new_n372), .A4(KEYINPUT82), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n368), .A2(new_n363), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(new_n356), .A3(new_n360), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n330), .A2(new_n335), .A3(new_n362), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n369), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n359), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n383), .A2(new_n386), .A3(KEYINPUT5), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n381), .A2(new_n388), .ZN(new_n389));
  XOR2_X1   g188(.A(G1gat), .B(G29gat), .Z(new_n390));
  XNOR2_X1  g189(.A(G57gat), .B(G85gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n389), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n387), .B1(new_n379), .B2(new_n380), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT6), .B1(new_n397), .B2(new_n394), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n389), .A2(KEYINPUT6), .A3(new_n395), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT35), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT24), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n404), .A2(G183gat), .A3(G190gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(G183gat), .B(G190gat), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n405), .B1(new_n406), .B2(new_n404), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT67), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(G169gat), .A2(G176gat), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT23), .B1(new_n410), .B2(KEYINPUT66), .ZN(new_n411));
  NAND2_X1  g210(.A1(G169gat), .A2(G176gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT25), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n410), .A2(KEYINPUT66), .A3(KEYINPUT23), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n409), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT65), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n407), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n413), .A2(new_n415), .ZN(new_n420));
  OAI211_X1 g219(.A(KEYINPUT65), .B(new_n405), .C1(new_n406), .C2(new_n404), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n414), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n417), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT69), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT27), .B(G183gat), .ZN(new_n426));
  INV_X1    g225(.A(G190gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT28), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n429), .A2(KEYINPUT68), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G183gat), .A2(G190gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT26), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n410), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n435), .B1(new_n410), .B2(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n438));
  OAI21_X1  g237(.A(new_n437), .B1(new_n428), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n425), .B1(new_n433), .B2(new_n439), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n428), .A2(new_n438), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n428), .A2(new_n430), .B1(G183gat), .B2(G190gat), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT69), .A4(new_n437), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n424), .A2(new_n328), .A3(new_n440), .A4(new_n443), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n409), .A2(new_n416), .B1(new_n422), .B2(new_n414), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n440), .A2(new_n443), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n366), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(G227gat), .A2(G233gat), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n448), .B(KEYINPUT64), .Z(new_n449));
  NAND3_X1  g248(.A1(new_n444), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  XOR2_X1   g249(.A(G71gat), .B(G99gat), .Z(new_n451));
  XNOR2_X1  g250(.A(G15gat), .B(G43gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT33), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n450), .A2(KEYINPUT32), .A3(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(KEYINPUT73), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n450), .A2(KEYINPUT32), .ZN(new_n457));
  INV_X1    g256(.A(new_n450), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n457), .B(new_n453), .C1(new_n458), .C2(KEYINPUT33), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n447), .ZN(new_n461));
  INV_X1    g260(.A(new_n449), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT34), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n464), .B1(new_n462), .B2(KEYINPUT74), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n461), .B(new_n462), .C1(KEYINPUT74), .C2(new_n464), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n460), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n468), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n456), .A2(new_n459), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(G197gat), .B(G204gat), .ZN(new_n473));
  INV_X1    g272(.A(G211gat), .ZN(new_n474));
  INV_X1    g273(.A(G218gat), .ZN(new_n475));
  OAI22_X1  g274(.A1(new_n474), .A2(new_n475), .B1(KEYINPUT75), .B2(KEYINPUT22), .ZN(new_n476));
  AND2_X1   g275(.A1(KEYINPUT75), .A2(KEYINPUT22), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(G211gat), .B(G218gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT29), .B1(new_n353), .B2(new_n354), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n483), .B2(KEYINPUT86), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(KEYINPUT86), .B2(new_n483), .ZN(new_n485));
  INV_X1    g284(.A(G228gat), .ZN(new_n486));
  INV_X1    g285(.A(G233gat), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n354), .B1(new_n480), .B2(KEYINPUT29), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n489), .A2(KEYINPUT85), .A3(new_n362), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n362), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT85), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n485), .A2(new_n488), .A3(new_n490), .A4(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n491), .B1(new_n481), .B2(new_n482), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n495), .B1(new_n486), .B2(new_n487), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n209), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n494), .A2(new_n496), .A3(new_n209), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G78gat), .B(G106gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT31), .B(G50gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT87), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n503), .B1(new_n497), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n498), .A2(new_n504), .A3(new_n499), .A4(new_n503), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G226gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n510), .A2(new_n487), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(KEYINPUT29), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n441), .A2(new_n442), .A3(new_n437), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n513), .B1(new_n424), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n511), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n445), .A2(new_n446), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n481), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n424), .A2(new_n511), .A3(new_n514), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n512), .B1(new_n445), .B2(new_n446), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n520), .A3(new_n480), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G8gat), .B(G36gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(G64gat), .B(G92gat), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n523), .B(new_n524), .Z(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n518), .A2(new_n521), .A3(new_n525), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(KEYINPUT30), .A3(new_n528), .ZN(new_n529));
  OR3_X1    g328(.A1(new_n522), .A2(KEYINPUT30), .A3(new_n526), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NOR4_X1   g330(.A1(new_n403), .A2(new_n472), .A3(new_n509), .A4(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT83), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n389), .A2(new_n533), .A3(new_n395), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT83), .B1(new_n397), .B2(new_n394), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n398), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(new_n400), .ZN(new_n537));
  INV_X1    g336(.A(new_n531), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT84), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT84), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n537), .A2(new_n541), .A3(new_n538), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n472), .A2(new_n509), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n532), .B1(new_n544), .B2(KEYINPUT35), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n541), .B1(new_n537), .B2(new_n538), .ZN(new_n547));
  AOI211_X1 g346(.A(KEYINPUT84), .B(new_n531), .C1(new_n536), .C2(new_n400), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n509), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT36), .ZN(new_n550));
  INV_X1    g349(.A(new_n471), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n470), .B1(new_n456), .B2(new_n459), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n469), .A2(KEYINPUT36), .A3(new_n471), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n384), .A2(new_n360), .A3(new_n369), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT39), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT89), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n376), .A2(new_n372), .A3(new_n356), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n359), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(KEYINPUT88), .B(KEYINPUT39), .Z(new_n562));
  NAND3_X1  g361(.A1(new_n559), .A2(new_n359), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n394), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT40), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n561), .A2(KEYINPUT40), .A3(new_n394), .A4(new_n563), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n531), .A2(new_n566), .A3(new_n396), .A4(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT37), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n519), .A2(new_n520), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT90), .B1(new_n570), .B2(new_n481), .ZN(new_n571));
  NOR3_X1   g370(.A1(new_n515), .A2(new_n517), .A3(new_n481), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(KEYINPUT90), .A3(new_n481), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n569), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT38), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n576), .B(new_n526), .C1(new_n522), .C2(KEYINPUT37), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n526), .B1(new_n522), .B2(KEYINPUT37), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n578), .B1(KEYINPUT37), .B2(new_n522), .ZN(new_n579));
  OAI221_X1 g378(.A(new_n528), .B1(new_n575), .B2(new_n577), .C1(new_n579), .C2(new_n576), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n508), .B(new_n568), .C1(new_n580), .C2(new_n401), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n549), .A2(new_n555), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n300), .B1(new_n546), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n537), .ZN(new_n584));
  OR2_X1    g383(.A1(KEYINPUT102), .A2(G57gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(KEYINPUT102), .A2(G57gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(G64gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G71gat), .A2(G78gat), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT9), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n585), .A2(G64gat), .A3(new_n586), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n589), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(G71gat), .ZN(new_n595));
  INV_X1    g394(.A(G78gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT101), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n597), .B1(new_n598), .B2(new_n590), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n599), .B1(new_n598), .B2(new_n590), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n590), .B1(new_n597), .B2(new_n591), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT103), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(G57gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(G64gat), .ZN(new_n604));
  AOI22_X1  g403(.A1(new_n594), .A2(new_n600), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT104), .B(KEYINPUT21), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n607), .B(new_n608), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(new_n311), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n605), .A2(KEYINPUT21), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n225), .A2(new_n263), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n610), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT105), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G155gat), .ZN(new_n616));
  XOR2_X1   g415(.A(G183gat), .B(G211gat), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n613), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G99gat), .A2(G106gat), .ZN(new_n620));
  INV_X1    g419(.A(G85gat), .ZN(new_n621));
  INV_X1    g420(.A(G92gat), .ZN(new_n622));
  AOI22_X1  g421(.A1(KEYINPUT8), .A2(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND4_X1  g422(.A1(KEYINPUT106), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n624));
  NAND3_X1  g423(.A1(KEYINPUT106), .A2(G85gat), .A3(G92gat), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT7), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n623), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT108), .ZN(new_n629));
  XNOR2_X1  g428(.A(G99gat), .B(G106gat), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n628), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n629), .B1(new_n628), .B2(new_n631), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n623), .A2(new_n630), .A3(new_n624), .A4(new_n627), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT107), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n639), .B1(new_n270), .B2(new_n276), .ZN(new_n640));
  XOR2_X1   g439(.A(G190gat), .B(G218gat), .Z(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n628), .A2(new_n631), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(KEYINPUT108), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n632), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n636), .B(KEYINPUT107), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n259), .ZN(new_n648));
  NAND2_X1  g447(.A1(G232gat), .A2(G233gat), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT41), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n640), .A2(new_n642), .A3(new_n648), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n259), .A2(KEYINPUT17), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n272), .A2(new_n275), .A3(new_n271), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n647), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n651), .B1(new_n260), .B2(new_n639), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n641), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n650), .A2(KEYINPUT41), .ZN(new_n658));
  XNOR2_X1  g457(.A(G134gat), .B(G162gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n652), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n660), .B1(new_n652), .B2(new_n657), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n619), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT111), .ZN(new_n666));
  XNOR2_X1  g465(.A(G120gat), .B(G148gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(G176gat), .B(G204gat), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n667), .B(new_n668), .Z(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(G230gat), .A2(G233gat), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(KEYINPUT109), .Z(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n605), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(new_n645), .B2(new_n646), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n638), .A2(new_n605), .A3(new_n643), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n673), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n670), .B1(new_n677), .B2(KEYINPUT110), .ZN(new_n678));
  INV_X1    g477(.A(new_n676), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n605), .B1(new_n635), .B2(new_n638), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n672), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT110), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT10), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n675), .A2(new_n685), .A3(new_n676), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n635), .A2(new_n605), .A3(new_n638), .A4(KEYINPUT10), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n672), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n666), .B1(new_n684), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n688), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n690), .A2(new_n678), .A3(KEYINPUT111), .A4(new_n683), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n670), .B1(new_n688), .B2(new_n677), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n665), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n583), .A2(new_n584), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g496(.A1(new_n583), .A2(new_n695), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n698), .A2(new_n538), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT16), .B(G8gat), .Z(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(KEYINPUT42), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(G8gat), .B1(new_n698), .B2(new_n538), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT113), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n699), .A2(new_n700), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n706), .A2(KEYINPUT112), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(KEYINPUT112), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n701), .B(new_n703), .C1(new_n707), .C2(new_n708), .ZN(G1325gat));
  OAI21_X1  g508(.A(G15gat), .B1(new_n698), .B2(new_n555), .ZN(new_n710));
  INV_X1    g509(.A(new_n472), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n211), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n698), .B2(new_n712), .ZN(G1326gat));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n508), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT43), .B(G22gat), .Z(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  XNOR2_X1  g515(.A(new_n298), .B(KEYINPUT100), .ZN(new_n717));
  INV_X1    g516(.A(new_n619), .ZN(new_n718));
  INV_X1    g517(.A(new_n694), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n664), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n580), .A2(new_n401), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n568), .A2(new_n508), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n555), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n540), .A2(new_n542), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n725), .B2(new_n509), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n717), .B(new_n721), .C1(new_n545), .C2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n728), .A2(new_n226), .A3(new_n584), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT45), .ZN(new_n730));
  INV_X1    g529(.A(new_n298), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n720), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT114), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(new_n545), .B2(new_n726), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n547), .A2(new_n548), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n402), .B1(new_n736), .B2(new_n543), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n582), .B(KEYINPUT114), .C1(new_n737), .C2(new_n532), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n664), .A2(KEYINPUT44), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n735), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n663), .B1(new_n545), .B2(new_n726), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT44), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n733), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(new_n584), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n730), .B1(new_n744), .B2(new_n226), .ZN(G1328gat));
  NOR3_X1   g544(.A1(new_n727), .A2(G36gat), .A3(new_n538), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT46), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n743), .A2(new_n531), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n227), .ZN(G1329gat));
  INV_X1    g548(.A(KEYINPUT47), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n472), .A2(G43gat), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n728), .B2(new_n751), .ZN(new_n752));
  AOI211_X1 g551(.A(new_n555), .B(new_n733), .C1(new_n740), .C2(new_n742), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n753), .B2(new_n238), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n583), .A2(KEYINPUT116), .A3(new_n721), .A4(new_n751), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT116), .ZN(new_n756));
  INV_X1    g555(.A(new_n751), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n727), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n740), .A2(new_n742), .ZN(new_n760));
  INV_X1    g559(.A(new_n555), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n760), .A2(new_n761), .A3(new_n732), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n759), .B1(new_n762), .B2(G43gat), .ZN(new_n763));
  XOR2_X1   g562(.A(KEYINPUT115), .B(KEYINPUT47), .Z(new_n764));
  OAI21_X1  g563(.A(new_n754), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT117), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n754), .B(KEYINPUT117), .C1(new_n763), .C2(new_n764), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(G1330gat));
  NOR3_X1   g568(.A1(new_n727), .A2(G50gat), .A3(new_n508), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n743), .A2(new_n509), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n772), .B2(new_n236), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT48), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1331gat));
  AND2_X1   g574(.A1(new_n735), .A2(new_n738), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n665), .A2(new_n298), .A3(new_n719), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n537), .ZN(new_n779));
  XOR2_X1   g578(.A(new_n779), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g579(.A1(new_n778), .A2(new_n538), .ZN(new_n781));
  NOR2_X1   g580(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n782));
  AND2_X1   g581(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n781), .B2(new_n782), .ZN(G1333gat));
  OAI21_X1  g584(.A(G71gat), .B1(new_n778), .B2(new_n555), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n711), .A2(new_n595), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n778), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(G1334gat));
  NOR2_X1   g589(.A1(new_n778), .A2(new_n508), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(new_n596), .ZN(G1335gat));
  NOR2_X1   g591(.A1(new_n619), .A2(new_n298), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT118), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n760), .A2(new_n694), .A3(new_n794), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n795), .A2(new_n584), .ZN(new_n796));
  INV_X1    g595(.A(new_n741), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n794), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n797), .A2(KEYINPUT51), .A3(new_n794), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n694), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n584), .A2(new_n621), .ZN(new_n804));
  OAI22_X1  g603(.A1(new_n796), .A2(new_n621), .B1(new_n803), .B2(new_n804), .ZN(G1336gat));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  AND4_X1   g605(.A1(new_n531), .A2(new_n760), .A3(new_n694), .A4(new_n794), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n531), .A2(new_n622), .ZN(new_n808));
  OAI221_X1 g607(.A(new_n806), .B1(new_n807), .B2(new_n622), .C1(new_n803), .C2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n807), .A2(new_n622), .ZN(new_n810));
  AOI211_X1 g609(.A(new_n719), .B(new_n808), .C1(new_n800), .C2(new_n801), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT52), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n809), .A2(new_n812), .ZN(G1337gat));
  AND2_X1   g612(.A1(new_n795), .A2(new_n761), .ZN(new_n814));
  INV_X1    g613(.A(G99gat), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n711), .A2(new_n815), .ZN(new_n816));
  OAI22_X1  g615(.A1(new_n814), .A2(new_n815), .B1(new_n803), .B2(new_n816), .ZN(G1338gat));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818));
  AND4_X1   g617(.A1(new_n509), .A2(new_n760), .A3(new_n694), .A4(new_n794), .ZN(new_n819));
  INV_X1    g618(.A(G106gat), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n509), .A2(new_n820), .ZN(new_n821));
  OAI221_X1 g620(.A(new_n818), .B1(new_n819), .B2(new_n820), .C1(new_n803), .C2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n819), .A2(new_n820), .ZN(new_n823));
  AOI211_X1 g622(.A(new_n719), .B(new_n821), .C1(new_n800), .C2(new_n801), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT53), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n822), .A2(new_n825), .ZN(G1339gat));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n686), .A2(new_n672), .A3(new_n687), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n828), .A2(new_n688), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n686), .A2(new_n687), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n829), .A3(new_n673), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n670), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n827), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n669), .B1(new_n688), .B2(new_n829), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n690), .A2(KEYINPUT54), .ZN(new_n836));
  OAI211_X1 g635(.A(KEYINPUT55), .B(new_n835), .C1(new_n836), .C2(new_n828), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n692), .A2(new_n834), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n280), .A2(new_n264), .A3(new_n204), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n203), .B1(new_n277), .B2(new_n280), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n285), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n277), .A2(new_n280), .ZN(new_n845));
  INV_X1    g644(.A(new_n203), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n839), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(KEYINPUT119), .A3(new_n285), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n288), .A2(KEYINPUT99), .A3(new_n289), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT99), .B1(new_n288), .B2(new_n289), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI22_X1  g651(.A1(new_n844), .A2(new_n849), .B1(new_n852), .B2(new_n287), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n838), .A2(new_n853), .A3(new_n854), .A4(new_n663), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT119), .B1(new_n848), .B2(new_n285), .ZN(new_n856));
  INV_X1    g655(.A(new_n285), .ZN(new_n857));
  AOI211_X1 g656(.A(new_n843), .B(new_n857), .C1(new_n847), .C2(new_n839), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n294), .B(new_n663), .C1(new_n856), .C2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n692), .A2(new_n834), .A3(new_n837), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT120), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n298), .A2(new_n692), .A3(new_n834), .A4(new_n837), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n844), .A2(new_n849), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n694), .A2(new_n294), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n663), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n718), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n619), .A2(new_n731), .A3(new_n664), .A4(new_n719), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n868), .B1(new_n867), .B2(new_n869), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n537), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n538), .A3(new_n543), .ZN(new_n875));
  OAI21_X1  g674(.A(G113gat), .B1(new_n875), .B2(new_n300), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n731), .A2(new_n331), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n875), .B2(new_n877), .ZN(G1340gat));
  NOR2_X1   g677(.A1(new_n875), .A2(new_n719), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(new_n325), .ZN(G1341gat));
  NOR2_X1   g679(.A1(new_n875), .A2(new_n718), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(new_n311), .ZN(G1342gat));
  NOR3_X1   g681(.A1(new_n531), .A2(G134gat), .A3(new_n664), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n874), .A2(new_n543), .A3(new_n883), .ZN(new_n884));
  XOR2_X1   g683(.A(new_n884), .B(KEYINPUT56), .Z(new_n885));
  OAI21_X1  g684(.A(G134gat), .B1(new_n875), .B2(new_n664), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1343gat));
  AND2_X1   g686(.A1(new_n509), .A2(KEYINPUT57), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n865), .B1(new_n300), .B2(new_n860), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n664), .ZN(new_n890));
  INV_X1    g689(.A(new_n862), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n619), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n869), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n888), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n870), .A2(new_n871), .A3(new_n508), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n895), .B2(KEYINPUT57), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n555), .A2(new_n584), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n538), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(G141gat), .B1(new_n901), .B2(new_n300), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT58), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n300), .A2(G141gat), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n895), .A2(new_n538), .A3(new_n898), .A4(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n896), .A2(new_n298), .A3(new_n900), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n907), .A2(new_n908), .A3(G141gat), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT58), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n905), .A2(KEYINPUT122), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n911), .B1(new_n907), .B2(G141gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n906), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n906), .B(KEYINPUT123), .C1(new_n910), .C2(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1344gat));
  INV_X1    g716(.A(KEYINPUT125), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n899), .A2(new_n719), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n895), .A2(new_n345), .A3(new_n919), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT124), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n901), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n694), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n345), .A2(KEYINPUT59), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT59), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n872), .A2(new_n888), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n717), .A2(new_n838), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n663), .B1(new_n929), .B2(new_n865), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n859), .A2(new_n860), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n718), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n695), .A2(new_n300), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT57), .B1(new_n934), .B2(new_n509), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n919), .B1(new_n928), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n927), .B1(new_n936), .B2(G148gat), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n918), .B(new_n922), .C1(new_n926), .C2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n937), .B1(new_n924), .B2(new_n925), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT125), .B1(new_n939), .B2(new_n921), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1345gat));
  INV_X1    g740(.A(G155gat), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n901), .A2(new_n942), .A3(new_n718), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n895), .A2(new_n898), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n538), .A3(new_n619), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n943), .B1(new_n942), .B2(new_n945), .ZN(G1346gat));
  NAND2_X1  g745(.A1(new_n923), .A2(new_n663), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n531), .A2(G162gat), .A3(new_n664), .ZN(new_n948));
  AOI22_X1  g747(.A1(new_n947), .A2(G162gat), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT126), .ZN(G1347gat));
  NAND2_X1  g749(.A1(new_n537), .A2(new_n531), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n951), .A2(new_n472), .A3(new_n509), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n872), .A2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n954), .A2(G169gat), .A3(new_n717), .ZN(new_n955));
  AOI21_X1  g754(.A(G169gat), .B1(new_n954), .B2(new_n298), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n955), .A2(new_n956), .ZN(G1348gat));
  NAND2_X1  g756(.A1(new_n954), .A2(new_n694), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g758(.A1(new_n954), .A2(new_n619), .ZN(new_n960));
  INV_X1    g759(.A(G183gat), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n962), .B1(new_n426), .B2(new_n960), .ZN(new_n963));
  XOR2_X1   g762(.A(new_n963), .B(KEYINPUT60), .Z(G1350gat));
  OAI22_X1  g763(.A1(new_n953), .A2(new_n664), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n965));
  NAND2_X1  g764(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n965), .B(new_n966), .ZN(G1351gat));
  NOR2_X1   g766(.A1(new_n928), .A2(new_n935), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n968), .A2(new_n761), .A3(new_n951), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(G197gat), .B1(new_n970), .B2(new_n300), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n761), .A2(new_n508), .A3(new_n951), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n872), .A2(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n974), .A2(G197gat), .A3(new_n731), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT127), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n971), .A2(new_n976), .ZN(G1352gat));
  OAI21_X1  g776(.A(G204gat), .B1(new_n970), .B2(new_n719), .ZN(new_n978));
  NOR3_X1   g777(.A1(new_n974), .A2(G204gat), .A3(new_n719), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(KEYINPUT62), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(G1353gat));
  NAND3_X1  g780(.A1(new_n973), .A2(new_n474), .A3(new_n619), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n969), .A2(new_n619), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n983), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n984));
  AOI21_X1  g783(.A(KEYINPUT63), .B1(new_n983), .B2(G211gat), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(G1354gat));
  OAI21_X1  g785(.A(G218gat), .B1(new_n970), .B2(new_n664), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n973), .A2(new_n475), .A3(new_n663), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(G1355gat));
endmodule


