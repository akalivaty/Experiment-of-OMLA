//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n809, new_n810, new_n812, new_n813, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G141gat), .B(G148gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  OR2_X1    g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(KEYINPUT2), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n205), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n207), .B(new_n206), .C1(new_n204), .C2(KEYINPUT2), .ZN(new_n211));
  AND2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT4), .ZN(new_n213));
  INV_X1    g012(.A(G127gat), .ZN(new_n214));
  NOR3_X1   g013(.A1(new_n214), .A2(KEYINPUT67), .A3(G134gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(G127gat), .B(G134gat), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(KEYINPUT67), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT1), .ZN(new_n218));
  INV_X1    g017(.A(G120gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(G113gat), .ZN(new_n220));
  INV_X1    g019(.A(G113gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(G120gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n218), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT68), .B1(new_n219), .B2(G113gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(new_n221), .A3(G120gat), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n224), .B(new_n226), .C1(new_n221), .C2(G120gat), .ZN(new_n227));
  INV_X1    g026(.A(G134gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G127gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n214), .A2(G134gat), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n229), .A2(new_n230), .A3(new_n218), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n217), .A2(new_n223), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n212), .A2(new_n213), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n215), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n229), .A2(new_n230), .A3(KEYINPUT67), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n223), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n227), .A2(new_n231), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n210), .A2(new_n211), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT4), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n203), .B1(new_n233), .B2(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n238), .A2(KEYINPUT76), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT76), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n232), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n239), .A2(KEYINPUT3), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n210), .A2(new_n211), .A3(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n243), .A2(new_n245), .A3(new_n246), .A4(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(KEYINPUT77), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT77), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n236), .A2(new_n237), .A3(new_n244), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n244), .B1(new_n236), .B2(new_n237), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n210), .A2(new_n211), .A3(new_n247), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n247), .B1(new_n210), .B2(new_n211), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n251), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n241), .B(new_n242), .C1(new_n250), .C2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n233), .A2(new_n240), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n202), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n249), .A2(KEYINPUT77), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n254), .A2(new_n251), .A3(new_n257), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n242), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n238), .A2(new_n239), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n266), .B1(new_n254), .B2(new_n239), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n265), .B1(new_n267), .B2(new_n202), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n259), .B1(new_n264), .B2(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(KEYINPUT79), .B(KEYINPUT0), .Z(new_n270));
  XNOR2_X1  g069(.A(G1gat), .B(G29gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G57gat), .B(G85gat), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n272), .B(new_n273), .Z(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n269), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n259), .B(new_n274), .C1(new_n264), .C2(new_n268), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n278), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n269), .A2(new_n275), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G15gat), .B(G22gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT86), .ZN(new_n284));
  INV_X1    g083(.A(G1gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(G8gat), .B1(new_n286), .B2(KEYINPUT87), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT86), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n283), .B(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT16), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n289), .B1(new_n290), .B2(G1gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n286), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n291), .B(new_n286), .C1(KEYINPUT87), .C2(G8gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G71gat), .B(G78gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(KEYINPUT92), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(G57gat), .B(G64gat), .ZN(new_n299));
  NOR3_X1   g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(KEYINPUT92), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g101(.A(KEYINPUT92), .B(new_n296), .C1(new_n299), .C2(new_n298), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT21), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n295), .A2(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(KEYINPUT93), .B(KEYINPUT94), .Z(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n309));
  NAND2_X1  g108(.A1(G231gat), .A2(G233gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n308), .B(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n304), .A2(KEYINPUT21), .ZN(new_n313));
  XOR2_X1   g112(.A(G127gat), .B(G155gat), .Z(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(G183gat), .B(G211gat), .Z(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(new_n317), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G29gat), .ZN(new_n322));
  INV_X1    g121(.A(G36gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT14), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT14), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n325), .B1(G29gat), .B2(G36gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT85), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n322), .A2(new_n323), .ZN(new_n329));
  XNOR2_X1  g128(.A(G43gat), .B(G50gat), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n329), .B1(new_n330), .B2(KEYINPUT15), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(KEYINPUT15), .B2(new_n330), .ZN(new_n332));
  OR2_X1    g131(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g132(.A(KEYINPUT15), .B(new_n330), .C1(new_n327), .C2(new_n329), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT17), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n333), .A2(KEYINPUT17), .A3(new_n334), .ZN(new_n338));
  NAND2_X1  g137(.A1(G85gat), .A2(G92gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT7), .ZN(new_n340));
  NAND2_X1  g139(.A1(G99gat), .A2(G106gat), .ZN(new_n341));
  INV_X1    g140(.A(G85gat), .ZN(new_n342));
  INV_X1    g141(.A(G92gat), .ZN(new_n343));
  AOI22_X1  g142(.A1(KEYINPUT8), .A2(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(G99gat), .B(G106gat), .Z(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n345), .B(new_n347), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n348), .A2(KEYINPUT95), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(KEYINPUT95), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n337), .A2(new_n338), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  AND2_X1   g150(.A1(G232gat), .A2(G233gat), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n335), .A2(new_n348), .B1(KEYINPUT41), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G134gat), .B(G162gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n354), .B(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n352), .A2(KEYINPUT41), .ZN(new_n358));
  XNOR2_X1  g157(.A(G190gat), .B(G218gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n357), .B(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n321), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G230gat), .ZN(new_n363));
  INV_X1    g162(.A(G233gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT96), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n346), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n304), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n348), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n302), .A2(new_n303), .B1(new_n366), .B2(new_n346), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n348), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n304), .A2(KEYINPUT10), .A3(new_n348), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n365), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n372), .B(new_n369), .ZN(new_n377));
  INV_X1    g176(.A(new_n365), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT98), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G176gat), .B(G204gat), .ZN(new_n381));
  INV_X1    g180(.A(G148gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT97), .B(G120gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  OR2_X1    g185(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n380), .A2(new_n386), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n362), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT72), .ZN(new_n394));
  XOR2_X1   g193(.A(G211gat), .B(G218gat), .Z(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT73), .ZN(new_n396));
  XNOR2_X1  g195(.A(G197gat), .B(G204gat), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n394), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT73), .ZN(new_n399));
  INV_X1    g198(.A(new_n395), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT29), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n399), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n403), .A2(new_n394), .A3(new_n396), .A4(new_n397), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n401), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n212), .B1(new_n405), .B2(new_n247), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(G50gat), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n401), .A2(new_n404), .B1(new_n402), .B2(new_n248), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n407), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(G50gat), .B1(new_n406), .B2(new_n409), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n409), .A2(KEYINPUT81), .ZN(new_n414));
  INV_X1    g213(.A(G228gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n415), .A2(new_n364), .ZN(new_n416));
  OAI21_X1  g215(.A(G22gat), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G22gat), .ZN(new_n418));
  OAI221_X1 g217(.A(new_n418), .B1(new_n415), .B2(new_n364), .C1(new_n409), .C2(KEYINPUT81), .ZN(new_n419));
  XNOR2_X1  g218(.A(G78gat), .B(G106gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT31), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n417), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n422), .B1(new_n417), .B2(new_n419), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n413), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n417), .A2(new_n419), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n421), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n428), .A2(new_n412), .A3(new_n411), .A4(new_n423), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n401), .A2(new_n404), .ZN(new_n431));
  NAND2_X1  g230(.A1(G169gat), .A2(G176gat), .ZN(new_n432));
  NOR2_X1   g231(.A1(G169gat), .A2(G176gat), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT26), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NOR3_X1   g234(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(G183gat), .A2(G190gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  XOR2_X1   g238(.A(KEYINPUT27), .B(G183gat), .Z(new_n440));
  INV_X1    g239(.A(KEYINPUT28), .ZN(new_n441));
  OR3_X1    g240(.A1(new_n440), .A2(new_n441), .A3(G190gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n443));
  AOI21_X1  g242(.A(G190gat), .B1(new_n443), .B2(KEYINPUT27), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n444), .B1(KEYINPUT27), .B2(new_n443), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n441), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n439), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G169gat), .ZN(new_n448));
  INV_X1    g247(.A(G176gat), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT23), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT64), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n433), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT23), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n454), .B1(G169gat), .B2(G176gat), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n452), .A2(new_n453), .A3(new_n432), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT65), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n455), .A2(new_n432), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT65), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n458), .A2(new_n459), .A3(new_n453), .A4(new_n452), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT24), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(G183gat), .A3(G190gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(G183gat), .B(G190gat), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n462), .B1(new_n463), .B2(new_n461), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n457), .A2(new_n460), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT25), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n458), .A2(KEYINPUT25), .A3(new_n450), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n469), .A2(new_n464), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n447), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(G226gat), .A2(G233gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n473), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n442), .A2(new_n446), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n476), .A2(new_n438), .A3(new_n437), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n464), .B1(new_n456), .B2(KEYINPUT65), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT25), .B1(new_n478), .B2(new_n460), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n477), .B1(new_n479), .B2(new_n470), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n475), .B1(new_n480), .B2(new_n402), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n431), .B1(new_n474), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n473), .B1(new_n472), .B2(KEYINPUT29), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n431), .B1(new_n480), .B2(new_n475), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G8gat), .B(G36gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(G92gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT74), .B(G64gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n482), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(KEYINPUT75), .B(KEYINPUT30), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n482), .A2(new_n485), .A3(KEYINPUT30), .A4(new_n490), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n482), .A2(new_n485), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n489), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n260), .B1(new_n250), .B2(new_n258), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT39), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n499), .A3(new_n203), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n499), .B1(new_n267), .B2(new_n202), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n233), .A2(new_n240), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n502), .B1(new_n262), .B2(new_n263), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n501), .B1(new_n503), .B2(new_n202), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n500), .A2(new_n504), .A3(KEYINPUT40), .A4(new_n274), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n500), .A2(new_n504), .A3(new_n274), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT40), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n506), .A2(new_n507), .B1(new_n275), .B2(new_n269), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n497), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT37), .ZN(new_n510));
  INV_X1    g309(.A(new_n431), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n511), .B1(new_n472), .B2(new_n473), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n510), .B1(new_n512), .B2(new_n481), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n480), .A2(new_n475), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n511), .B1(new_n483), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n489), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n510), .B1(new_n482), .B2(new_n485), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT38), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n518), .A2(new_n281), .A3(new_n279), .A4(new_n491), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT82), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n490), .A2(KEYINPUT38), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(new_n513), .B2(new_n515), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n520), .B1(new_n522), .B2(new_n517), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n495), .A2(KEYINPUT37), .ZN(new_n524));
  INV_X1    g323(.A(new_n521), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT37), .B1(new_n483), .B2(new_n484), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n525), .B1(new_n526), .B2(new_n482), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n524), .A2(KEYINPUT82), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n430), .B(new_n509), .C1(new_n519), .C2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n470), .B1(new_n466), .B2(new_n467), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n232), .B1(new_n531), .B2(new_n447), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n477), .B(new_n238), .C1(new_n479), .C2(new_n470), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n532), .A2(G227gat), .A3(G233gat), .A4(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT32), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT33), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G15gat), .B(G43gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(G71gat), .B(G99gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n535), .B1(new_n541), .B2(KEYINPUT33), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n537), .A2(new_n541), .B1(new_n534), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n532), .A2(new_n533), .ZN(new_n544));
  NAND2_X1  g343(.A1(G227gat), .A2(G233gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT34), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n546), .A2(KEYINPUT69), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(KEYINPUT69), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n544), .A2(new_n545), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n532), .A2(new_n533), .B1(G227gat), .B2(G233gat), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n549), .B1(new_n550), .B2(new_n548), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n543), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n544), .A2(new_n545), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(KEYINPUT69), .A3(new_n546), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n534), .A2(new_n542), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n540), .B1(new_n534), .B2(new_n536), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n549), .B(new_n554), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT70), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT71), .B1(new_n552), .B2(new_n557), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n560), .B(KEYINPUT36), .C1(new_n559), .C2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT36), .ZN(new_n563));
  INV_X1    g362(.A(new_n558), .ZN(new_n564));
  OAI211_X1 g363(.A(KEYINPUT70), .B(new_n563), .C1(new_n564), .C2(KEYINPUT71), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n282), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n426), .A2(new_n429), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n530), .A2(new_n562), .A3(new_n565), .A4(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n568), .A2(new_n558), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT35), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n571), .A2(new_n572), .A3(new_n282), .A4(new_n566), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n430), .A2(new_n552), .A3(new_n557), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT35), .B1(new_n567), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n570), .A2(KEYINPUT83), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT83), .B1(new_n570), .B2(new_n576), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT90), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n295), .A2(new_n337), .A3(new_n338), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n293), .A2(new_n335), .A3(new_n294), .ZN(new_n582));
  NAND2_X1  g381(.A1(G229gat), .A2(G233gat), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT18), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n587));
  XNOR2_X1  g386(.A(G113gat), .B(G141gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G169gat), .B(G197gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n591), .B(KEYINPUT12), .Z(new_n592));
  NAND2_X1  g391(.A1(new_n586), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n581), .A2(KEYINPUT18), .A3(new_n582), .A4(new_n583), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n583), .B(KEYINPUT88), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT13), .ZN(new_n596));
  INV_X1    g395(.A(new_n582), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n335), .B1(new_n293), .B2(new_n294), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n580), .B1(new_n593), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n592), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n602), .B1(new_n584), .B2(new_n585), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n603), .A2(KEYINPUT90), .A3(new_n599), .A4(new_n594), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n586), .B1(new_n600), .B2(KEYINPUT89), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT89), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n607), .B1(new_n594), .B2(new_n599), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n602), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT91), .B1(new_n579), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT91), .ZN(new_n612));
  INV_X1    g411(.A(new_n610), .ZN(new_n613));
  NOR4_X1   g412(.A1(new_n577), .A2(new_n578), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n392), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n570), .A2(new_n576), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT83), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n570), .A2(new_n576), .A3(KEYINPUT83), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n612), .B1(new_n622), .B2(new_n613), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n579), .A2(KEYINPUT91), .A3(new_n610), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(KEYINPUT99), .A3(new_n392), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n282), .B1(new_n617), .B2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(new_n285), .ZN(G1324gat));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT16), .B(G8gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT100), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT42), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT99), .B1(new_n625), .B2(new_n392), .ZN(new_n634));
  AOI211_X1 g433(.A(new_n616), .B(new_n391), .C1(new_n623), .C2(new_n624), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n497), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n566), .B1(new_n617), .B2(new_n626), .ZN(new_n637));
  INV_X1    g436(.A(G8gat), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n631), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT42), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n629), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n497), .B1(new_n634), .B2(new_n635), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n632), .B1(new_n643), .B2(new_n631), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(G8gat), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n644), .A2(KEYINPUT101), .A3(new_n636), .A4(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n646), .ZN(G1325gat));
  INV_X1    g446(.A(G15gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n562), .A2(new_n565), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  AOI211_X1 g449(.A(new_n648), .B(new_n650), .C1(new_n617), .C2(new_n626), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n564), .B1(new_n634), .B2(new_n635), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n648), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n652), .A2(KEYINPUT102), .A3(new_n648), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n651), .B1(new_n655), .B2(new_n656), .ZN(G1326gat));
  AOI21_X1  g456(.A(new_n430), .B1(new_n617), .B2(new_n626), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT43), .B(G22gat), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1327gat));
  NAND3_X1  g459(.A1(new_n579), .A2(KEYINPUT44), .A3(new_n361), .ZN(new_n661));
  INV_X1    g460(.A(new_n361), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n662), .B1(new_n570), .B2(new_n576), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n663), .A2(KEYINPUT44), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n320), .A2(new_n613), .A3(new_n389), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n661), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(KEYINPUT103), .ZN(new_n667));
  INV_X1    g466(.A(new_n282), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n661), .A2(new_n669), .A3(new_n664), .A4(new_n665), .ZN(new_n670));
  AND3_X1   g469(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT45), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n321), .A2(new_n361), .A3(new_n390), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n623), .B2(new_n624), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n282), .A2(G29gat), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n674), .A2(new_n672), .A3(new_n675), .ZN(new_n677));
  OAI22_X1  g476(.A1(new_n671), .A2(new_n322), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT104), .ZN(G1328gat));
  NAND3_X1  g478(.A1(new_n667), .A2(new_n497), .A3(new_n670), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n323), .B1(new_n680), .B2(KEYINPUT105), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n681), .B1(KEYINPUT105), .B2(new_n680), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n674), .A2(new_n323), .A3(new_n497), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n683), .B(KEYINPUT46), .Z(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(G1329gat));
  INV_X1    g484(.A(G43gat), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n674), .A2(new_n686), .A3(new_n564), .ZN(new_n687));
  OAI21_X1  g486(.A(G43gat), .B1(new_n666), .B2(new_n650), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(new_n688), .A3(KEYINPUT47), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n667), .A2(new_n649), .A3(new_n670), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(G43gat), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n691), .A2(new_n687), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n689), .B1(new_n692), .B2(KEYINPUT47), .ZN(G1330gat));
  AND2_X1   g492(.A1(new_n661), .A2(new_n664), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(new_n568), .A3(new_n665), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n408), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n697), .B1(new_n696), .B2(new_n695), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n674), .A2(new_n408), .A3(new_n568), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(KEYINPUT48), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n699), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n667), .A2(new_n568), .A3(new_n670), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(G50gat), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n700), .B1(KEYINPUT48), .B2(new_n703), .ZN(G1331gat));
  NOR3_X1   g503(.A1(new_n321), .A2(new_n361), .A3(new_n390), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n618), .A2(new_n705), .A3(new_n613), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n282), .B(KEYINPUT107), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT108), .B(G57gat), .Z(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1332gat));
  XNOR2_X1  g509(.A(new_n706), .B(KEYINPUT109), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n497), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT49), .B(G64gat), .Z(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n712), .B2(new_n714), .ZN(G1333gat));
  NAND2_X1  g514(.A1(new_n711), .A2(new_n649), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n558), .A2(G71gat), .ZN(new_n717));
  AOI22_X1  g516(.A1(new_n716), .A2(G71gat), .B1(new_n706), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n718), .A2(new_n719), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT50), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  OR2_X1    g523(.A1(new_n718), .A2(new_n719), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT50), .B1(new_n725), .B2(new_n720), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n724), .A2(new_n726), .ZN(G1334gat));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n568), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g528(.A1(new_n320), .A2(new_n610), .A3(new_n390), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n694), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(G85gat), .B1(new_n731), .B2(new_n282), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n663), .A2(new_n613), .A3(new_n321), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT51), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n668), .A2(new_n389), .A3(new_n342), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT111), .Z(new_n739));
  OAI21_X1  g538(.A(new_n732), .B1(new_n737), .B2(new_n739), .ZN(G1336gat));
  OAI21_X1  g539(.A(G92gat), .B1(new_n731), .B2(new_n566), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n737), .A2(new_n390), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n742), .A2(new_n343), .A3(new_n497), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g544(.A(G99gat), .B1(new_n731), .B2(new_n650), .ZN(new_n746));
  INV_X1    g545(.A(G99gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n742), .A2(new_n747), .A3(new_n564), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(G1338gat));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n661), .A2(new_n568), .A3(new_n664), .A4(new_n730), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G106gat), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n430), .A2(G106gat), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n389), .B(new_n753), .C1(new_n735), .C2(new_n736), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n750), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(G106gat), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n756), .B1(new_n751), .B2(KEYINPUT112), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(KEYINPUT112), .B2(new_n751), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n754), .A2(new_n750), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n755), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1339gat));
  NAND2_X1  g561(.A1(new_n392), .A2(new_n613), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT54), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n386), .B1(new_n376), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n374), .A2(KEYINPUT114), .A3(new_n365), .A4(new_n375), .ZN(new_n766));
  INV_X1    g565(.A(new_n375), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n767), .B1(new_n377), .B2(new_n371), .ZN(new_n768));
  OAI211_X1 g567(.A(KEYINPUT54), .B(new_n766), .C1(new_n768), .C2(new_n365), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n374), .A2(new_n365), .A3(new_n375), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g571(.A(KEYINPUT55), .B(new_n765), .C1(new_n769), .C2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n374), .A2(new_n375), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n378), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n775), .B(new_n386), .C1(new_n378), .C2(new_n377), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n770), .A2(new_n771), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n778), .A2(new_n775), .A3(KEYINPUT54), .A4(new_n766), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n765), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT115), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783));
  AOI211_X1 g582(.A(new_n783), .B(KEYINPUT55), .C1(new_n779), .C2(new_n765), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n777), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n591), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n583), .B1(new_n581), .B2(new_n582), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n597), .A2(new_n598), .A3(new_n596), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n361), .A2(new_n605), .A3(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n605), .A2(new_n389), .A3(new_n789), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n785), .B2(new_n613), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n791), .B1(new_n793), .B2(new_n662), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n321), .B1(new_n794), .B2(KEYINPUT116), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n610), .B(new_n777), .C1(new_n782), .C2(new_n784), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n361), .B1(new_n796), .B2(new_n792), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n797), .A2(new_n798), .A3(new_n791), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n763), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n568), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n802), .A2(new_n668), .A3(new_n564), .A4(new_n566), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n803), .A2(new_n221), .A3(new_n613), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n800), .A2(new_n707), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n805), .A2(new_n497), .A3(new_n574), .ZN(new_n806));
  AOI21_X1  g605(.A(G113gat), .B1(new_n806), .B2(new_n610), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n804), .A2(new_n807), .ZN(G1340gat));
  NOR3_X1   g607(.A1(new_n803), .A2(new_n219), .A3(new_n390), .ZN(new_n809));
  AOI21_X1  g608(.A(G120gat), .B1(new_n806), .B2(new_n389), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(G1341gat));
  OAI21_X1  g610(.A(G127gat), .B1(new_n803), .B2(new_n321), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n806), .A2(new_n214), .A3(new_n320), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(G1342gat));
  NAND2_X1  g613(.A1(new_n361), .A2(new_n566), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT117), .ZN(new_n816));
  OR4_X1    g615(.A1(G134gat), .A2(new_n805), .A3(new_n574), .A4(new_n816), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n817), .A2(KEYINPUT56), .ZN(new_n818));
  OAI21_X1  g617(.A(G134gat), .B1(new_n803), .B2(new_n662), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(KEYINPUT56), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(G1343gat));
  NOR2_X1   g620(.A1(new_n649), .A2(new_n430), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n822), .B1(new_n805), .B2(KEYINPUT119), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n824), .B1(new_n800), .B2(new_n707), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n613), .A2(G141gat), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NOR4_X1   g626(.A1(new_n823), .A2(new_n497), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(KEYINPUT58), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n649), .A2(new_n282), .A3(new_n497), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT57), .B1(new_n800), .B2(new_n568), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n780), .A2(new_n781), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n610), .A2(new_n777), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n792), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n662), .ZN(new_n835));
  INV_X1    g634(.A(new_n791), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n320), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(new_n613), .B2(new_n392), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n430), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n830), .B1(new_n831), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G141gat), .B1(new_n843), .B2(new_n613), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(KEYINPUT118), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n847), .B(new_n830), .C1(new_n831), .C2(new_n842), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(new_n610), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n828), .B1(new_n849), .B2(G141gat), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT58), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n845), .B1(new_n850), .B2(new_n851), .ZN(G1344gat));
  NOR3_X1   g651(.A1(new_n823), .A2(new_n497), .A3(new_n825), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n382), .A3(new_n389), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n382), .A2(KEYINPUT59), .ZN(new_n855));
  INV_X1    g654(.A(new_n848), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n793), .A2(new_n662), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(KEYINPUT116), .A3(new_n836), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n798), .B1(new_n797), .B2(new_n791), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n858), .A2(new_n859), .A3(new_n321), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n430), .B1(new_n860), .B2(new_n763), .ZN(new_n861));
  OAI22_X1  g660(.A1(new_n861), .A2(KEYINPUT57), .B1(new_n841), .B2(new_n838), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n847), .B1(new_n862), .B2(new_n830), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n856), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n855), .B1(new_n864), .B2(new_n389), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n830), .A2(new_n389), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n839), .B1(new_n838), .B2(new_n430), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n800), .A2(new_n840), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT59), .B1(new_n869), .B2(new_n382), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g671(.A(KEYINPUT120), .B(KEYINPUT59), .C1(new_n869), .C2(new_n382), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n854), .B1(new_n865), .B2(new_n874), .ZN(G1345gat));
  NAND2_X1  g674(.A1(new_n846), .A2(new_n848), .ZN(new_n876));
  OAI21_X1  g675(.A(G155gat), .B1(new_n876), .B2(new_n321), .ZN(new_n877));
  INV_X1    g676(.A(G155gat), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n853), .A2(new_n878), .A3(new_n320), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(G1346gat));
  OAI21_X1  g679(.A(G162gat), .B1(new_n876), .B2(new_n662), .ZN(new_n881));
  OR4_X1    g680(.A1(G162gat), .A2(new_n823), .A3(new_n816), .A4(new_n825), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(G1347gat));
  NOR2_X1   g682(.A1(new_n801), .A2(new_n668), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n574), .A2(new_n566), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT121), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(G169gat), .B1(new_n887), .B2(new_n610), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n707), .A2(new_n566), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n564), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT122), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n802), .A2(new_n891), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n892), .A2(new_n448), .A3(new_n613), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n888), .A2(new_n893), .ZN(G1348gat));
  NAND3_X1  g693(.A1(new_n887), .A2(new_n449), .A3(new_n389), .ZN(new_n895));
  OAI21_X1  g694(.A(G176gat), .B1(new_n892), .B2(new_n390), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1349gat));
  NOR2_X1   g696(.A1(new_n321), .A2(new_n440), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n887), .A2(new_n898), .B1(new_n899), .B2(KEYINPUT60), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n899), .A2(KEYINPUT60), .ZN(new_n901));
  INV_X1    g700(.A(G183gat), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n800), .A2(new_n430), .A3(new_n891), .A4(new_n320), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(KEYINPUT123), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n904), .B1(KEYINPUT123), .B2(new_n903), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n900), .A2(new_n901), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n901), .B1(new_n900), .B2(new_n905), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(G1350gat));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n802), .A2(new_n361), .A3(new_n891), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(G190gat), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n662), .A2(G190gat), .ZN(new_n913));
  AOI22_X1  g712(.A1(new_n911), .A2(new_n912), .B1(new_n887), .B2(new_n913), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n911), .A2(new_n912), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n910), .A2(new_n909), .A3(G190gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(G1351gat));
  NOR3_X1   g716(.A1(new_n649), .A2(new_n566), .A3(new_n430), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n884), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(G197gat), .B1(new_n920), .B2(new_n610), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n867), .A2(new_n868), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT126), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT126), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n867), .A2(new_n868), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n650), .A2(new_n889), .ZN(new_n927));
  INV_X1    g726(.A(G197gat), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n927), .A2(new_n928), .A3(new_n613), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n921), .B1(new_n926), .B2(new_n929), .ZN(G1352gat));
  NOR2_X1   g729(.A1(new_n390), .A2(G204gat), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT127), .B1(new_n919), .B2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT62), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n884), .A2(new_n935), .A3(new_n918), .A4(new_n931), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n934), .B1(new_n933), .B2(new_n936), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n927), .B1(new_n923), .B2(new_n925), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n939), .A2(new_n389), .ZN(new_n940));
  INV_X1    g739(.A(G204gat), .ZN(new_n941));
  OAI22_X1  g740(.A1(new_n937), .A2(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G1353gat));
  INV_X1    g741(.A(G211gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n920), .A2(new_n943), .A3(new_n320), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n927), .A2(new_n321), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n943), .B1(new_n922), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT63), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n946), .A2(KEYINPUT63), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n944), .B1(new_n948), .B2(new_n949), .ZN(G1354gat));
  AOI21_X1  g749(.A(G218gat), .B1(new_n920), .B2(new_n361), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n361), .A2(G218gat), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n951), .B1(new_n939), .B2(new_n952), .ZN(G1355gat));
endmodule


