//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n211, new_n212, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G50), .ZN(new_n207));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT65), .ZN(G353));
  NOR2_X1   g0010(.A1(G97), .A2(G107), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G87), .ZN(G355));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT0), .Z(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT67), .B(G77), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  XOR2_X1   g0020(.A(KEYINPUT66), .B(G238), .Z(new_n221));
  OAI211_X1 g0021(.A(new_n219), .B(new_n220), .C1(new_n203), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT68), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n222), .A2(KEYINPUT68), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n214), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n206), .A2(G50), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n217), .B(new_n229), .C1(new_n232), .C2(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT69), .ZN(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G68), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n203), .A2(G50), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n247), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  INV_X1    g0055(.A(G45), .ZN(new_n256));
  AOI21_X1  g0056(.A(G1), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G274), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G1), .A3(G13), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(new_n257), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n263), .A2(G226), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT3), .B(G33), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(G222), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n218), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(G1698), .ZN(new_n269));
  INV_X1    g0069(.A(G223), .ZN(new_n270));
  OAI221_X1 g0070(.A(new_n267), .B1(new_n268), .B2(new_n265), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  AOI211_X1 g0071(.A(new_n259), .B(new_n264), .C1(new_n271), .C2(new_n262), .ZN(new_n272));
  INV_X1    g0072(.A(G200), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n274), .B1(G190), .B2(new_n272), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT10), .ZN(new_n276));
  XOR2_X1   g0076(.A(KEYINPUT8), .B(G58), .Z(new_n277));
  NAND2_X1  g0077(.A1(new_n231), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n277), .A2(new_n279), .B1(G150), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(new_n207), .B2(new_n231), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n230), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G1), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(G13), .A3(G20), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(G50), .ZN(new_n288));
  INV_X1    g0088(.A(new_n284), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n289), .B1(G1), .B2(new_n231), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n288), .B1(new_n291), .B2(G50), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n285), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT71), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n295), .A2(KEYINPUT9), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(KEYINPUT9), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n293), .A2(new_n295), .A3(KEYINPUT9), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AND3_X1   g0100(.A1(new_n275), .A2(new_n276), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n276), .B1(new_n275), .B2(new_n300), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G179), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n272), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n305), .B(new_n293), .C1(G169), .C2(new_n272), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n290), .A2(new_n208), .B1(new_n218), .B2(new_n287), .ZN(new_n307));
  XOR2_X1   g0107(.A(KEYINPUT15), .B(G87), .Z(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n279), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n218), .A2(G20), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT70), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n277), .B1(new_n311), .B2(new_n280), .ZN(new_n312));
  INV_X1    g0112(.A(new_n280), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(KEYINPUT70), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n309), .B(new_n310), .C1(new_n312), .C2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n307), .B1(new_n315), .B2(new_n284), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n265), .A2(G232), .A3(new_n266), .ZN(new_n317));
  INV_X1    g0117(.A(G107), .ZN(new_n318));
  OAI221_X1 g0118(.A(new_n317), .B1(new_n318), .B2(new_n265), .C1(new_n269), .C2(new_n221), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n262), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n263), .A2(G244), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n258), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G169), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n316), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n322), .B1(new_n319), .B2(new_n262), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n304), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n324), .A2(G200), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n327), .A2(G190), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(new_n331), .A3(new_n316), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n303), .A2(new_n306), .A3(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(KEYINPUT72), .B1(new_n313), .B2(new_n248), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n279), .A2(G77), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n203), .A2(G20), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  OR3_X1    g0138(.A1(new_n313), .A2(KEYINPUT72), .A3(new_n248), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n289), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT11), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT12), .ZN(new_n342));
  INV_X1    g0142(.A(new_n287), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n342), .B1(new_n343), .B2(new_n203), .ZN(new_n344));
  NOR3_X1   g0144(.A1(new_n287), .A2(KEYINPUT12), .A3(G68), .ZN(new_n345));
  OAI221_X1 g0145(.A(new_n341), .B1(new_n203), .B2(new_n290), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n340), .A2(KEYINPUT11), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT13), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n265), .A2(G232), .A3(G1698), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n265), .A2(G226), .A3(new_n266), .ZN(new_n352));
  INV_X1    g0152(.A(G33), .ZN(new_n353));
  INV_X1    g0153(.A(G97), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n351), .B(new_n352), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n262), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n259), .B1(new_n263), .B2(G238), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n350), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n356), .A2(new_n350), .A3(new_n357), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(G179), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n325), .B1(new_n359), .B2(new_n360), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT14), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n360), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n363), .B(G169), .C1(new_n365), .C2(new_n358), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n349), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n365), .A2(new_n358), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G190), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n348), .B(new_n370), .C1(new_n273), .C2(new_n369), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G190), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n286), .B1(G41), .B2(G45), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n261), .A2(G232), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n258), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n353), .A2(KEYINPUT3), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT3), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G33), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n377), .A2(new_n379), .A3(G226), .A4(G1698), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n377), .A2(new_n379), .A3(G223), .A4(new_n266), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G33), .A2(G87), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  AOI211_X1 g0183(.A(new_n373), .B(new_n376), .C1(new_n262), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n262), .ZN(new_n385));
  INV_X1    g0185(.A(new_n376), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n273), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n277), .A2(new_n343), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n389), .B1(new_n290), .B2(new_n277), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n265), .B2(G20), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT73), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n378), .A2(G33), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n353), .A2(KEYINPUT3), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT7), .B(new_n231), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n393), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  AOI211_X1 g0198(.A(new_n392), .B(G20), .C1(new_n377), .C2(new_n379), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT73), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(G68), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G58), .A2(G68), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n204), .A2(new_n205), .A3(new_n402), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n403), .A2(G20), .B1(G159), .B2(new_n280), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT16), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n377), .A2(new_n379), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT7), .B1(new_n406), .B2(new_n231), .ZN(new_n407));
  OAI21_X1  g0207(.A(G68), .B1(new_n407), .B2(new_n399), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(KEYINPUT16), .A3(new_n404), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n284), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n388), .B(new_n391), .C1(new_n405), .C2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT17), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n401), .A2(new_n404), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT16), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n203), .B1(new_n393), .B2(new_n397), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n403), .A2(G20), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n280), .A2(G159), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n289), .B1(new_n420), .B2(KEYINPUT16), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT17), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n422), .A2(new_n423), .A3(new_n391), .A4(new_n388), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n412), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n390), .B1(new_n415), .B2(new_n421), .ZN(new_n427));
  AOI211_X1 g0227(.A(new_n304), .B(new_n376), .C1(new_n262), .C2(new_n383), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n325), .B1(new_n385), .B2(new_n386), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT18), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n391), .B1(new_n410), .B2(new_n405), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT18), .ZN(new_n433));
  INV_X1    g0233(.A(new_n430), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n426), .A2(new_n437), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n334), .A2(new_n372), .A3(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n377), .A2(new_n379), .A3(G244), .A4(new_n266), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT4), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n265), .A2(KEYINPUT4), .A3(G244), .A4(new_n266), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n265), .A2(G250), .A3(G1698), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G33), .A2(G283), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n442), .A2(new_n443), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n262), .ZN(new_n447));
  AND2_X1   g0247(.A1(KEYINPUT5), .A2(G41), .ZN(new_n448));
  NOR2_X1   g0248(.A1(KEYINPUT5), .A2(G41), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n286), .A2(G45), .A3(G274), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g0252(.A(KEYINPUT5), .B(G41), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n256), .A2(G1), .ZN(new_n454));
  INV_X1    g0254(.A(new_n230), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n453), .A2(new_n454), .B1(new_n455), .B2(new_n260), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n452), .B1(new_n456), .B2(G257), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n447), .A2(G179), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n325), .B1(new_n447), .B2(new_n457), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n211), .A2(KEYINPUT6), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT6), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G97), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n318), .A2(KEYINPUT75), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT75), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G107), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n461), .A2(new_n463), .A3(new_n465), .A4(new_n467), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(G20), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n280), .A2(G77), .ZN(new_n472));
  XOR2_X1   g0272(.A(new_n472), .B(KEYINPUT74), .Z(new_n473));
  AND2_X1   g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n398), .A2(G107), .A3(new_n400), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n289), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n287), .A2(G97), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n286), .A2(G33), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n287), .A2(new_n479), .A3(new_n230), .A4(new_n283), .ZN(new_n480));
  XNOR2_X1  g0280(.A(new_n480), .B(KEYINPUT76), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n478), .B1(new_n481), .B2(new_n354), .ZN(new_n482));
  OAI22_X1  g0282(.A1(new_n459), .A2(new_n460), .B1(new_n476), .B2(new_n482), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n398), .A2(G107), .A3(new_n400), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n471), .A2(new_n473), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n284), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n482), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n447), .A2(new_n373), .A3(new_n457), .ZN(new_n488));
  AOI21_X1  g0288(.A(G200), .B1(new_n447), .B2(new_n457), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n486), .B(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n483), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n377), .A2(new_n379), .A3(G244), .A4(G1698), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n377), .A2(new_n379), .A3(G238), .A4(new_n266), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G116), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n262), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n286), .A2(G45), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n261), .A2(G250), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n451), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT77), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n498), .A2(KEYINPUT77), .A3(new_n451), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n496), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(KEYINPUT78), .B1(new_n503), .B2(G179), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n498), .A2(KEYINPUT77), .A3(new_n451), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT77), .B1(new_n498), .B2(new_n451), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT78), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n507), .A2(new_n508), .A3(new_n304), .A4(new_n496), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n503), .A2(new_n325), .ZN(new_n510));
  NAND3_X1  g0310(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n231), .ZN(new_n512));
  XNOR2_X1  g0312(.A(KEYINPUT79), .B(G87), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(new_n212), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n377), .A2(new_n379), .A3(new_n231), .A4(G68), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT19), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n278), .B2(new_n354), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n284), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n308), .A2(new_n287), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n308), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n520), .B(new_n522), .C1(new_n523), .C2(new_n481), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n504), .A2(new_n509), .A3(new_n510), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n503), .A2(G200), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n507), .A2(G190), .A3(new_n496), .ZN(new_n527));
  INV_X1    g0327(.A(new_n519), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n289), .B1(new_n528), .B2(new_n514), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n529), .A2(new_n521), .ZN(new_n530));
  INV_X1    g0330(.A(new_n481), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G87), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n526), .A2(new_n527), .A3(new_n530), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n491), .A2(KEYINPUT80), .A3(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT80), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n483), .A2(new_n490), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(new_n534), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n377), .A2(new_n379), .A3(G257), .A4(new_n266), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n377), .A2(new_n379), .A3(G264), .A4(G1698), .ZN(new_n541));
  INV_X1    g0341(.A(G303), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n540), .B(new_n541), .C1(new_n542), .C2(new_n265), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n262), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n452), .B1(new_n456), .B2(G270), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(G116), .ZN(new_n547));
  OR2_X1    g0347(.A1(new_n480), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n343), .A2(new_n547), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n283), .A2(new_n230), .B1(G20), .B2(new_n547), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n445), .B(new_n231), .C1(G33), .C2(new_n354), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n550), .A2(KEYINPUT20), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT20), .B1(new_n550), .B2(new_n551), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n548), .B(new_n549), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n546), .A2(new_n554), .A3(G169), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT21), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n554), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n544), .A2(new_n545), .A3(G190), .ZN(new_n559));
  INV_X1    g0359(.A(new_n546), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n558), .B(new_n559), .C1(new_n560), .C2(new_n273), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n546), .A2(new_n554), .A3(KEYINPUT21), .A4(G169), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n554), .A2(G179), .A3(new_n544), .A4(new_n545), .ZN(new_n563));
  AND4_X1   g0363(.A1(new_n557), .A2(new_n561), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n287), .A2(G107), .ZN(new_n565));
  XNOR2_X1  g0365(.A(new_n565), .B(KEYINPUT25), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n481), .B2(new_n318), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT23), .B1(new_n231), .B2(G107), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT23), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(new_n318), .A3(G20), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n231), .A2(G33), .A3(G116), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT82), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n568), .A2(new_n570), .A3(new_n571), .A4(KEYINPUT82), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AND2_X1   g0376(.A1(KEYINPUT81), .A2(G87), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n265), .A2(new_n231), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT22), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n265), .A2(KEYINPUT22), .A3(new_n231), .A4(new_n577), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n576), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT24), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n289), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n576), .A2(KEYINPUT24), .A3(new_n580), .A4(new_n581), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n567), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n377), .A2(new_n379), .A3(G250), .A4(new_n266), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT83), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT83), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n265), .A2(new_n590), .A3(G250), .A4(new_n266), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G294), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n265), .A2(G257), .A3(G1698), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n589), .A2(new_n591), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n262), .ZN(new_n595));
  INV_X1    g0395(.A(new_n452), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n454), .B1(new_n448), .B2(new_n449), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n597), .A2(G264), .A3(new_n261), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n595), .A2(new_n304), .A3(new_n596), .A4(new_n599), .ZN(new_n600));
  AOI211_X1 g0400(.A(new_n452), .B(new_n598), .C1(new_n594), .C2(new_n262), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n600), .B1(new_n601), .B2(G169), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n587), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n595), .A2(new_n596), .A3(new_n599), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G200), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n586), .B(new_n606), .C1(new_n373), .C2(new_n605), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n564), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  AND4_X1   g0408(.A1(new_n439), .A2(new_n536), .A3(new_n539), .A4(new_n608), .ZN(G372));
  AND4_X1   g0409(.A1(new_n532), .A2(new_n526), .A3(new_n530), .A4(new_n527), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT76), .ZN(new_n611));
  OR2_X1    g0411(.A1(new_n480), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n480), .A2(new_n611), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n523), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n614), .A2(new_n529), .A3(new_n521), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n507), .A2(new_n304), .A3(new_n496), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n510), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT84), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n615), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n510), .A2(new_n616), .A3(KEYINPUT84), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n610), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n562), .A2(new_n563), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n622), .B(new_n557), .C1(new_n586), .C2(new_n602), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n491), .A2(new_n621), .A3(new_n623), .A4(new_n607), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT85), .B1(new_n459), .B2(new_n460), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n486), .A2(new_n487), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT85), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n447), .A2(new_n457), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n627), .B(new_n458), .C1(new_n628), .C2(new_n325), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n625), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n621), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n503), .A2(G179), .ZN(new_n633));
  AOI21_X1  g0433(.A(G169), .B1(new_n507), .B2(new_n496), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n618), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n635), .A2(new_n620), .A3(new_n524), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n458), .B1(new_n628), .B2(new_n325), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n525), .A2(new_n637), .A3(new_n626), .A4(new_n533), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n636), .B1(KEYINPUT26), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n624), .A2(new_n632), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n439), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n306), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n368), .A2(new_n329), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n426), .A2(new_n371), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n437), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n642), .B1(new_n645), .B2(new_n303), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n641), .A2(new_n646), .ZN(G369));
  NAND2_X1  g0447(.A1(new_n622), .A2(new_n557), .ZN(new_n648));
  INV_X1    g0448(.A(G13), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(G20), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n286), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT27), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n650), .A2(new_n653), .A3(new_n286), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n652), .A2(G213), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT86), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n655), .B(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n657), .A2(G343), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n648), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n587), .A2(new_n603), .A3(new_n658), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT87), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n604), .B(new_n607), .C1(new_n586), .C2(new_n659), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT88), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n660), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n604), .A2(new_n658), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n659), .A2(new_n558), .ZN(new_n674));
  MUX2_X1   g0474(.A(new_n564), .B(new_n648), .S(new_n674), .Z(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G330), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n672), .A2(new_n679), .ZN(G399));
  NOR2_X1   g0480(.A1(new_n513), .A2(new_n212), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n547), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n215), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G41), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n683), .A2(G1), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n233), .B2(new_n686), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT89), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT28), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n640), .A2(new_n659), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(KEYINPUT29), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n534), .A2(new_n483), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n636), .B1(new_n693), .B2(new_n631), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n635), .A2(new_n620), .A3(new_n524), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n533), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n625), .A2(new_n629), .A3(new_n626), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT26), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT90), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT90), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n694), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(new_n624), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n659), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n692), .B1(new_n704), .B2(KEYINPUT29), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n608), .A2(new_n536), .A3(new_n539), .A4(new_n659), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT31), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n628), .A2(G179), .A3(new_n560), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT30), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n595), .A2(new_n507), .A3(new_n496), .A4(new_n599), .ZN(new_n710));
  OR3_X1    g0510(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n503), .A2(new_n304), .ZN(new_n712));
  OR4_X1    g0512(.A1(new_n628), .A2(new_n601), .A3(new_n712), .A4(new_n560), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n709), .B1(new_n708), .B2(new_n710), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n711), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n707), .B1(new_n715), .B2(new_n658), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n706), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n715), .A2(new_n707), .A3(new_n658), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n717), .A2(G330), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n705), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n690), .B1(new_n722), .B2(G1), .ZN(G364));
  AOI21_X1  g0523(.A(new_n286), .B1(new_n650), .B2(G45), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n685), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n678), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n676), .A2(new_n677), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G13), .A2(G33), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n231), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT92), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n676), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n230), .B1(G20), .B2(new_n325), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G179), .A2(G200), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n231), .B1(new_n736), .B2(G190), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n373), .A2(G20), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n304), .A2(new_n273), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI221_X1 g0541(.A(new_n265), .B1(new_n737), .B2(new_n354), .C1(new_n741), .C2(new_n203), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n304), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n231), .A2(new_n373), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n273), .A2(G179), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n745), .A2(new_n218), .B1(new_n749), .B2(new_n513), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n739), .A2(new_n747), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n746), .A2(new_n740), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n752), .A2(KEYINPUT95), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(KEYINPUT95), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n750), .B1(new_n318), .B2(new_n751), .C1(new_n756), .C2(new_n248), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n739), .A2(new_n736), .ZN(new_n758));
  INV_X1    g0558(.A(G159), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XOR2_X1   g0560(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n761));
  XNOR2_X1  g0561(.A(new_n760), .B(new_n761), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n746), .A2(new_n743), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n763), .A2(KEYINPUT94), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(KEYINPUT94), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n202), .ZN(new_n768));
  OR4_X1    g0568(.A1(new_n742), .A2(new_n757), .A3(new_n762), .A4(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n766), .A2(G322), .B1(new_n755), .B2(G326), .ZN(new_n770));
  INV_X1    g0570(.A(new_n758), .ZN(new_n771));
  AOI22_X1  g0571(.A1(G329), .A2(new_n771), .B1(new_n745), .B2(G311), .ZN(new_n772));
  INV_X1    g0572(.A(new_n741), .ZN(new_n773));
  XNOR2_X1  g0573(.A(KEYINPUT33), .B(G317), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n749), .A2(G303), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G283), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n406), .B1(new_n751), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n737), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n777), .B1(G294), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n770), .A2(new_n772), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n735), .B1(new_n769), .B2(new_n780), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n726), .B(KEYINPUT91), .Z(new_n782));
  NAND3_X1  g0582(.A1(G355), .A2(new_n265), .A3(new_n215), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n253), .A2(new_n256), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n684), .A2(new_n265), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(new_n233), .B2(G45), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n783), .B1(G116), .B2(new_n215), .C1(new_n784), .C2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n732), .A2(new_n734), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n782), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g0589(.A1(new_n789), .A2(KEYINPUT93), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(KEYINPUT93), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n781), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n727), .A2(new_n728), .B1(new_n733), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(G396));
  NAND2_X1  g0594(.A1(new_n315), .A2(new_n284), .ZN(new_n795));
  INV_X1    g0595(.A(new_n307), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n658), .A2(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n332), .A2(new_n798), .B1(new_n328), .B2(new_n326), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n329), .A2(new_n658), .ZN(new_n800));
  OAI21_X1  g0600(.A(KEYINPUT99), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT99), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n659), .A2(new_n328), .A3(new_n326), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n797), .B1(G190), .B2(new_n327), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n804), .A2(new_n330), .B1(new_n797), .B2(new_n658), .ZN(new_n805));
  INV_X1    g0605(.A(new_n329), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n802), .B(new_n803), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n801), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n691), .B(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n726), .B1(new_n809), .B2(new_n719), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n719), .B2(new_n809), .ZN(new_n811));
  INV_X1    g0611(.A(new_n782), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n734), .A2(new_n729), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT97), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n812), .B1(new_n815), .B2(G77), .ZN(new_n816));
  INV_X1    g0616(.A(G87), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n751), .A2(new_n817), .B1(new_n748), .B2(new_n318), .ZN(new_n818));
  INV_X1    g0618(.A(G311), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n406), .B1(new_n737), .B2(new_n354), .C1(new_n758), .C2(new_n819), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n818), .B(new_n820), .C1(G116), .C2(new_n745), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n766), .A2(G294), .B1(new_n755), .B2(G303), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n773), .A2(KEYINPUT98), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n773), .A2(KEYINPUT98), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n821), .B(new_n822), .C1(new_n776), .C2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(G150), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n741), .A2(new_n827), .B1(new_n744), .B2(new_n759), .ZN(new_n828));
  INV_X1    g0628(.A(G137), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n756), .A2(new_n829), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n828), .B(new_n830), .C1(G143), .C2(new_n766), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n831), .A2(KEYINPUT34), .ZN(new_n832));
  INV_X1    g0632(.A(G132), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n265), .B1(new_n758), .B2(new_n833), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n751), .A2(new_n203), .B1(new_n748), .B2(new_n248), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n834), .B(new_n835), .C1(G58), .C2(new_n778), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n831), .B2(KEYINPUT34), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n826), .B1(new_n832), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n816), .B1(new_n838), .B2(new_n734), .ZN(new_n839));
  INV_X1    g0639(.A(new_n729), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n808), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n811), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G384));
  OAI21_X1  g0643(.A(new_n414), .B1(new_n416), .B2(new_n419), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n409), .A2(new_n844), .A3(new_n284), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT101), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n845), .A2(new_n846), .A3(new_n391), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n846), .B1(new_n845), .B2(new_n391), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n657), .A2(new_n428), .A3(new_n429), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n411), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT37), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT37), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n411), .B(new_n853), .C1(new_n427), .C2(new_n849), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n655), .B(KEYINPUT86), .ZN(new_n856));
  NOR3_X1   g0656(.A1(new_n847), .A2(new_n848), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n425), .B2(new_n436), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n855), .A2(new_n858), .A3(KEYINPUT38), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT104), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT104), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n855), .A2(new_n858), .A3(new_n861), .A4(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n427), .A2(new_n856), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n425), .B2(new_n436), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n411), .B1(new_n427), .B2(new_n849), .ZN(new_n866));
  OR3_X1    g0666(.A1(new_n866), .A2(KEYINPUT102), .A3(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(KEYINPUT37), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(KEYINPUT102), .A3(new_n854), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n865), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT103), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n871), .B1(new_n870), .B2(new_n872), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n863), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n349), .A2(new_n658), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n368), .A2(new_n371), .A3(new_n876), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n349), .B(new_n658), .C1(new_n364), .C2(new_n367), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n877), .A2(new_n878), .B1(new_n801), .B2(new_n807), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n717), .A3(new_n718), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT40), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n875), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n717), .A2(new_n718), .ZN(new_n884));
  INV_X1    g0684(.A(new_n859), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT38), .B1(new_n855), .B2(new_n858), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n881), .B1(new_n887), .B2(new_n880), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n883), .A2(new_n439), .A3(new_n884), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n870), .A2(new_n872), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT103), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n891), .A2(new_n892), .B1(new_n860), .B2(new_n862), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n884), .A2(KEYINPUT40), .A3(new_n879), .ZN(new_n894));
  OAI211_X1 g0694(.A(G330), .B(new_n888), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n439), .A2(new_n719), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n889), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n439), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n646), .B1(new_n705), .B2(new_n900), .ZN(new_n901));
  XOR2_X1   g0701(.A(new_n899), .B(new_n901), .Z(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n863), .B(new_n903), .C1(new_n874), .C2(new_n873), .ZN(new_n904));
  INV_X1    g0704(.A(new_n886), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n859), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT39), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n368), .A2(new_n658), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n877), .A2(new_n878), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n640), .A2(new_n659), .A3(new_n808), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT100), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n912), .A2(new_n913), .A3(new_n803), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n913), .B1(new_n912), .B2(new_n803), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n906), .B(new_n911), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n436), .A2(new_n856), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n910), .A2(KEYINPUT105), .A3(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT105), .ZN(new_n920));
  INV_X1    g0720(.A(new_n909), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n904), .B2(new_n907), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n916), .A2(new_n917), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n919), .A2(new_n924), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n902), .A2(new_n925), .B1(new_n286), .B2(new_n650), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n925), .B2(new_n902), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n469), .A2(new_n470), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n928), .A2(KEYINPUT35), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(KEYINPUT35), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n929), .A2(G116), .A3(new_n232), .A4(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT36), .Z(new_n932));
  NAND3_X1  g0732(.A1(new_n234), .A2(new_n218), .A3(new_n402), .ZN(new_n933));
  AOI211_X1 g0733(.A(new_n286), .B(G13), .C1(new_n933), .C2(new_n249), .ZN(new_n934));
  OR3_X1    g0734(.A1(new_n927), .A2(new_n932), .A3(new_n934), .ZN(G367));
  INV_X1    g0735(.A(new_n660), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n673), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n671), .ZN(new_n938));
  INV_X1    g0738(.A(new_n626), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n491), .B1(new_n939), .B2(new_n659), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n630), .A2(new_n658), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n937), .A2(new_n938), .A3(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT45), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n672), .A2(KEYINPUT45), .A3(new_n942), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT44), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n672), .B2(new_n942), .ZN(new_n949));
  INV_X1    g0749(.A(new_n942), .ZN(new_n950));
  OAI211_X1 g0750(.A(KEYINPUT44), .B(new_n950), .C1(new_n670), .C2(new_n671), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n947), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n679), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n947), .A2(new_n952), .A3(new_n679), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n668), .A2(new_n669), .A3(new_n660), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n937), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n678), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n958), .B(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n960), .A2(new_n721), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n955), .A2(new_n956), .A3(new_n961), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n962), .A2(KEYINPUT106), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(KEYINPUT106), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n722), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n685), .B(KEYINPUT41), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n725), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n670), .A2(new_n942), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n968), .A2(KEYINPUT42), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n950), .A2(new_n938), .B1(new_n483), .B2(new_n658), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n968), .B2(KEYINPUT42), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n530), .A2(new_n532), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n658), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n621), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n695), .B2(new_n973), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n969), .A2(new_n971), .B1(KEYINPUT43), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n976), .B(new_n977), .Z(new_n978));
  NOR2_X1   g0778(.A1(new_n679), .A2(new_n950), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n978), .B(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n975), .A2(new_n731), .ZN(new_n982));
  INV_X1    g0782(.A(new_n785), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n239), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n788), .B1(new_n215), .B2(new_n523), .ZN(new_n985));
  INV_X1    g0785(.A(new_n825), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n986), .A2(G159), .B1(new_n755), .B2(G143), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n268), .A2(new_n751), .B1(new_n744), .B2(new_n248), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n265), .B1(new_n737), .B2(new_n203), .C1(new_n758), .C2(new_n829), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n988), .B(new_n989), .C1(G58), .C2(new_n749), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n987), .B(new_n990), .C1(new_n827), .C2(new_n767), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n986), .A2(G294), .B1(G303), .B2(new_n766), .ZN(new_n992));
  INV_X1    g0792(.A(G317), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n406), .B1(new_n758), .B2(new_n993), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n354), .A2(new_n751), .B1(new_n744), .B2(new_n776), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(new_n755), .C2(G311), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n749), .A2(KEYINPUT46), .A3(G116), .ZN(new_n997));
  AOI21_X1  g0797(.A(KEYINPUT46), .B1(new_n749), .B2(G116), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G107), .B2(new_n778), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n992), .A2(new_n996), .A3(new_n997), .A4(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n991), .A2(new_n1000), .A3(KEYINPUT47), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n734), .ZN(new_n1002));
  AOI21_X1  g0802(.A(KEYINPUT47), .B1(new_n991), .B2(new_n1000), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n812), .B1(new_n984), .B2(new_n985), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT107), .Z(new_n1005));
  OAI22_X1  g0805(.A1(new_n967), .A2(new_n981), .B1(new_n982), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT108), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1005), .A2(new_n982), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n955), .A2(new_n956), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT106), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1010), .A2(new_n1011), .A3(new_n961), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n962), .A2(KEYINPUT106), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n721), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n966), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n724), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1009), .B1(new_n1016), .B2(new_n980), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(KEYINPUT108), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1008), .A2(new_n1018), .ZN(G387));
  INV_X1    g0819(.A(new_n960), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n668), .A2(new_n669), .A3(new_n732), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n785), .B1(new_n243), .B2(new_n256), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n682), .A2(new_n215), .A3(new_n265), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n277), .A2(new_n248), .ZN(new_n1025));
  XOR2_X1   g0825(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n1026));
  XNOR2_X1  g0826(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1027), .A2(new_n683), .A3(new_n1028), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n1024), .A2(new_n1029), .B1(new_n318), .B2(new_n684), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n788), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n812), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(KEYINPUT110), .B(G150), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n744), .A2(new_n203), .B1(new_n758), .B2(new_n1033), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n767), .A2(new_n248), .B1(new_n756), .B2(new_n759), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n277), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1036), .A2(new_n741), .B1(new_n268), .B2(new_n748), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n265), .B1(new_n751), .B2(new_n354), .C1(new_n523), .C2(new_n737), .ZN(new_n1038));
  OR4_X1    g0838(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n766), .A2(G317), .B1(new_n755), .B2(G322), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n542), .B2(new_n744), .C1(new_n819), .C2(new_n825), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT48), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n749), .A2(G294), .B1(new_n778), .B2(G283), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT111), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT49), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n406), .B1(new_n751), .B2(new_n547), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G326), .B2(new_n771), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1039), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1032), .B1(new_n1052), .B2(new_n734), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n1020), .A2(new_n725), .B1(new_n1021), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n685), .B1(new_n960), .B2(new_n721), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1020), .A2(new_n722), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1054), .B1(new_n1055), .B2(new_n1056), .ZN(G393));
  NOR2_X1   g0857(.A1(new_n1010), .A2(KEYINPUT112), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1058), .A2(new_n724), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1010), .A2(KEYINPUT112), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n950), .A2(new_n732), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n247), .A2(new_n983), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n788), .B1(new_n354), .B2(new_n215), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n812), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n766), .A2(G159), .B1(new_n755), .B2(G150), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT51), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n771), .A2(G143), .B1(new_n749), .B2(G68), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1067), .B(new_n265), .C1(new_n817), .C2(new_n751), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT113), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n778), .A2(G77), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n1036), .B2(new_n744), .C1(new_n825), .C2(new_n248), .ZN(new_n1071));
  OR3_X1    g0871(.A1(new_n1066), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1072), .A2(KEYINPUT114), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(KEYINPUT114), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n766), .A2(G311), .B1(new_n755), .B2(G317), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n1075), .A2(KEYINPUT52), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(KEYINPUT52), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n986), .A2(G303), .ZN(new_n1078));
  INV_X1    g0878(.A(G322), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n758), .A2(new_n1079), .B1(new_n748), .B2(new_n776), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n406), .B1(new_n737), .B2(new_n547), .C1(new_n751), .C2(new_n318), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1080), .B(new_n1081), .C1(G294), .C2(new_n745), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .A4(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1073), .A2(new_n1074), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1064), .B1(new_n1084), .B2(new_n734), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1059), .A2(new_n1060), .B1(new_n1061), .B2(new_n1085), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n685), .B1(new_n1010), .B2(new_n961), .C1(new_n963), .C2(new_n964), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(G390));
  INV_X1    g0888(.A(new_n624), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n699), .B2(KEYINPUT90), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n658), .B1(new_n1090), .B2(new_n702), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n800), .B1(new_n1091), .B2(new_n808), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n911), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n921), .B(new_n875), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n912), .A2(new_n803), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(KEYINPUT100), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n912), .A2(new_n913), .A3(new_n803), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n909), .B1(new_n1098), .B2(new_n911), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1094), .B1(new_n1099), .B2(new_n908), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n880), .A2(new_n677), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1093), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n907), .B(new_n904), .C1(new_n1103), .C2(new_n909), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1101), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1104), .A2(new_n1105), .A3(new_n1094), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n646), .B(new_n897), .C1(new_n705), .C2(new_n900), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n911), .B1(new_n719), .B2(new_n808), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1098), .B1(new_n1108), .B2(new_n1101), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n719), .A2(new_n808), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1105), .B(new_n1092), .C1(new_n1110), .C2(new_n911), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1107), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1102), .A2(new_n1106), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(KEYINPUT115), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT115), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1102), .A2(new_n1115), .A3(new_n1112), .A4(new_n1106), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1111), .A2(new_n1109), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1107), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n686), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(KEYINPUT116), .B1(new_n1117), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1102), .A2(new_n725), .A3(new_n1106), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n986), .A2(G137), .B1(new_n755), .B2(G128), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n748), .A2(new_n1033), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT53), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1126), .B(new_n1128), .C1(new_n833), .C2(new_n767), .ZN(new_n1129));
  XOR2_X1   g0929(.A(KEYINPUT54), .B(G143), .Z(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(G125), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n1131), .A2(new_n744), .B1(new_n1132), .B2(new_n758), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n751), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n406), .B1(new_n1135), .B2(G50), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1134), .B(new_n1136), .C1(new_n759), .C2(new_n737), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n986), .A2(G107), .B1(new_n755), .B2(G283), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n547), .B2(new_n767), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n771), .A2(G294), .B1(new_n749), .B2(G87), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n265), .B1(new_n1135), .B2(G68), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n745), .A2(G97), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1140), .A2(new_n1141), .A3(new_n1070), .A4(new_n1142), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1129), .A2(new_n1137), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n734), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n782), .B1(new_n1036), .B2(new_n814), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1145), .B(new_n1146), .C1(new_n908), .C2(new_n840), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1125), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1148), .A2(KEYINPUT117), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT117), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n1125), .B2(new_n1147), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1117), .A2(new_n1122), .A3(KEYINPUT116), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1124), .A2(new_n1152), .A3(new_n1153), .ZN(G378));
  XNOR2_X1  g0954(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n294), .A2(new_n856), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n303), .A2(new_n306), .A3(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n306), .B1(new_n301), .B2(new_n302), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n1156), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1155), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1158), .A2(new_n1160), .A3(new_n1155), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n729), .A3(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n265), .A2(G41), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G50), .B(new_n1165), .C1(new_n353), .C2(new_n255), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1165), .B1(new_n203), .B2(new_n737), .C1(new_n268), .C2(new_n748), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n741), .A2(new_n354), .B1(new_n758), .B2(new_n776), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n523), .A2(new_n744), .B1(new_n751), .B2(new_n202), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n547), .B2(new_n756), .C1(new_n318), .C2(new_n767), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT58), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1166), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n766), .A2(G128), .B1(new_n755), .B2(G125), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n741), .A2(new_n833), .B1(new_n744), .B2(new_n829), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n749), .B2(new_n1130), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1174), .B(new_n1176), .C1(new_n827), .C2(new_n737), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(KEYINPUT59), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1135), .A2(G159), .ZN(new_n1179));
  AOI211_X1 g0979(.A(G33), .B(G41), .C1(new_n771), .C2(G124), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1177), .A2(KEYINPUT59), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1173), .B1(new_n1172), .B2(new_n1171), .C1(new_n1181), .C2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n734), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n725), .B(new_n685), .C1(new_n248), .C2(new_n813), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1164), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1162), .A2(KEYINPUT118), .A3(new_n1163), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n895), .A2(new_n1188), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n883), .A2(new_n1187), .A3(G330), .A4(new_n888), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(KEYINPUT105), .B1(new_n910), .B2(new_n918), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n922), .A2(new_n923), .A3(new_n920), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1191), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1191), .A2(KEYINPUT119), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n919), .A2(new_n924), .A3(new_n1190), .A4(new_n1189), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n925), .A2(KEYINPUT119), .A3(new_n1191), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1186), .B1(new_n1199), .B2(new_n725), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1104), .A2(new_n1105), .A3(new_n1094), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1105), .B1(new_n1104), .B2(new_n1094), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1115), .B1(new_n1203), .B2(new_n1112), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1116), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1120), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT57), .B1(new_n1206), .B2(new_n1199), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1107), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1194), .A2(KEYINPUT57), .A3(new_n1196), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n685), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1200), .B1(new_n1207), .B2(new_n1210), .ZN(G375));
  NAND3_X1  g1011(.A1(new_n1111), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1121), .A2(new_n966), .A3(new_n1212), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n744), .A2(new_n318), .B1(new_n758), .B2(new_n542), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n406), .B1(new_n354), .B2(new_n748), .C1(new_n523), .C2(new_n737), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(G77), .C2(new_n1135), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n755), .A2(G294), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n767), .B2(new_n776), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G116), .B2(new_n986), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n825), .A2(new_n1131), .B1(new_n756), .B2(new_n833), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G137), .B2(new_n766), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n744), .A2(new_n827), .B1(new_n748), .B2(new_n759), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n265), .B1(new_n737), .B2(new_n248), .C1(new_n751), .C2(new_n202), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(G128), .C2(new_n771), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1216), .A2(new_n1219), .B1(new_n1221), .B2(new_n1224), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n812), .B1(G68), .B2(new_n815), .C1(new_n1225), .C2(new_n735), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1093), .B2(new_n729), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1119), .B2(new_n725), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1213), .A2(new_n1228), .ZN(G381));
  INV_X1    g1029(.A(new_n1209), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n686), .B1(new_n1206), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT57), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1232), .B1(new_n1233), .B2(new_n1208), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1231), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1148), .B1(new_n1117), .B2(new_n1122), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n1200), .A3(new_n1236), .ZN(new_n1237));
  OR4_X1    g1037(.A1(G396), .A2(G393), .A3(G384), .A4(G381), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(G390), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1008), .A2(new_n1018), .A3(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT120), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1237), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1008), .A2(new_n1018), .A3(KEYINPUT120), .A4(new_n1239), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT121), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1242), .A2(KEYINPUT121), .A3(new_n1243), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(G407));
  INV_X1    g1047(.A(G213), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1237), .ZN(new_n1249));
  OR3_X1    g1049(.A1(new_n1248), .A2(KEYINPUT122), .A3(G343), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT122), .B1(new_n1248), .B2(G343), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1248), .B1(new_n1249), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1255));
  AND4_X1   g1055(.A1(KEYINPUT121), .A2(new_n1255), .A3(new_n1243), .A4(new_n1249), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1254), .B1(new_n1256), .B2(new_n1244), .ZN(G409));
  NAND3_X1  g1057(.A1(G378), .A2(new_n1235), .A3(new_n1200), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1233), .A2(new_n1208), .A3(new_n1015), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1194), .A2(new_n725), .A3(new_n1196), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1186), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1236), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1258), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT60), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1212), .A2(new_n1265), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1111), .A2(new_n1107), .A3(KEYINPUT60), .A4(new_n1109), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1266), .A2(new_n685), .A3(new_n1121), .A4(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(G384), .B1(new_n1268), .B2(new_n1228), .ZN(new_n1269));
  OR2_X1    g1069(.A1(new_n1269), .A2(KEYINPUT124), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1228), .ZN(new_n1271));
  OR3_X1    g1071(.A1(new_n1271), .A2(KEYINPUT123), .A3(new_n842), .ZN(new_n1272));
  OAI21_X1  g1072(.A(KEYINPUT123), .B1(new_n1271), .B2(new_n842), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1269), .A2(KEYINPUT124), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1270), .A2(new_n1272), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1264), .A2(new_n1252), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  OR2_X1    g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(G393), .B(G396), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G390), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1007), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1086), .A2(new_n1282), .A3(new_n1087), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1284), .B(new_n1006), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1252), .A2(KEYINPUT125), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1253), .A2(G2897), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1276), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G2897), .B(new_n1253), .C1(new_n1275), .C2(new_n1286), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1264), .A2(new_n1252), .ZN(new_n1292));
  AOI21_X1  g1092(.A(KEYINPUT61), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1279), .A2(new_n1285), .A3(new_n1293), .A4(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT62), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1264), .A2(new_n1296), .A3(new_n1252), .A4(new_n1276), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1277), .A2(KEYINPUT62), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1293), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1295), .B1(new_n1299), .B2(new_n1285), .ZN(G405));
  INV_X1    g1100(.A(new_n1153), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(new_n1301), .A2(new_n1123), .A3(new_n1302), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(G375), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1236), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1305), .B1(new_n1235), .B2(new_n1200), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1276), .B1(new_n1304), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(G375), .A2(new_n1236), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1308), .A2(new_n1258), .A3(new_n1275), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1307), .A2(KEYINPUT126), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(KEYINPUT127), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT127), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1307), .A2(KEYINPUT126), .A3(new_n1312), .A4(new_n1309), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT126), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1284), .B(new_n1017), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1314), .A2(new_n1319), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1311), .A2(new_n1317), .A3(new_n1318), .A4(new_n1313), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(G402));
endmodule


