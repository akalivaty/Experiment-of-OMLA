

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772;

  NAND2_X2 U377 ( .A1(n397), .A2(n396), .ZN(n395) );
  NOR2_X1 U378 ( .A1(n364), .A2(n593), .ZN(n386) );
  AND2_X2 U379 ( .A1(n394), .A2(n399), .ZN(n398) );
  INV_X2 U380 ( .A(n636), .ZN(n637) );
  XNOR2_X2 U381 ( .A(n612), .B(KEYINPUT1), .ZN(n685) );
  XNOR2_X2 U382 ( .A(n542), .B(KEYINPUT102), .ZN(n531) );
  XNOR2_X2 U383 ( .A(n432), .B(n431), .ZN(n542) );
  INV_X2 U384 ( .A(G953), .ZN(n760) );
  NOR2_X1 U385 ( .A1(n771), .A2(n730), .ZN(n604) );
  XNOR2_X1 U386 ( .A(n407), .B(KEYINPUT32), .ZN(n771) );
  INV_X1 U387 ( .A(n594), .ZN(n619) );
  XNOR2_X1 U388 ( .A(G113), .B(KEYINPUT3), .ZN(n367) );
  XNOR2_X1 U389 ( .A(G116), .B(G122), .ZN(n405) );
  XNOR2_X1 U390 ( .A(n386), .B(n385), .ZN(n769) );
  NAND2_X1 U391 ( .A1(n685), .A2(n686), .ZN(n617) );
  OR2_X1 U392 ( .A1(n555), .A2(n570), .ZN(n734) );
  XNOR2_X1 U393 ( .A(n367), .B(G119), .ZN(n471) );
  XNOR2_X1 U394 ( .A(n405), .B(G107), .ZN(n514) );
  XNOR2_X1 U395 ( .A(KEYINPUT66), .B(G101), .ZN(n481) );
  NOR2_X2 U396 ( .A1(G953), .A2(G237), .ZN(n498) );
  AND2_X1 U397 ( .A1(n403), .A2(n413), .ZN(n402) );
  AND2_X1 U398 ( .A1(n409), .A2(n650), .ZN(n408) );
  NAND2_X1 U399 ( .A1(n772), .A2(n410), .ZN(n409) );
  NOR2_X1 U400 ( .A1(n582), .A2(n617), .ZN(n583) );
  NOR2_X1 U401 ( .A1(n589), .A2(n588), .ZN(n591) );
  XNOR2_X1 U402 ( .A(n550), .B(n549), .ZN(n589) );
  BUF_X1 U403 ( .A(n746), .Z(n354) );
  NOR2_X2 U404 ( .A1(n653), .A2(G902), .ZN(n449) );
  XNOR2_X2 U405 ( .A(n757), .B(n424), .ZN(n463) );
  XNOR2_X2 U406 ( .A(n422), .B(n423), .ZN(n757) );
  NOR2_X1 U407 ( .A1(n769), .A2(KEYINPUT44), .ZN(n363) );
  NOR2_X1 U408 ( .A1(n411), .A2(n558), .ZN(n403) );
  INV_X1 U409 ( .A(n769), .ZN(n406) );
  NAND2_X1 U410 ( .A1(n361), .A2(n604), .ZN(n360) );
  INV_X1 U411 ( .A(KEYINPUT67), .ZN(n362) );
  INV_X1 U412 ( .A(KEYINPUT73), .ZN(n420) );
  XOR2_X1 U413 ( .A(G131), .B(G140), .Z(n493) );
  XNOR2_X1 U414 ( .A(n458), .B(KEYINPUT90), .ZN(n459) );
  INV_X1 U415 ( .A(G107), .ZN(n458) );
  XOR2_X1 U416 ( .A(G110), .B(G104), .Z(n473) );
  XNOR2_X1 U417 ( .A(n488), .B(n366), .ZN(n672) );
  NAND2_X1 U418 ( .A1(n633), .A2(n746), .ZN(n359) );
  INV_X1 U419 ( .A(KEYINPUT82), .ZN(n631) );
  XNOR2_X1 U420 ( .A(n575), .B(KEYINPUT109), .ZN(n545) );
  XNOR2_X1 U421 ( .A(n365), .B(KEYINPUT34), .ZN(n364) );
  OR2_X1 U422 ( .A1(n615), .A2(n700), .ZN(n365) );
  INV_X1 U423 ( .A(KEYINPUT46), .ZN(n400) );
  INV_X1 U424 ( .A(n649), .ZN(n412) );
  INV_X1 U425 ( .A(KEYINPUT83), .ZN(n410) );
  INV_X1 U426 ( .A(KEYINPUT18), .ZN(n373) );
  INV_X1 U427 ( .A(KEYINPUT77), .ZN(n374) );
  XNOR2_X1 U428 ( .A(KEYINPUT12), .B(KEYINPUT95), .ZN(n496) );
  XNOR2_X1 U429 ( .A(KEYINPUT11), .B(KEYINPUT96), .ZN(n495) );
  XOR2_X1 U430 ( .A(G122), .B(G104), .Z(n502) );
  XNOR2_X1 U431 ( .A(G113), .B(G143), .ZN(n501) );
  NAND2_X1 U432 ( .A1(G234), .A2(G237), .ZN(n452) );
  XNOR2_X1 U433 ( .A(n492), .B(KEYINPUT38), .ZN(n705) );
  INV_X1 U434 ( .A(KEYINPUT15), .ZN(n445) );
  XNOR2_X1 U435 ( .A(G902), .B(KEYINPUT87), .ZN(n446) );
  INV_X1 U436 ( .A(G237), .ZN(n433) );
  XNOR2_X1 U437 ( .A(n509), .B(n508), .ZN(n569) );
  INV_X1 U438 ( .A(G902), .ZN(n517) );
  XNOR2_X1 U439 ( .A(G119), .B(G128), .ZN(n435) );
  XNOR2_X1 U440 ( .A(G137), .B(KEYINPUT23), .ZN(n437) );
  XOR2_X1 U441 ( .A(G146), .B(G125), .Z(n443) );
  INV_X1 U442 ( .A(G134), .ZN(n416) );
  XNOR2_X1 U443 ( .A(n360), .B(KEYINPUT70), .ZN(n628) );
  XNOR2_X1 U444 ( .A(n475), .B(n474), .ZN(n366) );
  XNOR2_X1 U445 ( .A(KEYINPUT72), .B(KEYINPUT16), .ZN(n472) );
  XNOR2_X1 U446 ( .A(n462), .B(n461), .ZN(n464) );
  XNOR2_X1 U447 ( .A(n460), .B(n459), .ZN(n461) );
  AND2_X1 U448 ( .A1(n548), .A2(n685), .ZN(n744) );
  INV_X1 U449 ( .A(KEYINPUT35), .ZN(n385) );
  AND2_X1 U450 ( .A1(n607), .A2(n603), .ZN(n407) );
  XOR2_X1 U451 ( .A(KEYINPUT24), .B(KEYINPUT91), .Z(n355) );
  NOR2_X1 U452 ( .A1(n555), .A2(n570), .ZN(n738) );
  AND2_X1 U453 ( .A1(n580), .A2(KEYINPUT83), .ZN(n356) );
  XOR2_X1 U454 ( .A(n383), .B(n643), .Z(n357) );
  XNOR2_X1 U455 ( .A(KEYINPUT122), .B(n638), .ZN(n358) );
  NOR2_X1 U456 ( .A1(n760), .A2(G952), .ZN(n675) );
  NAND2_X1 U457 ( .A1(n359), .A2(n635), .ZN(n636) );
  NAND2_X1 U458 ( .A1(n683), .A2(n359), .ZN(n721) );
  XNOR2_X1 U459 ( .A(n363), .B(n362), .ZN(n361) );
  XNOR2_X1 U460 ( .A(n366), .B(G101), .ZN(n753) );
  NAND2_X1 U461 ( .A1(n418), .A2(n417), .ZN(n368) );
  NAND2_X1 U462 ( .A1(n418), .A2(n417), .ZN(n371) );
  AND2_X1 U463 ( .A1(n392), .A2(n390), .ZN(n369) );
  NAND2_X1 U464 ( .A1(n391), .A2(n356), .ZN(n390) );
  NAND2_X1 U465 ( .A1(n573), .A2(n705), .ZN(n415) );
  XNOR2_X1 U466 ( .A(n470), .B(n469), .ZN(n573) );
  NAND2_X1 U467 ( .A1(n398), .A2(n395), .ZN(n370) );
  NAND2_X1 U468 ( .A1(n398), .A2(n395), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n672), .B(n671), .ZN(n673) );
  NOR2_X1 U470 ( .A1(n600), .A2(n601), .ZN(n607) );
  NAND2_X1 U471 ( .A1(n370), .A2(n402), .ZN(n372) );
  NAND2_X1 U472 ( .A1(n404), .A2(n402), .ZN(n401) );
  NAND2_X1 U473 ( .A1(KEYINPUT18), .A2(n374), .ZN(n375) );
  NAND2_X1 U474 ( .A1(n373), .A2(KEYINPUT77), .ZN(n376) );
  NAND2_X1 U475 ( .A1(n375), .A2(n376), .ZN(n478) );
  BUF_X1 U476 ( .A(n680), .Z(n759) );
  XNOR2_X1 U477 ( .A(n514), .B(n471), .ZN(n475) );
  BUF_X1 U478 ( .A(n521), .Z(n377) );
  BUF_X1 U479 ( .A(n542), .Z(n616) );
  XNOR2_X1 U480 ( .A(n657), .B(n656), .ZN(n658) );
  AND2_X1 U481 ( .A1(n555), .A2(n570), .ZN(n740) );
  NOR2_X1 U482 ( .A1(G902), .A2(n657), .ZN(n509) );
  NOR2_X2 U483 ( .A1(n531), .A2(n527), .ZN(n434) );
  XNOR2_X2 U484 ( .A(n449), .B(n378), .ZN(n606) );
  XNOR2_X1 U485 ( .A(KEYINPUT25), .B(n448), .ZN(n378) );
  BUF_X1 U486 ( .A(n757), .Z(n379) );
  XNOR2_X1 U487 ( .A(n372), .B(KEYINPUT48), .ZN(n380) );
  INV_X1 U488 ( .A(n397), .ZN(n381) );
  XNOR2_X1 U489 ( .A(G143), .B(G128), .ZN(n382) );
  BUF_X1 U490 ( .A(n644), .Z(n383) );
  XNOR2_X1 U491 ( .A(n401), .B(KEYINPUT48), .ZN(n393) );
  XNOR2_X1 U492 ( .A(n524), .B(n523), .ZN(n651) );
  NAND2_X1 U493 ( .A1(n384), .A2(n628), .ZN(n629) );
  XNOR2_X1 U494 ( .A(n627), .B(KEYINPUT85), .ZN(n384) );
  INV_X1 U495 ( .A(KEYINPUT2), .ZN(n417) );
  XNOR2_X1 U496 ( .A(n463), .B(n464), .ZN(n666) );
  XNOR2_X2 U497 ( .A(KEYINPUT99), .B(n556), .ZN(n702) );
  AND2_X2 U498 ( .A1(n637), .A2(n368), .ZN(n663) );
  NAND2_X1 U499 ( .A1(n387), .A2(n637), .ZN(n659) );
  AND2_X1 U500 ( .A1(n371), .A2(G475), .ZN(n387) );
  NAND2_X1 U501 ( .A1(n388), .A2(n637), .ZN(n674) );
  AND2_X1 U502 ( .A1(n371), .A2(G210), .ZN(n388) );
  NAND2_X1 U503 ( .A1(n663), .A2(G478), .ZN(n639) );
  NAND2_X1 U504 ( .A1(n663), .A2(G472), .ZN(n645) );
  AND2_X2 U505 ( .A1(n389), .A2(n408), .ZN(n392) );
  NAND2_X1 U506 ( .A1(n393), .A2(n410), .ZN(n389) );
  NAND2_X2 U507 ( .A1(n392), .A2(n390), .ZN(n630) );
  INV_X1 U508 ( .A(n380), .ZN(n391) );
  NAND2_X1 U509 ( .A1(n651), .A2(n400), .ZN(n394) );
  NOR2_X1 U510 ( .A1(n652), .A2(n400), .ZN(n396) );
  INV_X1 U511 ( .A(n651), .ZN(n397) );
  NAND2_X1 U512 ( .A1(n652), .A2(n400), .ZN(n399) );
  NAND2_X1 U513 ( .A1(n577), .A2(n701), .ZN(n550) );
  XNOR2_X2 U514 ( .A(n491), .B(n490), .ZN(n577) );
  NAND2_X1 U515 ( .A1(n604), .A2(n406), .ZN(n605) );
  NAND2_X1 U516 ( .A1(n568), .A2(n412), .ZN(n411) );
  INV_X1 U517 ( .A(n744), .ZN(n413) );
  INV_X1 U518 ( .A(n601), .ZN(n582) );
  NAND2_X1 U519 ( .A1(n414), .A2(n601), .ZN(n575) );
  NOR2_X1 U520 ( .A1(n544), .A2(n734), .ZN(n414) );
  INV_X1 U521 ( .A(n377), .ZN(n581) );
  XNOR2_X2 U522 ( .A(n415), .B(KEYINPUT39), .ZN(n521) );
  INV_X1 U523 ( .A(n423), .ZN(n513) );
  XNOR2_X2 U524 ( .A(n477), .B(n416), .ZN(n423) );
  XNOR2_X2 U525 ( .A(G143), .B(G128), .ZN(n477) );
  NAND2_X1 U526 ( .A1(n419), .A2(n746), .ZN(n418) );
  XNOR2_X2 U527 ( .A(n629), .B(KEYINPUT45), .ZN(n746) );
  XNOR2_X1 U528 ( .A(n680), .B(n420), .ZN(n419) );
  XNOR2_X2 U529 ( .A(n630), .B(KEYINPUT81), .ZN(n680) );
  OR2_X1 U530 ( .A1(n455), .A2(G900), .ZN(n421) );
  XNOR2_X1 U531 ( .A(n500), .B(n499), .ZN(n504) );
  INV_X1 U532 ( .A(G475), .ZN(n506) );
  XNOR2_X1 U533 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U534 ( .A(n507), .B(n506), .ZN(n508) );
  AND2_X1 U535 ( .A1(n510), .A2(G221), .ZN(n441) );
  XNOR2_X1 U536 ( .A(n632), .B(n631), .ZN(n633) );
  BUF_X1 U537 ( .A(n594), .Z(n615) );
  INV_X1 U538 ( .A(n675), .ZN(n646) );
  XNOR2_X1 U539 ( .A(n645), .B(n357), .ZN(n647) );
  XNOR2_X2 U540 ( .A(KEYINPUT69), .B(KEYINPUT4), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(G137), .ZN(n422) );
  XNOR2_X1 U542 ( .A(n481), .B(G146), .ZN(n424) );
  NAND2_X1 U543 ( .A1(n498), .A2(G210), .ZN(n425) );
  XNOR2_X1 U544 ( .A(n425), .B(G131), .ZN(n427) );
  XNOR2_X1 U545 ( .A(G116), .B(KEYINPUT5), .ZN(n426) );
  XNOR2_X1 U546 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U547 ( .A(n428), .B(n471), .ZN(n429) );
  XNOR2_X1 U548 ( .A(n463), .B(n429), .ZN(n644) );
  OR2_X2 U549 ( .A1(n644), .A2(G902), .ZN(n432) );
  XNOR2_X1 U550 ( .A(KEYINPUT92), .B(G472), .ZN(n430) );
  XNOR2_X1 U551 ( .A(n430), .B(KEYINPUT71), .ZN(n431) );
  NAND2_X1 U552 ( .A1(n517), .A2(n433), .ZN(n489) );
  NAND2_X1 U553 ( .A1(n489), .A2(G214), .ZN(n701) );
  INV_X1 U554 ( .A(n701), .ZN(n527) );
  XNOR2_X1 U555 ( .A(n434), .B(KEYINPUT30), .ZN(n468) );
  XOR2_X1 U556 ( .A(G140), .B(G110), .Z(n436) );
  XNOR2_X1 U557 ( .A(n436), .B(n435), .ZN(n439) );
  XNOR2_X1 U558 ( .A(n355), .B(n437), .ZN(n438) );
  XOR2_X1 U559 ( .A(n439), .B(n438), .Z(n442) );
  NAND2_X1 U560 ( .A1(G234), .A2(n760), .ZN(n440) );
  XOR2_X1 U561 ( .A(KEYINPUT8), .B(n440), .Z(n510) );
  XNOR2_X1 U562 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U563 ( .A(n443), .B(KEYINPUT10), .ZN(n494) );
  XNOR2_X1 U564 ( .A(n444), .B(n494), .ZN(n653) );
  XNOR2_X1 U565 ( .A(n446), .B(n445), .ZN(n634) );
  NAND2_X1 U566 ( .A1(G234), .A2(n634), .ZN(n447) );
  XNOR2_X1 U567 ( .A(KEYINPUT20), .B(n447), .ZN(n450) );
  NAND2_X1 U568 ( .A1(n450), .A2(G217), .ZN(n448) );
  NAND2_X1 U569 ( .A1(n450), .A2(G221), .ZN(n451) );
  XNOR2_X1 U570 ( .A(n451), .B(KEYINPUT21), .ZN(n688) );
  INV_X1 U571 ( .A(n688), .ZN(n533) );
  NAND2_X1 U572 ( .A1(n606), .A2(n533), .ZN(n611) );
  XNOR2_X1 U573 ( .A(n452), .B(KEYINPUT88), .ZN(n453) );
  XNOR2_X1 U574 ( .A(KEYINPUT14), .B(n453), .ZN(n454) );
  NAND2_X1 U575 ( .A1(G952), .A2(n454), .ZN(n713) );
  NOR2_X1 U576 ( .A1(n713), .A2(G953), .ZN(n587) );
  INV_X1 U577 ( .A(n587), .ZN(n456) );
  NAND2_X1 U578 ( .A1(G902), .A2(n454), .ZN(n585) );
  OR2_X1 U579 ( .A1(n760), .A2(n585), .ZN(n455) );
  NAND2_X1 U580 ( .A1(n456), .A2(n421), .ZN(n532) );
  INV_X1 U581 ( .A(n532), .ZN(n457) );
  NOR2_X1 U582 ( .A1(n611), .A2(n457), .ZN(n466) );
  XOR2_X1 U583 ( .A(n473), .B(n493), .Z(n462) );
  NAND2_X1 U584 ( .A1(G227), .A2(n760), .ZN(n460) );
  NAND2_X1 U585 ( .A1(n666), .A2(n517), .ZN(n465) );
  XNOR2_X2 U586 ( .A(n465), .B(G469), .ZN(n612) );
  AND2_X1 U587 ( .A1(n466), .A2(n612), .ZN(n467) );
  NAND2_X1 U588 ( .A1(n468), .A2(n467), .ZN(n470) );
  INV_X1 U589 ( .A(KEYINPUT74), .ZN(n469) );
  XNOR2_X1 U590 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U591 ( .A(G146), .B(G125), .ZN(n476) );
  XOR2_X1 U592 ( .A(n476), .B(KEYINPUT17), .Z(n480) );
  XNOR2_X1 U593 ( .A(n382), .B(n478), .ZN(n479) );
  XNOR2_X1 U594 ( .A(n480), .B(n479), .ZN(n487) );
  XNOR2_X1 U595 ( .A(n482), .B(n481), .ZN(n485) );
  NAND2_X1 U596 ( .A1(G224), .A2(n760), .ZN(n483) );
  XNOR2_X1 U597 ( .A(n483), .B(KEYINPUT76), .ZN(n484) );
  XNOR2_X1 U598 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U599 ( .A(n487), .B(n486), .ZN(n488) );
  NAND2_X1 U600 ( .A1(n672), .A2(n634), .ZN(n491) );
  AND2_X1 U601 ( .A1(n489), .A2(G210), .ZN(n490) );
  INV_X1 U602 ( .A(n577), .ZN(n492) );
  XNOR2_X1 U603 ( .A(n494), .B(n493), .ZN(n756) );
  INV_X1 U604 ( .A(n495), .ZN(n497) );
  XNOR2_X1 U605 ( .A(n497), .B(n496), .ZN(n500) );
  NAND2_X1 U606 ( .A1(n498), .A2(G214), .ZN(n499) );
  XNOR2_X1 U607 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U608 ( .A(n756), .B(n505), .ZN(n657) );
  INV_X1 U609 ( .A(KEYINPUT13), .ZN(n507) );
  XNOR2_X1 U610 ( .A(n569), .B(KEYINPUT97), .ZN(n555) );
  XOR2_X1 U611 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n512) );
  NAND2_X1 U612 ( .A1(G217), .A2(n510), .ZN(n511) );
  XNOR2_X1 U613 ( .A(n512), .B(n511), .ZN(n516) );
  XNOR2_X1 U614 ( .A(n513), .B(n514), .ZN(n515) );
  XNOR2_X1 U615 ( .A(n516), .B(n515), .ZN(n638) );
  NAND2_X1 U616 ( .A1(n638), .A2(n517), .ZN(n519) );
  XNOR2_X1 U617 ( .A(KEYINPUT98), .B(G478), .ZN(n518) );
  XNOR2_X1 U618 ( .A(n519), .B(n518), .ZN(n570) );
  INV_X1 U619 ( .A(n734), .ZN(n520) );
  NAND2_X1 U620 ( .A1(n521), .A2(n520), .ZN(n524) );
  INV_X1 U621 ( .A(KEYINPUT106), .ZN(n522) );
  XNOR2_X1 U622 ( .A(n522), .B(KEYINPUT40), .ZN(n523) );
  INV_X1 U623 ( .A(n569), .ZN(n526) );
  INV_X1 U624 ( .A(n570), .ZN(n525) );
  NAND2_X1 U625 ( .A1(n526), .A2(n525), .ZN(n703) );
  OR2_X1 U626 ( .A1(n703), .A2(n527), .ZN(n707) );
  INV_X1 U627 ( .A(n705), .ZN(n528) );
  NOR2_X1 U628 ( .A1(n707), .A2(n528), .ZN(n530) );
  INV_X1 U629 ( .A(KEYINPUT41), .ZN(n529) );
  XNOR2_X1 U630 ( .A(n530), .B(n529), .ZN(n715) );
  INV_X1 U631 ( .A(n531), .ZN(n597) );
  NAND2_X1 U632 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U633 ( .A1(n606), .A2(n534), .ZN(n541) );
  NAND2_X1 U634 ( .A1(n597), .A2(n541), .ZN(n536) );
  XNOR2_X1 U635 ( .A(KEYINPUT105), .B(KEYINPUT28), .ZN(n535) );
  XNOR2_X1 U636 ( .A(n536), .B(n535), .ZN(n537) );
  AND2_X1 U637 ( .A1(n537), .A2(n612), .ZN(n552) );
  NAND2_X1 U638 ( .A1(n715), .A2(n552), .ZN(n540) );
  XNOR2_X1 U639 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n538) );
  XNOR2_X1 U640 ( .A(n538), .B(KEYINPUT107), .ZN(n539) );
  XNOR2_X1 U641 ( .A(n540), .B(n539), .ZN(n652) );
  INV_X1 U642 ( .A(n541), .ZN(n544) );
  XNOR2_X1 U643 ( .A(KEYINPUT100), .B(KEYINPUT6), .ZN(n543) );
  XNOR2_X1 U644 ( .A(n616), .B(n543), .ZN(n601) );
  INV_X1 U645 ( .A(n545), .ZN(n546) );
  NOR2_X1 U646 ( .A1(n546), .A2(n550), .ZN(n547) );
  XNOR2_X1 U647 ( .A(n547), .B(KEYINPUT36), .ZN(n548) );
  XNOR2_X1 U648 ( .A(KEYINPUT75), .B(KEYINPUT19), .ZN(n549) );
  INV_X1 U649 ( .A(n589), .ZN(n551) );
  NAND2_X1 U650 ( .A1(n552), .A2(n551), .ZN(n735) );
  NOR2_X1 U651 ( .A1(n735), .A2(KEYINPUT47), .ZN(n553) );
  NAND2_X1 U652 ( .A1(KEYINPUT68), .A2(n553), .ZN(n554) );
  NAND2_X1 U653 ( .A1(n554), .A2(KEYINPUT80), .ZN(n557) );
  NOR2_X1 U654 ( .A1(n740), .A2(n738), .ZN(n556) );
  AND2_X1 U655 ( .A1(n557), .A2(n702), .ZN(n558) );
  INV_X1 U656 ( .A(KEYINPUT68), .ZN(n559) );
  AND2_X1 U657 ( .A1(n702), .A2(n559), .ZN(n561) );
  INV_X1 U658 ( .A(KEYINPUT47), .ZN(n560) );
  NOR2_X1 U659 ( .A1(n561), .A2(n560), .ZN(n565) );
  INV_X1 U660 ( .A(KEYINPUT80), .ZN(n562) );
  NOR2_X1 U661 ( .A1(n702), .A2(n562), .ZN(n563) );
  NOR2_X1 U662 ( .A1(n563), .A2(n735), .ZN(n564) );
  NAND2_X1 U663 ( .A1(n565), .A2(n564), .ZN(n567) );
  NAND2_X1 U664 ( .A1(n560), .A2(KEYINPUT80), .ZN(n566) );
  NAND2_X1 U665 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U666 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U667 ( .A(n571), .B(KEYINPUT103), .ZN(n592) );
  AND2_X1 U668 ( .A1(n577), .A2(n592), .ZN(n572) );
  AND2_X1 U669 ( .A1(n573), .A2(n572), .ZN(n649) );
  INV_X1 U670 ( .A(n685), .ZN(n608) );
  NAND2_X1 U671 ( .A1(n608), .A2(n701), .ZN(n574) );
  NOR2_X1 U672 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U673 ( .A(n576), .B(KEYINPUT43), .ZN(n578) );
  NOR2_X1 U674 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U675 ( .A(n579), .B(KEYINPUT104), .ZN(n772) );
  INV_X1 U676 ( .A(n772), .ZN(n580) );
  INV_X1 U677 ( .A(n740), .ZN(n731) );
  OR2_X1 U678 ( .A1(n581), .A2(n731), .ZN(n650) );
  INV_X1 U679 ( .A(n611), .ZN(n686) );
  XNOR2_X1 U680 ( .A(KEYINPUT33), .B(n583), .ZN(n700) );
  NOR2_X1 U681 ( .A1(G898), .A2(n760), .ZN(n584) );
  XNOR2_X1 U682 ( .A(KEYINPUT89), .B(n584), .ZN(n752) );
  NOR2_X1 U683 ( .A1(n585), .A2(n752), .ZN(n586) );
  NOR2_X1 U684 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U685 ( .A(KEYINPUT0), .B(KEYINPUT86), .Z(n590) );
  XNOR2_X1 U686 ( .A(n591), .B(n590), .ZN(n594) );
  XOR2_X1 U687 ( .A(n592), .B(KEYINPUT78), .Z(n593) );
  NOR2_X1 U688 ( .A1(n703), .A2(n688), .ZN(n595) );
  NAND2_X1 U689 ( .A1(n619), .A2(n595), .ZN(n596) );
  XNOR2_X1 U690 ( .A(n596), .B(KEYINPUT22), .ZN(n600) );
  NOR2_X1 U691 ( .A1(n597), .A2(n606), .ZN(n598) );
  NAND2_X1 U692 ( .A1(n608), .A2(n598), .ZN(n599) );
  NOR2_X1 U693 ( .A1(n600), .A2(n599), .ZN(n730) );
  INV_X1 U694 ( .A(n606), .ZN(n602) );
  AND2_X1 U695 ( .A1(n685), .A2(n602), .ZN(n603) );
  NAND2_X1 U696 ( .A1(n605), .A2(KEYINPUT44), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n607), .A2(n608), .ZN(n609) );
  NOR2_X1 U698 ( .A1(n602), .A2(n609), .ZN(n610) );
  XOR2_X1 U699 ( .A(KEYINPUT101), .B(n610), .Z(n770) );
  INV_X1 U700 ( .A(n702), .ZN(n623) );
  INV_X1 U701 ( .A(n616), .ZN(n693) );
  NOR2_X1 U702 ( .A1(n611), .A2(n693), .ZN(n613) );
  NAND2_X1 U703 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U704 ( .A1(n615), .A2(n614), .ZN(n725) );
  NOR2_X1 U705 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U706 ( .A(KEYINPUT93), .B(n618), .Z(n696) );
  NAND2_X1 U707 ( .A1(n696), .A2(n619), .ZN(n620) );
  XNOR2_X1 U708 ( .A(n620), .B(KEYINPUT94), .ZN(n621) );
  XNOR2_X1 U709 ( .A(KEYINPUT31), .B(n621), .ZN(n741) );
  NOR2_X1 U710 ( .A1(n725), .A2(n741), .ZN(n622) );
  NOR2_X1 U711 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U712 ( .A1(n770), .A2(n624), .ZN(n625) );
  NAND2_X1 U713 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U714 ( .A1(n369), .A2(KEYINPUT2), .ZN(n632) );
  INV_X1 U715 ( .A(n634), .ZN(n635) );
  XNOR2_X1 U716 ( .A(n639), .B(n358), .ZN(n640) );
  NAND2_X1 U717 ( .A1(n640), .A2(n646), .ZN(n641) );
  XNOR2_X1 U718 ( .A(n641), .B(KEYINPUT123), .ZN(G63) );
  XOR2_X1 U719 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n642) );
  XNOR2_X1 U720 ( .A(n642), .B(KEYINPUT62), .ZN(n643) );
  NAND2_X1 U721 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U722 ( .A(n648), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U723 ( .A(n649), .B(G143), .Z(G45) );
  XNOR2_X1 U724 ( .A(n650), .B(G134), .ZN(G36) );
  XOR2_X1 U725 ( .A(n381), .B(G131), .Z(G33) );
  XOR2_X1 U726 ( .A(G137), .B(n652), .Z(G39) );
  NAND2_X1 U727 ( .A1(n663), .A2(G217), .ZN(n654) );
  XNOR2_X1 U728 ( .A(n654), .B(n653), .ZN(n655) );
  NOR2_X1 U729 ( .A1(n655), .A2(n675), .ZN(G66) );
  XOR2_X1 U730 ( .A(KEYINPUT64), .B(KEYINPUT59), .Z(n656) );
  XNOR2_X1 U731 ( .A(n659), .B(n658), .ZN(n660) );
  NOR2_X2 U732 ( .A1(n660), .A2(n675), .ZN(n662) );
  XOR2_X1 U733 ( .A(KEYINPUT65), .B(KEYINPUT60), .Z(n661) );
  XNOR2_X1 U734 ( .A(n662), .B(n661), .ZN(G60) );
  NAND2_X1 U735 ( .A1(n663), .A2(G469), .ZN(n668) );
  XOR2_X1 U736 ( .A(KEYINPUT121), .B(KEYINPUT57), .Z(n664) );
  XNOR2_X1 U737 ( .A(n664), .B(KEYINPUT58), .ZN(n665) );
  XNOR2_X1 U738 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U739 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X1 U740 ( .A1(n669), .A2(n675), .ZN(G54) );
  XOR2_X1 U741 ( .A(KEYINPUT119), .B(KEYINPUT54), .Z(n670) );
  XNOR2_X1 U742 ( .A(n670), .B(KEYINPUT55), .ZN(n671) );
  XNOR2_X1 U743 ( .A(n674), .B(n673), .ZN(n676) );
  NOR2_X2 U744 ( .A1(n676), .A2(n675), .ZN(n679) );
  XNOR2_X1 U745 ( .A(KEYINPUT120), .B(KEYINPUT56), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n677), .B(KEYINPUT84), .ZN(n678) );
  XNOR2_X1 U747 ( .A(n679), .B(n678), .ZN(G51) );
  NAND2_X1 U748 ( .A1(n746), .A2(n759), .ZN(n681) );
  NAND2_X1 U749 ( .A1(n681), .A2(n417), .ZN(n682) );
  XOR2_X1 U750 ( .A(KEYINPUT79), .B(n682), .Z(n683) );
  XNOR2_X1 U751 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n684) );
  XNOR2_X1 U752 ( .A(n684), .B(KEYINPUT51), .ZN(n698) );
  NOR2_X1 U753 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U754 ( .A(KEYINPUT50), .B(n687), .Z(n692) );
  NAND2_X1 U755 ( .A1(n688), .A2(n602), .ZN(n689) );
  XNOR2_X1 U756 ( .A(n689), .B(KEYINPUT115), .ZN(n690) );
  XNOR2_X1 U757 ( .A(KEYINPUT49), .B(n690), .ZN(n691) );
  NAND2_X1 U758 ( .A1(n692), .A2(n691), .ZN(n694) );
  NOR2_X1 U759 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U760 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U761 ( .A(n698), .B(n697), .Z(n699) );
  NAND2_X1 U762 ( .A1(n699), .A2(n715), .ZN(n711) );
  INV_X1 U763 ( .A(n700), .ZN(n716) );
  NAND2_X1 U764 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U765 ( .A1(n704), .A2(n703), .ZN(n706) );
  NAND2_X1 U766 ( .A1(n706), .A2(n705), .ZN(n708) );
  NAND2_X1 U767 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U768 ( .A1(n716), .A2(n709), .ZN(n710) );
  NAND2_X1 U769 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U770 ( .A(KEYINPUT52), .B(n712), .Z(n714) );
  NOR2_X1 U771 ( .A1(n714), .A2(n713), .ZN(n719) );
  NAND2_X1 U772 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U773 ( .A1(n717), .A2(n760), .ZN(n718) );
  NOR2_X1 U774 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U775 ( .A1(n721), .A2(n720), .ZN(n723) );
  XOR2_X1 U776 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n722) );
  XNOR2_X1 U777 ( .A(n723), .B(n722), .ZN(G75) );
  NAND2_X1 U778 ( .A1(n725), .A2(n738), .ZN(n724) );
  XNOR2_X1 U779 ( .A(n724), .B(G104), .ZN(G6) );
  XNOR2_X1 U780 ( .A(G107), .B(KEYINPUT27), .ZN(n729) );
  XOR2_X1 U781 ( .A(KEYINPUT112), .B(KEYINPUT26), .Z(n727) );
  NAND2_X1 U782 ( .A1(n725), .A2(n740), .ZN(n726) );
  XNOR2_X1 U783 ( .A(n727), .B(n726), .ZN(n728) );
  XNOR2_X1 U784 ( .A(n729), .B(n728), .ZN(G9) );
  XOR2_X1 U785 ( .A(G110), .B(n730), .Z(G12) );
  NOR2_X1 U786 ( .A1(n735), .A2(n731), .ZN(n733) );
  XNOR2_X1 U787 ( .A(G128), .B(KEYINPUT29), .ZN(n732) );
  XNOR2_X1 U788 ( .A(n733), .B(n732), .ZN(G30) );
  NOR2_X1 U789 ( .A1(n735), .A2(n734), .ZN(n737) );
  XNOR2_X1 U790 ( .A(G146), .B(KEYINPUT113), .ZN(n736) );
  XNOR2_X1 U791 ( .A(n737), .B(n736), .ZN(G48) );
  NAND2_X1 U792 ( .A1(n741), .A2(n738), .ZN(n739) );
  XNOR2_X1 U793 ( .A(n739), .B(G113), .ZN(G15) );
  NAND2_X1 U794 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U795 ( .A(n742), .B(KEYINPUT114), .ZN(n743) );
  XNOR2_X1 U796 ( .A(G116), .B(n743), .ZN(G18) );
  XNOR2_X1 U797 ( .A(G125), .B(n744), .ZN(n745) );
  XNOR2_X1 U798 ( .A(n745), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U799 ( .A1(n354), .A2(n760), .ZN(n747) );
  XNOR2_X1 U800 ( .A(n747), .B(KEYINPUT124), .ZN(n751) );
  NAND2_X1 U801 ( .A1(G953), .A2(G224), .ZN(n748) );
  XNOR2_X1 U802 ( .A(KEYINPUT61), .B(n748), .ZN(n749) );
  NAND2_X1 U803 ( .A1(n749), .A2(G898), .ZN(n750) );
  NAND2_X1 U804 ( .A1(n751), .A2(n750), .ZN(n755) );
  NAND2_X1 U805 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U806 ( .A(n755), .B(n754), .Z(G69) );
  XOR2_X1 U807 ( .A(n379), .B(n756), .Z(n762) );
  XNOR2_X1 U808 ( .A(n762), .B(KEYINPUT125), .ZN(n758) );
  XNOR2_X1 U809 ( .A(n759), .B(n758), .ZN(n761) );
  NAND2_X1 U810 ( .A1(n761), .A2(n760), .ZN(n768) );
  XNOR2_X1 U811 ( .A(n762), .B(G227), .ZN(n763) );
  XNOR2_X1 U812 ( .A(n763), .B(KEYINPUT126), .ZN(n764) );
  NAND2_X1 U813 ( .A1(G900), .A2(n764), .ZN(n765) );
  XOR2_X1 U814 ( .A(KEYINPUT127), .B(n765), .Z(n766) );
  NAND2_X1 U815 ( .A1(G953), .A2(n766), .ZN(n767) );
  NAND2_X1 U816 ( .A1(n768), .A2(n767), .ZN(G72) );
  XOR2_X1 U817 ( .A(n769), .B(G122), .Z(G24) );
  XOR2_X1 U818 ( .A(G101), .B(n770), .Z(G3) );
  XOR2_X1 U819 ( .A(G119), .B(n771), .Z(G21) );
  XOR2_X1 U820 ( .A(G140), .B(n772), .Z(G42) );
endmodule

