//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1218, new_n1219,
    new_n1220, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291, new_n1292;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n204), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G68), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n206), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n209), .B(new_n214), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G226), .B(G232), .Z(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XOR2_X1   g0039(.A(G50), .B(G58), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  INV_X1    g0045(.A(KEYINPUT74), .ZN(new_n246));
  AND2_X1   g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NOR2_X1   g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g0049(.A(KEYINPUT7), .B1(new_n249), .B2(new_n204), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n253), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(G68), .B1(new_n250), .B2(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(G58), .A2(G68), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G58), .A2(G68), .ZN(new_n259));
  OAI21_X1  g0059(.A(G20), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G159), .ZN(new_n261));
  NOR4_X1   g0061(.A1(new_n261), .A2(KEYINPUT73), .A3(G20), .A4(G33), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT73), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G20), .A2(G33), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n263), .B1(new_n264), .B2(G159), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n260), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(KEYINPUT16), .B1(new_n257), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n212), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n253), .A2(new_n204), .A3(new_n254), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT7), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n224), .B1(new_n273), .B2(new_n255), .ZN(new_n274));
  OAI211_X1 g0074(.A(KEYINPUT16), .B(new_n260), .C1(new_n262), .C2(new_n265), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n270), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n246), .B1(new_n268), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n270), .ZN(new_n278));
  INV_X1    g0078(.A(new_n275), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n278), .B1(new_n257), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT16), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(new_n274), .B2(new_n266), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n280), .A2(KEYINPUT74), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n203), .A2(G20), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n278), .A2(new_n289), .ZN(new_n290));
  OAI22_X1  g0090(.A1(new_n288), .A2(new_n290), .B1(new_n289), .B2(new_n286), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G274), .ZN(new_n297));
  AND2_X1   g0097(.A1(G1), .A2(G13), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G41), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n296), .A2(G232), .B1(new_n295), .B2(new_n300), .ZN(new_n301));
  OR2_X1    g0101(.A1(G223), .A2(G1698), .ZN(new_n302));
  INV_X1    g0102(.A(G226), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G1698), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n302), .B(new_n304), .C1(new_n247), .C2(new_n248), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G87), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n293), .ZN(new_n308));
  AOI21_X1  g0108(.A(G200), .B1(new_n301), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n300), .A2(new_n295), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n298), .A2(new_n299), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n294), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n310), .B1(new_n223), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n311), .B1(new_n305), .B2(new_n306), .ZN(new_n314));
  INV_X1    g0114(.A(G190), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n315), .A2(KEYINPUT75), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(KEYINPUT75), .ZN(new_n317));
  OR2_X1    g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n313), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n309), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n284), .A2(new_n292), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT17), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n291), .B1(new_n277), .B2(new_n283), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT17), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(new_n325), .A3(new_n321), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G179), .ZN(new_n328));
  NOR3_X1   g0128(.A1(new_n313), .A2(new_n314), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n301), .A2(new_n308), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n329), .B1(new_n330), .B2(G169), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT18), .B1(new_n324), .B2(new_n331), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n268), .A2(new_n276), .A3(new_n246), .ZN(new_n333));
  AOI21_X1  g0133(.A(KEYINPUT74), .B1(new_n280), .B2(new_n282), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n292), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT18), .ZN(new_n336));
  INV_X1    g0136(.A(new_n331), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n327), .A2(new_n332), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n289), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n341), .A2(new_n270), .ZN(new_n342));
  INV_X1    g0142(.A(G50), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(new_n203), .B2(G20), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n342), .A2(new_n344), .B1(new_n343), .B2(new_n341), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n204), .A2(G33), .ZN(new_n346));
  INV_X1    g0146(.A(G150), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n204), .A2(new_n252), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n285), .A2(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT65), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n349), .A2(new_n350), .ZN(new_n352));
  NOR2_X1   g0152(.A1(G50), .A2(G58), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n204), .B1(new_n353), .B2(new_n224), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT66), .ZN(new_n355));
  NOR3_X1   g0155(.A1(new_n351), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n345), .B1(new_n356), .B2(new_n278), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n357), .B(KEYINPUT9), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n253), .A2(new_n254), .ZN(new_n359));
  INV_X1    g0159(.A(G1698), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G222), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G223), .A2(G1698), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n359), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(new_n293), .C1(G77), .C2(new_n359), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n364), .B(new_n310), .C1(new_n303), .C2(new_n312), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n365), .A2(new_n315), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(G200), .B2(new_n365), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n358), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n368), .B(KEYINPUT10), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n365), .A2(G179), .ZN(new_n370));
  INV_X1    g0170(.A(G169), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n370), .B1(new_n371), .B2(new_n365), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n357), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT69), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n290), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n342), .A2(KEYINPUT69), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n379), .A2(G68), .A3(new_n287), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT70), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT70), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n379), .A2(new_n382), .A3(G68), .A4(new_n287), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT71), .B1(new_n289), .B2(G68), .ZN(new_n385));
  XOR2_X1   g0185(.A(new_n385), .B(KEYINPUT12), .Z(new_n386));
  INV_X1    g0186(.A(KEYINPUT11), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n348), .A2(new_n343), .B1(new_n204), .B2(G68), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n346), .A2(new_n216), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n270), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n386), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(new_n387), .B2(new_n390), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n384), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT14), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n371), .A2(KEYINPUT72), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n223), .A2(G1698), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n359), .B(new_n396), .C1(G226), .C2(G1698), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G33), .A2(G97), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n311), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n310), .B1(new_n312), .B2(new_n225), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT13), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n399), .A2(KEYINPUT13), .A3(new_n400), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n394), .B(new_n395), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n403), .A2(new_n404), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n405), .B1(new_n407), .B2(new_n328), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n394), .B1(new_n407), .B2(new_n395), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n393), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n407), .A2(G200), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n406), .A2(G190), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n412), .A2(new_n384), .A3(new_n392), .A4(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n379), .A2(G77), .A3(new_n287), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(G77), .B2(new_n289), .ZN(new_n418));
  XNOR2_X1  g0218(.A(KEYINPUT15), .B(G87), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT67), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n420), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n421), .A2(new_n204), .A3(G33), .A4(new_n422), .ZN(new_n423));
  OR2_X1    g0223(.A1(new_n423), .A2(KEYINPUT68), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n285), .A2(new_n348), .B1(new_n204), .B2(new_n216), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n423), .B2(KEYINPUT68), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n278), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n418), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G238), .A2(G1698), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n359), .B(new_n429), .C1(new_n223), .C2(G1698), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n430), .B(new_n293), .C1(G107), .C2(new_n359), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n431), .B(new_n310), .C1(new_n217), .C2(new_n312), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n371), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(G179), .B2(new_n432), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n428), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n432), .A2(G200), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n315), .B2(new_n432), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n437), .A2(new_n427), .A3(new_n418), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  AND4_X1   g0239(.A1(new_n340), .A2(new_n375), .A3(new_n416), .A4(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G41), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n203), .B(G45), .C1(new_n442), .C2(KEYINPUT5), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n442), .A2(KEYINPUT5), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(new_n293), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G257), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n300), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G283), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n359), .A2(G250), .A3(G1698), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n217), .A2(G1698), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n359), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n451), .B(new_n452), .C1(new_n454), .C2(KEYINPUT4), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n359), .A2(KEYINPUT4), .A3(new_n453), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT77), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n454), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n455), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n450), .B1(new_n460), .B2(new_n311), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n371), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(new_n458), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n452), .A2(new_n451), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT4), .B1(new_n359), .B2(new_n453), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n449), .B1(new_n467), .B2(new_n293), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n328), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n462), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G97), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n341), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n203), .A2(G33), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n342), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n472), .B1(new_n474), .B2(new_n471), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT6), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n476), .A2(new_n471), .A3(G107), .ZN(new_n477));
  XNOR2_X1  g0277(.A(G97), .B(G107), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n477), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  OAI22_X1  g0279(.A1(new_n479), .A2(new_n204), .B1(new_n216), .B2(new_n348), .ZN(new_n480));
  INV_X1    g0280(.A(G107), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(new_n273), .B2(new_n255), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n270), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT76), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT76), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n485), .B(new_n270), .C1(new_n480), .C2(new_n482), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n475), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT78), .B1(new_n470), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n487), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT78), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n489), .A2(new_n490), .A3(new_n462), .A4(new_n469), .ZN(new_n491));
  XOR2_X1   g0291(.A(KEYINPUT79), .B(G87), .Z(new_n492));
  NOR2_X1   g0292(.A1(G97), .A2(G107), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n398), .A2(new_n204), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(KEYINPUT19), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n359), .A2(new_n204), .A3(G68), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n346), .A2(new_n471), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n496), .B(new_n497), .C1(KEYINPUT19), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n270), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n421), .A2(new_n422), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n341), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n474), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n503), .B1(G87), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n203), .A2(new_n297), .A3(G45), .ZN(new_n506));
  INV_X1    g0306(.A(G45), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n219), .B1(new_n507), .B2(G1), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n311), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(G116), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n252), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(G238), .A2(G1698), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n512), .B1(new_n217), .B2(G1698), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n511), .B1(new_n513), .B2(new_n359), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n509), .B1(new_n514), .B2(new_n311), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(new_n315), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n516), .B1(G200), .B2(new_n515), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n500), .B(new_n502), .C1(new_n501), .C2(new_n474), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n515), .A2(G179), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n519), .B1(new_n371), .B2(new_n515), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n505), .A2(new_n517), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n461), .A2(G200), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n487), .B(new_n522), .C1(new_n315), .C2(new_n461), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n488), .A2(new_n491), .A3(new_n521), .A4(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n451), .B(new_n204), .C1(G33), .C2(new_n471), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n510), .A2(G20), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(new_n270), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT20), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT81), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT81), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n528), .A2(new_n531), .A3(KEYINPUT20), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n530), .B(new_n532), .C1(KEYINPUT20), .C2(new_n528), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n341), .A2(new_n510), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n510), .B1(new_n203), .B2(G33), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n377), .A2(new_n378), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G264), .A2(G1698), .ZN(new_n538));
  INV_X1    g0338(.A(G257), .ZN(new_n539));
  OAI221_X1 g0339(.A(new_n538), .B1(new_n539), .B2(G1698), .C1(new_n247), .C2(new_n248), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n540), .B(new_n293), .C1(G303), .C2(new_n359), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n311), .B(G270), .C1(new_n443), .C2(new_n444), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n448), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT80), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n541), .A2(new_n448), .A3(KEYINPUT80), .A4(new_n542), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n537), .A2(new_n547), .A3(KEYINPUT21), .A4(G169), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n536), .A2(new_n534), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n528), .A2(KEYINPUT20), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(KEYINPUT81), .B2(new_n529), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n549), .B1(new_n551), .B2(new_n532), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n545), .A2(G200), .A3(new_n546), .ZN(new_n553));
  INV_X1    g0353(.A(new_n318), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n552), .B(new_n553), .C1(new_n547), .C2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n543), .A2(new_n328), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n537), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT21), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n545), .A2(G169), .A3(new_n546), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n552), .B2(new_n559), .ZN(new_n560));
  AND4_X1   g0360(.A1(new_n548), .A2(new_n555), .A3(new_n557), .A4(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n359), .A2(new_n204), .A3(G87), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n562), .B(KEYINPUT22), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT24), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT23), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n204), .B2(G107), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n481), .A2(KEYINPUT23), .A3(G20), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n566), .A2(new_n567), .B1(new_n511), .B2(new_n204), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n563), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n564), .B1(new_n563), .B2(new_n568), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n270), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n341), .A2(new_n481), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n572), .B(KEYINPUT25), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n504), .B2(G107), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n446), .A2(G264), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n359), .A2(G250), .A3(new_n360), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G294), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT82), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n539), .A2(new_n360), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n359), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n359), .A2(new_n581), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT82), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n579), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n448), .B(new_n576), .C1(new_n585), .C2(new_n311), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G200), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n584), .A2(new_n582), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n577), .A2(new_n578), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n590), .A2(new_n293), .B1(G264), .B2(new_n446), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(G190), .A3(new_n448), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n575), .A2(new_n587), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n571), .A2(new_n574), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n586), .A2(G169), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n590), .A2(new_n293), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n596), .A2(G179), .A3(new_n448), .A4(new_n576), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n595), .A2(KEYINPUT83), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT83), .B1(new_n595), .B2(new_n597), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n594), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n561), .A2(new_n593), .A3(new_n600), .ZN(new_n601));
  NOR3_X1   g0401(.A1(new_n441), .A2(new_n524), .A3(new_n601), .ZN(G372));
  AND4_X1   g0402(.A1(new_n325), .A2(new_n284), .A3(new_n292), .A4(new_n321), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n325), .B1(new_n324), .B2(new_n321), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n435), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n410), .B1(new_n415), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n605), .B1(new_n607), .B2(KEYINPUT84), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(KEYINPUT84), .B2(new_n607), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n338), .A2(new_n332), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n612), .A2(new_n369), .B1(new_n357), .B2(new_n372), .ZN(new_n613));
  INV_X1    g0413(.A(new_n593), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n560), .A2(new_n557), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n548), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n595), .A2(new_n597), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n594), .A2(new_n618), .ZN(new_n619));
  AOI211_X1 g0419(.A(new_n614), .B(new_n524), .C1(new_n617), .C2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n470), .A2(new_n487), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n621), .A2(new_n521), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n518), .A2(new_n520), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n488), .A2(new_n491), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n626), .A2(new_n521), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n624), .B(new_n625), .C1(new_n627), .C2(new_n623), .ZN(new_n628));
  OR2_X1    g0428(.A1(new_n620), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n613), .B1(new_n441), .B2(new_n630), .ZN(G369));
  NAND3_X1  g0431(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n633));
  XOR2_X1   g0433(.A(new_n633), .B(KEYINPUT85), .Z(new_n634));
  OAI21_X1  g0434(.A(G213), .B1(new_n632), .B2(KEYINPUT27), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(G343), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(new_n552), .ZN(new_n641));
  MUX2_X1   g0441(.A(new_n561), .B(new_n616), .S(new_n641), .Z(new_n642));
  XNOR2_X1  g0442(.A(KEYINPUT86), .B(G330), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g0444(.A(new_n644), .B(KEYINPUT87), .Z(new_n645));
  OAI211_X1 g0445(.A(new_n600), .B(new_n593), .C1(new_n575), .C2(new_n640), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(KEYINPUT88), .ZN(new_n647));
  INV_X1    g0447(.A(new_n600), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n647), .B1(new_n648), .B2(new_n639), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n617), .A2(new_n639), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n619), .B2(new_n639), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n650), .A2(new_n653), .ZN(G399));
  INV_X1    g0454(.A(new_n207), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(G41), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G1), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n492), .A2(new_n510), .A3(new_n493), .ZN(new_n659));
  OAI22_X1  g0459(.A1(new_n658), .A2(new_n659), .B1(new_n210), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT28), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n629), .A2(new_n640), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT29), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n625), .B1(new_n622), .B2(new_n623), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n665), .B1(new_n623), .B2(new_n627), .ZN(new_n666));
  AND4_X1   g0466(.A1(new_n488), .A2(new_n491), .A3(new_n523), .A4(new_n521), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n667), .B(new_n593), .C1(new_n616), .C2(new_n648), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n639), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT29), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n664), .A2(new_n670), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n561), .A2(new_n593), .A3(new_n600), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(new_n667), .A3(new_n640), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n515), .A2(new_n328), .ZN(new_n674));
  AND4_X1   g0474(.A1(new_n461), .A2(new_n547), .A3(new_n586), .A4(new_n674), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n543), .A2(new_n515), .A3(new_n328), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n591), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT30), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n677), .A2(new_n678), .A3(new_n461), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT90), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n677), .B2(new_n461), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n468), .A2(KEYINPUT90), .A3(new_n591), .A4(new_n676), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(new_n678), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g0485(.A(KEYINPUT89), .B(KEYINPUT31), .Z(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(new_n639), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT91), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n682), .A2(new_n683), .A3(KEYINPUT91), .A4(new_n678), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(new_n690), .A3(new_n680), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n691), .A2(new_n639), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(KEYINPUT31), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n673), .B(new_n687), .C1(new_n693), .C2(KEYINPUT92), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n693), .A2(KEYINPUT92), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n643), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n671), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n661), .B1(new_n697), .B2(G1), .ZN(G364));
  AND2_X1   g0498(.A1(new_n204), .A2(G13), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G45), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G1), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n656), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g0502(.A(new_n702), .B(KEYINPUT93), .Z(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n645), .B(new_n704), .C1(new_n643), .C2(new_n642), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n655), .A2(new_n249), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G355), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(G116), .B2(new_n207), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n655), .A2(new_n359), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n710), .B1(new_n507), .B2(new_n211), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n241), .A2(G45), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n708), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(G13), .A2(G33), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G20), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n212), .B1(G20), .B2(new_n371), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n703), .B1(new_n713), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n204), .A2(new_n328), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G200), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n554), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT95), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n204), .A2(G179), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(G190), .A3(G200), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT96), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n725), .A2(G326), .B1(G303), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT94), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n721), .B(new_n730), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n554), .A2(new_n731), .A3(G200), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(G322), .ZN(new_n734));
  INV_X1    g0534(.A(G311), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n731), .A2(G190), .A3(G200), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI22_X1  g0537(.A1(new_n733), .A2(new_n734), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n315), .A2(G179), .A3(G200), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n204), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n722), .A2(G190), .ZN(new_n742));
  XNOR2_X1  g0542(.A(KEYINPUT33), .B(G317), .ZN(new_n743));
  AOI22_X1  g0543(.A1(G294), .A2(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G190), .A2(G200), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n726), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n359), .B1(new_n747), .B2(G329), .ZN(new_n748));
  INV_X1    g0548(.A(G283), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n726), .A2(new_n315), .A3(G200), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n744), .B(new_n748), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n738), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n729), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT97), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n492), .A2(new_n727), .B1(new_n750), .B2(new_n481), .ZN(new_n755));
  INV_X1    g0555(.A(new_n742), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n224), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n755), .B(new_n757), .C1(G50), .C2(new_n723), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT32), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(new_n746), .B2(new_n261), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n747), .A2(KEYINPUT32), .A3(G159), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n736), .A2(G77), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n732), .A2(G58), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n249), .B1(new_n741), .B2(G97), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n758), .A2(new_n762), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(KEYINPUT98), .B1(new_n754), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n717), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n754), .A2(KEYINPUT98), .A3(new_n765), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n720), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n716), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n770), .B1(new_n642), .B2(new_n771), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n705), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(G396));
  AOI21_X1  g0574(.A(new_n249), .B1(new_n747), .B2(G132), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n775), .B1(new_n222), .B2(new_n740), .C1(new_n224), .C2(new_n750), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n723), .A2(G137), .B1(G150), .B2(new_n742), .ZN(new_n777));
  INV_X1    g0577(.A(G143), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n777), .B1(new_n737), .B2(new_n261), .C1(new_n733), .C2(new_n778), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT34), .Z(new_n780));
  AOI211_X1 g0580(.A(new_n776), .B(new_n780), .C1(G50), .C2(new_n728), .ZN(new_n781));
  INV_X1    g0581(.A(new_n750), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n723), .A2(G303), .B1(G87), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n249), .B1(new_n746), .B2(new_n735), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(G97), .B2(new_n741), .ZN(new_n785));
  INV_X1    g0585(.A(G294), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n783), .B(new_n785), .C1(new_n733), .C2(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n736), .A2(G116), .B1(G283), .B2(new_n742), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT100), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n787), .B(new_n789), .C1(G107), .C2(new_n728), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n717), .B1(new_n781), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n717), .A2(new_n714), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT99), .Z(new_n793));
  OAI211_X1 g0593(.A(new_n791), .B(new_n703), .C1(G77), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n428), .A2(new_n640), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n795), .A2(new_n438), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n606), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n606), .A2(new_n639), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n794), .B1(new_n714), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n662), .A2(new_n800), .ZN(new_n802));
  INV_X1    g0602(.A(new_n800), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n640), .B(new_n803), .C1(new_n620), .C2(new_n628), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n805), .A2(new_n696), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n703), .B1(new_n805), .B2(new_n696), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n801), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G384));
  INV_X1    g0609(.A(new_n479), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n810), .A2(KEYINPUT35), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(KEYINPUT35), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n811), .A2(G116), .A3(new_n213), .A4(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT36), .Z(new_n814));
  OAI211_X1 g0614(.A(new_n211), .B(G77), .C1(new_n222), .C2(new_n224), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n343), .A2(G68), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n203), .B(G13), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n640), .B1(new_n384), .B2(new_n392), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(KEYINPUT101), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n393), .A2(new_n639), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT101), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n410), .A2(new_n820), .A3(new_n414), .A4(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n819), .B1(new_n408), .B2(new_n409), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n804), .B2(new_n799), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT102), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n274), .B2(new_n266), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n257), .A2(KEYINPUT102), .A3(new_n267), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n829), .A2(new_n830), .A3(new_n281), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n291), .B1(new_n831), .B2(new_n280), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n832), .A2(new_n637), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n322), .B1(new_n331), .B2(new_n832), .ZN(new_n834));
  OAI21_X1  g0634(.A(KEYINPUT37), .B1(new_n834), .B2(new_n833), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n335), .A2(new_n337), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n335), .A2(new_n636), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT37), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n836), .A2(new_n837), .A3(new_n838), .A4(new_n322), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n339), .A2(new_n833), .B1(new_n835), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT103), .B1(new_n840), .B2(KEYINPUT38), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n833), .B1(new_n605), .B2(new_n610), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n291), .B(new_n320), .C1(new_n277), .C2(new_n283), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n831), .A2(new_n280), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n331), .B1(new_n844), .B2(new_n292), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n843), .A2(new_n833), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n839), .B1(new_n846), .B2(new_n838), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT38), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT103), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n842), .A2(new_n847), .A3(KEYINPUT38), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n841), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n827), .A2(new_n852), .B1(new_n610), .B2(new_n637), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n851), .B1(new_n848), .B2(new_n849), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n840), .A2(KEYINPUT103), .A3(KEYINPUT38), .ZN(new_n856));
  OAI211_X1 g0656(.A(KEYINPUT104), .B(KEYINPUT39), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT104), .B1(new_n852), .B2(KEYINPUT39), .ZN(new_n859));
  INV_X1    g0659(.A(new_n837), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n605), .B2(new_n610), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n836), .A2(new_n837), .A3(new_n322), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT37), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n861), .A2(KEYINPUT105), .B1(new_n839), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT105), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n339), .A2(new_n865), .A3(new_n860), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT38), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n842), .A2(new_n847), .A3(KEYINPUT38), .ZN(new_n868));
  NOR4_X1   g0668(.A1(new_n867), .A2(KEYINPUT106), .A3(KEYINPUT39), .A4(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT106), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n861), .A2(KEYINPUT105), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n863), .A2(new_n839), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n871), .A2(new_n866), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n868), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT39), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n870), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n858), .A2(new_n859), .B1(new_n869), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT107), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT39), .B1(new_n855), .B2(new_n856), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT104), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n857), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n873), .A2(new_n874), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(new_n876), .A3(new_n851), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(KEYINPUT106), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n875), .A2(new_n870), .A3(new_n876), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT107), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n883), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n879), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n411), .A2(new_n640), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n854), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT108), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n664), .A2(new_n440), .A3(new_n670), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n613), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n895), .B(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n691), .A2(KEYINPUT31), .A3(new_n639), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n673), .B(new_n899), .C1(new_n692), .C2(new_n686), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n826), .A2(new_n800), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT40), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n875), .A2(KEYINPUT109), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT109), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n867), .B2(new_n868), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n902), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n824), .A2(new_n825), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n803), .A2(new_n907), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n601), .A2(new_n524), .A3(new_n639), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n686), .B1(new_n691), .B2(new_n639), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n908), .B1(new_n911), .B2(new_n899), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT40), .B1(new_n912), .B2(new_n852), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n906), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(new_n440), .A3(new_n900), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(new_n852), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT40), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n903), .A2(new_n905), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n918), .B1(new_n919), .B2(new_n902), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n440), .A2(new_n900), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n915), .A2(new_n922), .A3(new_n643), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n898), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n203), .B2(new_n699), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n898), .A2(new_n923), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n818), .B1(new_n925), .B2(new_n926), .ZN(G367));
  INV_X1    g0727(.A(new_n626), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n928), .B(new_n523), .C1(new_n487), .C2(new_n640), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n621), .A2(new_n639), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n928), .B1(new_n932), .B2(new_n600), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n931), .A2(new_n647), .A3(new_n651), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n933), .A2(new_n640), .B1(KEYINPUT42), .B2(new_n934), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n934), .A2(KEYINPUT42), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n505), .A2(new_n640), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n521), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n625), .B2(new_n937), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n935), .A2(new_n936), .B1(KEYINPUT43), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n940), .B(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n650), .A2(new_n931), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n942), .B(new_n943), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n656), .B(KEYINPUT41), .Z(new_n945));
  NAND2_X1  g0745(.A1(new_n653), .A2(new_n932), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT44), .Z(new_n947));
  NOR2_X1   g0747(.A1(new_n653), .A2(new_n932), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT45), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n650), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n947), .B(new_n949), .C1(new_n645), .C2(new_n649), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n649), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n652), .B1(new_n954), .B2(new_n651), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(new_n645), .Z(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n697), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n945), .B1(new_n958), .B2(new_n697), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n701), .B(KEYINPUT110), .Z(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n944), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n718), .B1(new_n207), .B2(new_n501), .C1(new_n710), .C2(new_n237), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n703), .A2(new_n963), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n725), .A2(G311), .B1(G303), .B2(new_n732), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT111), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n736), .A2(G283), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n728), .A2(KEYINPUT46), .A3(G116), .ZN(new_n968));
  INV_X1    g0768(.A(G317), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n249), .B1(new_n746), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G97), .B2(new_n782), .ZN(new_n971));
  AOI22_X1  g0771(.A1(G107), .A2(new_n741), .B1(new_n742), .B2(G294), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n967), .A2(new_n968), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n727), .ZN(new_n974));
  AOI21_X1  g0774(.A(KEYINPUT46), .B1(new_n974), .B2(G116), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT112), .Z(new_n976));
  NOR2_X1   g0776(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n782), .A2(G77), .ZN(new_n978));
  INV_X1    g0778(.A(G137), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n978), .B(new_n359), .C1(new_n979), .C2(new_n746), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n737), .A2(new_n343), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n980), .B(new_n981), .C1(G150), .C2(new_n732), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n741), .A2(G68), .B1(new_n974), .B2(G58), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n261), .B2(new_n756), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(new_n725), .B2(G143), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n966), .A2(new_n977), .B1(new_n982), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT47), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n964), .B1(new_n771), .B2(new_n939), .C1(new_n987), .C2(new_n767), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n962), .A2(new_n988), .ZN(G387));
  AOI22_X1  g0789(.A1(new_n736), .A2(G303), .B1(G311), .B2(new_n742), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n969), .B2(new_n733), .C1(new_n724), .C2(new_n734), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT48), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n992), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n741), .A2(G283), .B1(new_n974), .B2(G294), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT49), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n997), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n750), .A2(new_n510), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n359), .B(new_n1000), .C1(G326), .C2(new_n747), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n421), .A2(new_n741), .A3(new_n422), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n737), .B2(new_n224), .C1(new_n733), .C2(new_n343), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n974), .A2(G77), .B1(new_n747), .B2(G150), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1005), .A2(KEYINPUT113), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n723), .A2(G159), .B1(new_n286), .B2(new_n742), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(KEYINPUT113), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n249), .B1(new_n782), .B2(G97), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  NOR3_X1   g0810(.A1(new_n1004), .A2(new_n1006), .A3(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT114), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n767), .B1(new_n1002), .B2(new_n1012), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n234), .A2(new_n507), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n1014), .A2(new_n709), .B1(new_n659), .B2(new_n706), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n286), .A2(new_n343), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT50), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n507), .B1(new_n224), .B2(new_n216), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n1017), .A2(new_n659), .A3(new_n1018), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n1015), .A2(new_n1019), .B1(G107), .B2(new_n207), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n704), .B(new_n1013), .C1(new_n718), .C2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT115), .Z(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n649), .B2(new_n716), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n956), .B2(new_n961), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n657), .B1(new_n956), .B2(new_n697), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n697), .B2(new_n956), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1026), .ZN(G393));
  INV_X1    g0827(.A(KEYINPUT116), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n960), .B1(new_n953), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n951), .A2(KEYINPUT116), .A3(new_n952), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n932), .A2(new_n716), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n732), .A2(G311), .B1(new_n723), .B2(G317), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT52), .Z(new_n1033));
  OAI221_X1 g0833(.A(new_n249), .B1(new_n746), .B2(new_n734), .C1(new_n481), .C2(new_n750), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G116), .A2(new_n741), .B1(new_n742), .B2(G303), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n749), .B2(new_n727), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1034), .B(new_n1036), .C1(G294), .C2(new_n736), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1033), .A2(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n732), .A2(G159), .B1(new_n723), .B2(G150), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT51), .Z(new_n1040));
  OAI221_X1 g0840(.A(new_n359), .B1(new_n746), .B2(new_n778), .C1(new_n218), .C2(new_n750), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n741), .A2(G77), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n224), .B2(new_n727), .C1(new_n756), .C2(new_n343), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1041), .B(new_n1043), .C1(new_n286), .C2(new_n736), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n767), .B1(new_n1038), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n710), .A2(new_n244), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n719), .B(new_n1047), .C1(G97), .C2(new_n655), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1046), .A2(new_n704), .A3(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1029), .A2(new_n1030), .B1(new_n1031), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n953), .A2(new_n957), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n958), .A2(new_n656), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1052), .ZN(G390));
  INV_X1    g0853(.A(KEYINPUT119), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n827), .A2(new_n893), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n879), .A2(new_n890), .A3(new_n1055), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n643), .B(new_n901), .C1(new_n694), .C2(new_n695), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n798), .B1(new_n669), .B2(new_n797), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n892), .B1(new_n1058), .B2(new_n826), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1059), .A2(new_n919), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  AND3_X1   g0861(.A1(new_n1056), .A2(new_n1057), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(G330), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n911), .B2(new_n899), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n901), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n1062), .A2(new_n1066), .A3(new_n960), .ZN(new_n1067));
  AND3_X1   g0867(.A1(new_n883), .A2(new_n888), .A3(new_n889), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n889), .B1(new_n883), .B2(new_n888), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n714), .ZN(new_n1071));
  OAI21_X1  g0871(.A(KEYINPUT53), .B1(new_n727), .B2(new_n347), .ZN(new_n1072));
  INV_X1    g0872(.A(G132), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1072), .B1(new_n733), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n723), .A2(G128), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n249), .B1(new_n747), .B2(G125), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(KEYINPUT54), .B(G143), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1075), .B(new_n1076), .C1(new_n737), .C2(new_n1077), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n727), .A2(KEYINPUT53), .A3(new_n347), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n741), .A2(G159), .B1(new_n782), .B2(G50), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n979), .B2(new_n756), .ZN(new_n1081));
  NOR4_X1   g0881(.A1(new_n1074), .A2(new_n1078), .A3(new_n1079), .A4(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n733), .A2(new_n510), .B1(new_n737), .B2(new_n471), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n750), .A2(new_n224), .B1(new_n746), .B2(new_n786), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G87), .A2(new_n728), .B1(new_n1085), .B2(KEYINPUT118), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(KEYINPUT118), .B2(new_n1085), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n723), .A2(G283), .B1(G107), .B2(new_n742), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1088), .A2(new_n249), .A3(new_n1042), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n1083), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n717), .B1(new_n1082), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n793), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n704), .B1(new_n285), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1071), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1054), .B1(new_n1067), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1056), .A2(new_n1057), .A3(new_n1061), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1060), .B1(new_n1070), .B2(new_n1055), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n961), .B(new_n1097), .C1(new_n1098), .C2(new_n1065), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1099), .A2(KEYINPUT119), .A3(new_n1094), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n440), .A2(new_n1064), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n896), .A2(new_n613), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n826), .B1(new_n696), .B2(new_n800), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1103), .A2(new_n1065), .B1(new_n799), .B2(new_n804), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT117), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1064), .A2(new_n803), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1106), .B1(new_n1107), .B2(new_n826), .ZN(new_n1108));
  AOI211_X1 g0908(.A(KEYINPUT117), .B(new_n907), .C1(new_n1064), .C2(new_n803), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n1105), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1102), .B1(new_n1104), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n896), .A2(new_n613), .A3(new_n1101), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1103), .A2(new_n1065), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n804), .A2(new_n799), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  OR3_X1    g0916(.A1(new_n1105), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1113), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1097), .B(new_n1118), .C1(new_n1098), .C2(new_n1065), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1112), .A2(new_n1119), .A3(new_n656), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1096), .A2(new_n1100), .A3(new_n1120), .ZN(G378));
  XNOR2_X1  g0921(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n369), .B2(new_n373), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n369), .A2(new_n373), .A3(new_n1123), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1125), .A2(new_n357), .A3(new_n636), .A4(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n357), .A2(new_n636), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1126), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1128), .B1(new_n1129), .B2(new_n1124), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n714), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n703), .B1(G50), .B2(new_n793), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n222), .A2(new_n750), .B1(new_n727), .B2(new_n216), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n756), .A2(new_n471), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1135), .B(new_n1136), .C1(G116), .C2(new_n723), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n359), .A2(G41), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1138), .B1(new_n749), .B2(new_n746), .C1(new_n224), .C2(new_n740), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n732), .B2(G107), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1137), .B(new_n1140), .C1(new_n501), .C2(new_n737), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT58), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1138), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1144), .B(new_n343), .C1(G33), .C2(G41), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n723), .A2(G125), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n742), .A2(G132), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1149), .B1(new_n347), .B2(new_n740), .C1(new_n727), .C2(new_n1077), .ZN(new_n1150));
  INV_X1    g0950(.A(G128), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n733), .A2(new_n1151), .B1(new_n737), .B2(new_n979), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(KEYINPUT59), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n782), .A2(G159), .ZN(new_n1156));
  AOI211_X1 g0956(.A(G33), .B(G41), .C1(new_n747), .C2(G124), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1154), .A2(KEYINPUT59), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1146), .B1(new_n1142), .B2(new_n1141), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1134), .B1(new_n1160), .B2(new_n717), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1133), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1131), .B1(new_n914), .B2(G330), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n906), .A2(new_n1132), .A3(new_n913), .A4(new_n1063), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT120), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n894), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1132), .B1(new_n920), .B2(new_n1063), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n914), .A2(G330), .A3(new_n1131), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n892), .B1(new_n879), .B2(new_n890), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1170), .B(KEYINPUT120), .C1(new_n1171), .C2(new_n854), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1167), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1162), .B1(new_n1173), .B2(new_n960), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT57), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1062), .A2(new_n1066), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1113), .B1(new_n1176), .B2(new_n1118), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1175), .B1(new_n1177), .B2(new_n1173), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1119), .A2(new_n1102), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1170), .B1(new_n1171), .B2(new_n854), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n893), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1165), .A2(new_n1181), .A3(new_n853), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1175), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n657), .B1(new_n1179), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1174), .B1(new_n1178), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(G375));
  NOR2_X1   g0986(.A1(new_n1104), .A2(new_n1110), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n1113), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n945), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1188), .A2(new_n1189), .A3(new_n1111), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n703), .B1(G68), .B2(new_n793), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1003), .B1(new_n737), .B2(new_n481), .C1(new_n733), .C2(new_n749), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n723), .A2(G294), .B1(G116), .B2(new_n742), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n728), .A2(G97), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n359), .B1(new_n747), .B2(G303), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1193), .A2(new_n978), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n359), .B1(new_n746), .B2(new_n1151), .C1(new_n222), .C2(new_n750), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n732), .B2(G137), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n347), .B2(new_n737), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1077), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n723), .A2(G132), .B1(new_n742), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n728), .A2(G159), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(new_n343), .C2(new_n740), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n1192), .A2(new_n1196), .B1(new_n1199), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1191), .B1(new_n717), .B2(new_n1204), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT121), .Z(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n715), .B2(new_n907), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n1187), .B2(new_n960), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1190), .A2(new_n1209), .ZN(G381));
  NAND4_X1  g1010(.A1(new_n962), .A2(new_n988), .A3(new_n1050), .A4(new_n1052), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1067), .A2(new_n1095), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1213), .A2(new_n1120), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1024), .A2(new_n773), .A3(new_n1026), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n1215), .A2(G384), .A3(G381), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1212), .A2(new_n1185), .A3(new_n1214), .A4(new_n1216), .ZN(G407));
  NAND2_X1  g1017(.A1(new_n638), .A2(G213), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1185), .A2(new_n1214), .A3(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(G407), .A2(G213), .A3(new_n1220), .ZN(G409));
  INV_X1    g1021(.A(KEYINPUT126), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1219), .A2(G2897), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1187), .A2(KEYINPUT60), .A3(new_n1113), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1225), .A2(KEYINPUT123), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(KEYINPUT123), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1102), .A2(new_n1104), .A3(new_n1110), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n656), .B(new_n1111), .C1(new_n1229), .C2(KEYINPUT60), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1209), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1231), .A2(new_n808), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G384), .B(new_n1209), .C1(new_n1228), .C2(new_n1230), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1224), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1231), .A2(new_n808), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1236), .A2(new_n1233), .A3(new_n1223), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1119), .A2(new_n1102), .B1(new_n1167), .B2(new_n1172), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n1189), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1240), .B(new_n1162), .C1(new_n960), .C2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1214), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT122), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n1185), .B2(G378), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1062), .A2(new_n1066), .A3(new_n1111), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1183), .B1(new_n1246), .B2(new_n1113), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1247), .B(new_n656), .C1(new_n1239), .C2(KEYINPUT57), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1167), .A2(new_n1172), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1249), .A2(new_n961), .B1(new_n1133), .B2(new_n1161), .ZN(new_n1250));
  AND4_X1   g1050(.A1(new_n1244), .A2(new_n1248), .A3(G378), .A4(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1243), .B1(new_n1245), .B2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1238), .B1(new_n1252), .B2(new_n1218), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1222), .B1(new_n1253), .B2(KEYINPUT61), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT61), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1248), .A2(new_n1250), .A3(G378), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(KEYINPUT122), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1185), .A2(new_n1244), .A3(G378), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1219), .B1(new_n1259), .B2(new_n1243), .ZN(new_n1260));
  OAI211_X1 g1060(.A(KEYINPUT126), .B(new_n1255), .C1(new_n1260), .C2(new_n1238), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1260), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1252), .A2(new_n1218), .A3(new_n1262), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT127), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1265), .A2(new_n1266), .A3(KEYINPUT62), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1254), .A2(new_n1261), .A3(new_n1264), .A4(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G387), .A2(G390), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G393), .A2(G396), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT125), .B1(new_n1270), .B2(new_n1215), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1215), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT125), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1269), .B(new_n1211), .C1(new_n1271), .C2(new_n1274), .ZN(new_n1275));
  AND2_X1   g1075(.A1(G387), .A2(G390), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(new_n1212), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1275), .B1(new_n1277), .B2(new_n1274), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1268), .A2(new_n1279), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1257), .A2(new_n1258), .B1(new_n1214), .B2(new_n1242), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1237), .B(new_n1235), .C1(new_n1281), .C2(new_n1219), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1282), .A2(new_n1278), .A3(new_n1255), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1260), .A2(KEYINPUT63), .A3(new_n1262), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT63), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT124), .B1(new_n1265), .B2(new_n1285), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1265), .A2(KEYINPUT124), .A3(new_n1285), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1283), .B(new_n1284), .C1(new_n1286), .C2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1280), .A2(new_n1288), .ZN(G405));
  INV_X1    g1089(.A(new_n1214), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1259), .B1(new_n1185), .B2(new_n1290), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(new_n1262), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1292), .B(new_n1279), .ZN(G402));
endmodule


