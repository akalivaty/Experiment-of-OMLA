//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1245, new_n1246, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1305,
    new_n1306;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AND2_X1   g0009(.A1(G107), .A2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n211), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n210), .B(new_n215), .C1(G116), .C2(G270), .ZN(new_n216));
  XOR2_X1   g0016(.A(KEYINPUT64), .B(G244), .Z(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G77), .ZN(new_n218));
  AND2_X1   g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n202), .C2(new_n222), .ZN(new_n223));
  AND2_X1   g0023(.A1(G50), .A2(G226), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n206), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(G50), .B1(G58), .B2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n209), .B(new_n226), .C1(new_n229), .C2(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT65), .B(KEYINPUT66), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XOR2_X1   g0039(.A(G238), .B(G244), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  AOI21_X1  g0049(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n250));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT67), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT67), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G1), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G41), .ZN(new_n256));
  INV_X1    g0056(.A(G45), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n250), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(G274), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n259), .A2(G232), .B1(new_n251), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G179), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G223), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G1698), .ZN(new_n266));
  AND2_X1   g0066(.A1(G226), .A2(G1698), .ZN(new_n267));
  AND2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  OAI22_X1  g0069(.A1(new_n266), .A2(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(new_n213), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AND3_X1   g0073(.A1(new_n270), .A2(KEYINPUT74), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(KEYINPUT74), .B1(new_n270), .B2(new_n273), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n250), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT75), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT74), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n271), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G223), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G226), .A2(G1698), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n281), .A2(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n279), .B1(new_n286), .B2(new_n272), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n270), .A2(KEYINPUT74), .A3(new_n273), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(KEYINPUT75), .A3(new_n250), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n264), .B1(new_n278), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(G169), .B1(new_n276), .B2(new_n262), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT76), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(G58), .B(G68), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G20), .A2(G33), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n294), .A2(G20), .B1(G159), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n281), .A2(new_n228), .A3(new_n282), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT7), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n281), .A2(KEYINPUT7), .A3(new_n228), .A4(new_n282), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(KEYINPUT73), .B1(new_n301), .B2(G68), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT73), .ZN(new_n303));
  AOI211_X1 g0103(.A(new_n303), .B(new_n211), .C1(new_n299), .C2(new_n300), .ZN(new_n304));
  OAI211_X1 g0104(.A(KEYINPUT16), .B(new_n296), .C1(new_n302), .C2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n227), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n301), .A2(G68), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n296), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT16), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n305), .A2(new_n307), .A3(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT8), .B(G58), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT69), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n313), .B(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n307), .B1(new_n255), .B2(G20), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(new_n315), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n312), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n264), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT75), .B1(new_n289), .B2(new_n250), .ZN(new_n322));
  INV_X1    g0122(.A(new_n250), .ZN(new_n323));
  AOI211_X1 g0123(.A(new_n277), .B(new_n323), .C1(new_n287), .C2(new_n288), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n321), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT76), .ZN(new_n326));
  INV_X1    g0126(.A(new_n292), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n293), .A2(new_n320), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT18), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n293), .A2(new_n320), .A3(new_n328), .A4(KEYINPUT18), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(KEYINPUT77), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT77), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n329), .A2(new_n334), .A3(new_n330), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT17), .ZN(new_n336));
  AOI21_X1  g0136(.A(G200), .B1(new_n276), .B2(new_n262), .ZN(new_n337));
  AOI21_X1  g0137(.A(G190), .B1(new_n278), .B2(new_n290), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(new_n262), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT78), .B1(new_n339), .B2(new_n320), .ZN(new_n340));
  INV_X1    g0140(.A(G190), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(new_n262), .C1(new_n322), .C2(new_n324), .ZN(new_n342));
  INV_X1    g0142(.A(new_n337), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT78), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n344), .A2(new_n345), .A3(new_n312), .A4(new_n319), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n336), .B1(new_n340), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n344), .A2(new_n312), .A3(new_n319), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n348), .A2(KEYINPUT17), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n333), .B(new_n335), .C1(new_n347), .C2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT13), .ZN(new_n351));
  OAI211_X1 g0151(.A(G226), .B(new_n283), .C1(new_n268), .C2(new_n269), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT70), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n281), .A2(new_n282), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT70), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n354), .A2(new_n355), .A3(G226), .A4(new_n283), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G33), .A2(G97), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n354), .A2(G232), .A3(G1698), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n353), .A2(new_n356), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n250), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n261), .A2(new_n251), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n259), .A2(G238), .ZN(new_n362));
  AND4_X1   g0162(.A1(new_n351), .A2(new_n360), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n359), .A2(new_n250), .B1(G238), .B2(new_n259), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n351), .B1(new_n364), .B2(new_n361), .ZN(new_n365));
  OAI21_X1  g0165(.A(G169), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT14), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n363), .A2(new_n365), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G179), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT14), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n370), .B(G169), .C1(new_n363), .C2(new_n365), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n367), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n271), .A2(G20), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(G77), .B1(G20), .B2(new_n211), .ZN(new_n374));
  INV_X1    g0174(.A(G50), .ZN(new_n375));
  INV_X1    g0175(.A(new_n295), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT71), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n377), .A2(new_n378), .A3(new_n307), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n378), .B1(new_n377), .B2(new_n307), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT11), .ZN(new_n381));
  OR3_X1    g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT67), .B(G1), .ZN(new_n383));
  INV_X1    g0183(.A(G13), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n383), .A2(new_n384), .A3(new_n228), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(KEYINPUT12), .A3(new_n211), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT12), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n316), .B2(G68), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n318), .A2(G68), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n390), .A2(KEYINPUT72), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(KEYINPUT72), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n381), .B1(new_n379), .B2(new_n380), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n382), .A2(new_n391), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n372), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n394), .B1(new_n368), .B2(G190), .ZN(new_n396));
  INV_X1    g0196(.A(G200), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n396), .B1(new_n397), .B2(new_n368), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n350), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n318), .A2(G50), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n385), .A2(new_n375), .ZN(new_n402));
  INV_X1    g0202(.A(G150), .ZN(new_n403));
  NOR3_X1   g0203(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n403), .A2(new_n376), .B1(new_n404), .B2(new_n228), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n405), .B1(new_n315), .B2(new_n373), .ZN(new_n406));
  INV_X1    g0206(.A(new_n307), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n401), .B(new_n402), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT9), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n313), .B(KEYINPUT69), .ZN(new_n410));
  INV_X1    g0210(.A(new_n373), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n307), .B1(new_n412), .B2(new_n405), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT9), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n413), .A2(new_n414), .A3(new_n401), .A4(new_n402), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n409), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n259), .A2(G226), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n361), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT68), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n283), .A2(G222), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n354), .B(new_n420), .C1(new_n265), .C2(new_n283), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n421), .B(new_n250), .C1(G77), .C2(new_n354), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT68), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n417), .A2(new_n423), .A3(new_n361), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n419), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G200), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n419), .A2(new_n422), .A3(new_n424), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G190), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n416), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT10), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT10), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n416), .A2(new_n428), .A3(new_n431), .A4(new_n426), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n427), .A2(new_n263), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n434), .B(new_n408), .C1(G169), .C2(new_n427), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n268), .A2(new_n269), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(G238), .B2(G1698), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n221), .B2(G1698), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n438), .B(new_n250), .C1(G107), .C2(new_n354), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n259), .A2(new_n217), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(new_n361), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G200), .ZN(new_n442));
  INV_X1    g0242(.A(new_n313), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n443), .A2(new_n295), .B1(G20), .B2(G77), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT15), .B(G87), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n411), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G77), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n446), .A2(new_n307), .B1(new_n447), .B2(new_n385), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n318), .A2(G77), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n442), .B(new_n451), .C1(new_n341), .C2(new_n441), .ZN(new_n452));
  INV_X1    g0252(.A(G169), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n441), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n454), .B(new_n450), .C1(G179), .C2(new_n441), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n433), .A2(new_n435), .A3(new_n452), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(KEYINPUT79), .B1(new_n400), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT79), .ZN(new_n459));
  NOR4_X1   g0259(.A1(new_n350), .A2(new_n456), .A3(new_n399), .A4(new_n459), .ZN(new_n460));
  OR2_X1    g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n354), .A2(new_n228), .A3(G68), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n357), .A2(G20), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(KEYINPUT19), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(KEYINPUT19), .B1(new_n204), .B2(G87), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n465), .B1(new_n228), .B2(new_n357), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n307), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n255), .A2(G33), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n316), .A2(new_n407), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G87), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n385), .A2(new_n445), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n467), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n212), .A2(new_n283), .ZN(new_n474));
  OAI221_X1 g0274(.A(new_n474), .B1(G244), .B2(new_n283), .C1(new_n268), .C2(new_n269), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G116), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n250), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n214), .B1(new_n383), .B2(new_n257), .ZN(new_n479));
  INV_X1    g0279(.A(G274), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n255), .A2(G45), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(new_n481), .A3(new_n323), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G200), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n473), .B(new_n484), .C1(new_n341), .C2(new_n483), .ZN(new_n485));
  INV_X1    g0285(.A(new_n483), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n263), .ZN(new_n487));
  INV_X1    g0287(.A(new_n445), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n469), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n467), .A2(new_n489), .A3(new_n471), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n487), .B(new_n490), .C1(G169), .C2(new_n486), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n485), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT24), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n228), .B(G87), .C1(new_n268), .C2(new_n269), .ZN(new_n494));
  NAND2_X1  g0294(.A1(KEYINPUT87), .A2(KEYINPUT22), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT88), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT88), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(KEYINPUT87), .A3(KEYINPUT22), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g0299(.A(new_n494), .B(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT23), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n501), .B1(new_n228), .B2(G107), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n502), .A2(new_n503), .B1(new_n373), .B2(G116), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n493), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n499), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n507), .A2(new_n494), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n507), .A2(new_n494), .ZN(new_n509));
  OAI211_X1 g0309(.A(KEYINPUT24), .B(new_n504), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n506), .A2(new_n307), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n469), .A2(G107), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n316), .A2(G107), .ZN(new_n513));
  XNOR2_X1  g0313(.A(new_n513), .B(KEYINPUT25), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n511), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n222), .A2(G1698), .ZN(new_n516));
  OAI221_X1 g0316(.A(new_n516), .B1(G250), .B2(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n517));
  INV_X1    g0317(.A(G294), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n517), .B1(new_n271), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n250), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n256), .A2(KEYINPUT5), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n383), .A2(new_n257), .A3(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT5), .ZN(new_n523));
  OAI21_X1  g0323(.A(KEYINPUT81), .B1(new_n523), .B2(G41), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT81), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(new_n256), .A3(KEYINPUT5), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n522), .A2(G274), .A3(new_n323), .A4(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n257), .B1(new_n252), .B2(new_n254), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n523), .A2(G41), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(G264), .A3(new_n323), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n520), .A2(new_n528), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(new_n341), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n515), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(G200), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n492), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT21), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n316), .A2(new_n468), .A3(G116), .A4(new_n407), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G283), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT80), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(KEYINPUT80), .A2(G33), .A3(G283), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(G20), .B1(new_n271), .B2(G97), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(G116), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n306), .A2(new_n227), .B1(G20), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n548), .A3(KEYINPUT20), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT20), .B1(new_n546), .B2(new_n548), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n539), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n385), .A2(KEYINPUT86), .A3(new_n547), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT86), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n316), .B2(G116), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(G169), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n283), .A2(G257), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G264), .A2(G1698), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n558), .B(new_n559), .C1(new_n268), .C2(new_n269), .ZN(new_n560));
  XNOR2_X1  g0360(.A(KEYINPUT85), .B(G303), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n560), .B(new_n250), .C1(new_n354), .C2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n529), .A2(new_n527), .A3(G274), .A4(new_n530), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n562), .B1(new_n563), .B2(new_n250), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n531), .A2(G270), .A3(new_n323), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT84), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT84), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n531), .A2(new_n568), .A3(G270), .A4(new_n323), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n565), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n538), .B1(new_n557), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n553), .A2(new_n555), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n572), .B(new_n539), .C1(new_n551), .C2(new_n550), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n570), .A2(G179), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n565), .A2(new_n567), .A3(new_n569), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n573), .A2(new_n575), .A3(KEYINPUT21), .A4(G169), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n571), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n533), .A2(new_n453), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n520), .A2(new_n532), .A3(new_n528), .A4(new_n263), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n580), .A2(new_n515), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n567), .A2(new_n569), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(G190), .A3(new_n565), .ZN(new_n583));
  INV_X1    g0383(.A(new_n573), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n575), .A2(G200), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n577), .A2(new_n581), .A3(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(G244), .B(new_n283), .C1(new_n268), .C2(new_n269), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT4), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n354), .A2(KEYINPUT4), .A3(G244), .A4(new_n283), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n354), .A2(G250), .A3(G1698), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n593), .A2(new_n544), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n323), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n253), .A2(G1), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n251), .A2(KEYINPUT67), .ZN(new_n597));
  OAI211_X1 g0397(.A(G45), .B(new_n530), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n524), .A2(new_n526), .ZN(new_n599));
  OAI211_X1 g0399(.A(G257), .B(new_n323), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n528), .A2(new_n600), .ZN(new_n601));
  NOR3_X1   g0401(.A1(new_n595), .A2(KEYINPUT83), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT83), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n528), .A2(new_n600), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n590), .A2(new_n591), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n593), .A2(new_n544), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n250), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n603), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(G190), .B1(new_n602), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n203), .A2(KEYINPUT6), .A3(G97), .ZN(new_n610));
  XOR2_X1   g0410(.A(G97), .B(G107), .Z(new_n611));
  OAI21_X1  g0411(.A(new_n610), .B1(new_n611), .B2(KEYINPUT6), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n612), .A2(G20), .B1(G77), .B2(new_n295), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n301), .A2(G107), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n407), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n469), .A2(G97), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n316), .A2(G97), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT82), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n528), .A2(new_n600), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n619), .B1(new_n528), .B2(new_n600), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n607), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(G200), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n609), .A2(new_n618), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n618), .ZN(new_n625));
  OAI21_X1  g0425(.A(KEYINPUT83), .B1(new_n595), .B2(new_n601), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n604), .A2(new_n603), .A3(new_n607), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n627), .A3(new_n453), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n263), .B(new_n607), .C1(new_n620), .C2(new_n621), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n625), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  AND4_X1   g0431(.A1(new_n461), .A2(new_n537), .A3(new_n587), .A4(new_n631), .ZN(G372));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n487), .A2(new_n490), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT89), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n482), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT89), .A4(new_n323), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n478), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n453), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n634), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n639), .A2(G200), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n642), .B(new_n473), .C1(new_n341), .C2(new_n483), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT92), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n628), .A2(new_n629), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT91), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n628), .A2(KEYINPUT91), .A3(new_n629), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n646), .B1(new_n651), .B2(new_n625), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n628), .A2(KEYINPUT91), .A3(new_n629), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT91), .B1(new_n628), .B2(new_n629), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n646), .B(new_n625), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n633), .B(new_n645), .C1(new_n652), .C2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n577), .A2(KEYINPUT90), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT90), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n571), .A2(new_n574), .A3(new_n576), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n580), .A2(new_n515), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n535), .A2(new_n536), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n663), .A2(new_n664), .A3(new_n631), .A4(new_n645), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n492), .A2(new_n630), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n641), .B1(new_n666), .B2(new_n633), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n657), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n461), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n331), .A2(new_n332), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n340), .A2(new_n346), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n349), .B1(new_n672), .B2(KEYINPUT17), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n395), .B2(new_n455), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n671), .B1(new_n674), .B2(new_n398), .ZN(new_n675));
  INV_X1    g0475(.A(new_n433), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n435), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n670), .A2(new_n678), .ZN(G369));
  INV_X1    g0479(.A(new_n577), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n384), .A2(G20), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  OR3_X1    g0482(.A1(new_n383), .A2(new_n682), .A3(KEYINPUT27), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT27), .B1(new_n383), .B2(new_n682), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(new_n684), .A3(G213), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n584), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n680), .A2(new_n689), .ZN(new_n690));
  AOI211_X1 g0490(.A(new_n586), .B(new_n690), .C1(new_n661), .C2(new_n689), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G330), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n662), .A2(new_n687), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n515), .A2(new_n687), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n664), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n693), .B1(new_n695), .B2(new_n662), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n680), .A2(new_n687), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n696), .A2(new_n697), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n693), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n702), .ZN(G399));
  INV_X1    g0503(.A(new_n207), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G1), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n230), .B2(new_n706), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n680), .A2(new_n662), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n711), .A2(new_n631), .A3(new_n664), .A4(new_n645), .ZN(new_n712));
  INV_X1    g0512(.A(new_n641), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n713), .B1(new_n666), .B2(new_n633), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n625), .B1(new_n653), .B2(new_n654), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT92), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n644), .B1(new_n716), .B2(new_n655), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n712), .B(new_n714), .C1(new_n717), .C2(new_n633), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(KEYINPUT29), .A3(new_n688), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n667), .B1(new_n717), .B2(new_n633), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n687), .B1(new_n720), .B2(new_n665), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n719), .B1(new_n721), .B2(KEYINPUT29), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n587), .A2(new_n631), .A3(new_n537), .A4(new_n688), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n626), .A2(new_n627), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n565), .A2(new_n567), .A3(G179), .A4(new_n569), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n520), .A2(new_n478), .A3(new_n532), .A4(new_n482), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n725), .A2(new_n728), .A3(KEYINPUT30), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT30), .B1(new_n725), .B2(new_n728), .ZN(new_n730));
  AOI21_X1  g0530(.A(G179), .B1(new_n638), .B2(new_n478), .ZN(new_n731));
  AND4_X1   g0531(.A1(new_n533), .A2(new_n622), .A3(new_n575), .A4(new_n731), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n724), .B1(new_n733), .B2(new_n688), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n602), .A2(new_n608), .ZN(new_n736));
  INV_X1    g0536(.A(new_n727), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n737), .A2(new_n582), .A3(G179), .A4(new_n565), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n735), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n725), .A2(new_n728), .A3(KEYINPUT30), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n622), .A2(new_n731), .A3(new_n533), .A4(new_n575), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n723), .A2(new_n734), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G330), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n722), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n710), .B1(new_n746), .B2(G1), .ZN(G364));
  NAND2_X1  g0547(.A1(new_n681), .A2(G45), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n706), .A2(G1), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n692), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n691), .A2(G330), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n245), .A2(G45), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n704), .A2(new_n354), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n752), .B(new_n753), .C1(G45), .C2(new_n230), .ZN(new_n754));
  INV_X1    g0554(.A(G355), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n354), .A2(new_n207), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n754), .B1(G116), .B2(new_n207), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n228), .B1(KEYINPUT93), .B2(new_n453), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(KEYINPUT93), .B2(new_n453), .ZN(new_n759));
  INV_X1    g0559(.A(new_n227), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G13), .A2(G33), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n757), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n749), .ZN(new_n768));
  INV_X1    g0568(.A(new_n765), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n767), .B(new_n768), .C1(new_n691), .C2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n228), .A2(new_n263), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n772), .A2(new_n341), .A3(G200), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G322), .ZN(new_n775));
  INV_X1    g0575(.A(G283), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n228), .A2(G179), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n397), .A2(G190), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n774), .A2(new_n775), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G179), .A2(G200), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT94), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n782), .A2(G190), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n228), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n782), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G329), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n771), .A2(new_n778), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G317), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(KEYINPUT33), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n790), .A2(KEYINPUT33), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n789), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n784), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G294), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n341), .A2(new_n397), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n771), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n354), .B1(new_n798), .B2(G326), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n787), .A2(new_n793), .A3(new_n795), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n796), .A2(new_n777), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n780), .B(new_n800), .C1(G303), .C2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G311), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n772), .A2(G190), .A3(G200), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n803), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G159), .ZN(new_n808));
  OR3_X1    g0608(.A1(new_n785), .A2(KEYINPUT32), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n354), .B1(new_n788), .B2(new_n211), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(new_n794), .B2(G97), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n773), .A2(G58), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n802), .A2(G87), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n798), .A2(G50), .ZN(new_n814));
  INV_X1    g0614(.A(new_n779), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G107), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n812), .A2(new_n813), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G77), .B2(new_n805), .ZN(new_n818));
  OAI21_X1  g0618(.A(KEYINPUT32), .B1(new_n785), .B2(new_n808), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n809), .A2(new_n811), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n761), .B1(new_n807), .B2(new_n820), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n750), .A2(new_n751), .B1(new_n770), .B2(new_n821), .ZN(G396));
  OAI21_X1  g0622(.A(new_n452), .B1(new_n451), .B2(new_n688), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n455), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n455), .A2(new_n687), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n721), .B(new_n826), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(new_n745), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n749), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n784), .A2(new_n202), .B1(new_n518), .B2(new_n774), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT95), .Z(new_n831));
  AOI211_X1 g0631(.A(new_n354), .B(new_n831), .C1(G311), .C2(new_n786), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n798), .A2(G303), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n779), .A2(new_n213), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n806), .A2(new_n547), .B1(new_n801), .B2(new_n203), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n834), .B(new_n835), .C1(G283), .C2(new_n789), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n832), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT96), .Z(new_n838));
  NOR2_X1   g0638(.A1(new_n779), .A2(new_n211), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n840), .B(new_n354), .C1(new_n375), .C2(new_n801), .ZN(new_n841));
  XOR2_X1   g0641(.A(KEYINPUT97), .B(G143), .Z(new_n842));
  AOI22_X1  g0642(.A1(new_n842), .A2(new_n773), .B1(new_n805), .B2(G159), .ZN(new_n843));
  INV_X1    g0643(.A(G137), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n843), .B1(new_n844), .B2(new_n797), .C1(new_n403), .C2(new_n788), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT34), .Z(new_n846));
  AOI211_X1 g0646(.A(new_n841), .B(new_n846), .C1(G132), .C2(new_n786), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n220), .B2(new_n784), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n761), .B1(new_n838), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n762), .A2(new_n763), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n826), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n768), .B1(G77), .B2(new_n851), .C1(new_n852), .C2(new_n764), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n829), .A2(new_n854), .ZN(G384));
  INV_X1    g0655(.A(KEYINPUT102), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n742), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT31), .B1(new_n742), .B2(new_n687), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n856), .B1(new_n859), .B2(new_n723), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n723), .A2(new_n734), .A3(new_n856), .A4(new_n743), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT99), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n394), .A2(new_n687), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n372), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n864), .B1(new_n372), .B2(new_n866), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n395), .A2(new_n398), .A3(new_n865), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n826), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n302), .A2(new_n304), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT16), .B1(new_n872), .B2(new_n296), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n305), .A2(new_n307), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n319), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n685), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n333), .A2(new_n335), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n878), .B1(new_n879), .B2(new_n673), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n875), .A2(new_n328), .A3(new_n293), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n672), .A2(new_n877), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT37), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n320), .A2(new_n876), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n329), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT37), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(new_n886), .A3(new_n672), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n880), .A2(KEYINPUT38), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n880), .B2(new_n888), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n863), .B(new_n871), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT40), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n340), .A2(new_n346), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n329), .A2(new_n886), .A3(new_n884), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT100), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n329), .A2(new_n348), .A3(new_n884), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT37), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT100), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n885), .A2(new_n672), .A3(new_n899), .A4(new_n886), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n896), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n320), .B(new_n876), .C1(new_n673), .C2(new_n671), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT38), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n880), .A2(new_n888), .A3(KEYINPUT38), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n893), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n744), .A2(KEYINPUT102), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n871), .A2(new_n908), .A3(new_n861), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n891), .A2(new_n892), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n911), .A2(new_n461), .A3(new_n863), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n889), .A2(new_n890), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n892), .B1(new_n913), .B2(new_n909), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n905), .A2(new_n906), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n915), .A2(new_n910), .A3(KEYINPUT40), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n914), .A2(G330), .A3(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n863), .B(G330), .C1(new_n458), .C2(new_n460), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n912), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n395), .A2(new_n687), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT38), .B1(new_n901), .B2(new_n902), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n921), .B1(new_n889), .B2(new_n922), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n889), .A2(new_n890), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n920), .B(new_n923), .C1(new_n924), .C2(new_n921), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n671), .A2(new_n685), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n869), .A2(new_n870), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n669), .A2(new_n688), .A3(new_n852), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n927), .B1(new_n928), .B2(new_n825), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n924), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n925), .A2(new_n926), .A3(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n919), .B(new_n931), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n718), .A2(KEYINPUT29), .A3(new_n688), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT29), .B1(new_n669), .B2(new_n688), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n677), .B1(new_n935), .B2(new_n461), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n932), .B(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n255), .B2(new_n681), .ZN(new_n938));
  OAI211_X1 g0738(.A(G116), .B(new_n229), .C1(new_n612), .C2(KEYINPUT35), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT98), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n612), .A2(KEYINPUT35), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT36), .ZN(new_n943));
  OAI21_X1  g0743(.A(G77), .B1(new_n220), .B2(new_n211), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n944), .A2(new_n230), .B1(G50), .B2(new_n211), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(new_n384), .A3(new_n383), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n938), .A2(new_n943), .A3(new_n946), .ZN(G367));
  NAND2_X1  g0747(.A1(new_n701), .A2(new_n631), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT42), .Z(new_n949));
  OAI21_X1  g0749(.A(new_n631), .B1(new_n618), .B2(new_n688), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n651), .A2(new_n625), .A3(new_n687), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n630), .B1(new_n953), .B2(new_n662), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n688), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n949), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n472), .A2(new_n687), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n713), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n644), .B2(new_n957), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT103), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n956), .A2(new_n963), .B1(KEYINPUT43), .B2(new_n961), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n963), .B2(new_n956), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n700), .A2(new_n953), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n965), .A2(new_n966), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT105), .Z(new_n969));
  XNOR2_X1  g0769(.A(new_n705), .B(KEYINPUT41), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n701), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(KEYINPUT106), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n692), .A2(new_n698), .ZN(new_n974));
  AND3_X1   g0774(.A1(new_n700), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n973), .B1(new_n700), .B2(new_n974), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n746), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT107), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n978), .B(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n702), .A2(new_n952), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT45), .Z(new_n982));
  NOR2_X1   g0782(.A1(new_n702), .A2(new_n952), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT44), .ZN(new_n984));
  AND3_X1   g0784(.A1(new_n982), .A2(new_n700), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n700), .B1(new_n982), .B2(new_n984), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n980), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n971), .B1(new_n988), .B2(new_n746), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n748), .A2(G1), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n967), .B(new_n969), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n766), .B1(new_n207), .B2(new_n445), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n237), .B2(new_n753), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n794), .A2(G68), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n773), .A2(G150), .B1(G159), .B2(new_n789), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(new_n375), .C2(new_n806), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n785), .A2(new_n844), .B1(new_n447), .B2(new_n779), .ZN(new_n997));
  INV_X1    g0797(.A(new_n842), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n354), .B1(new_n998), .B2(new_n797), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n996), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n220), .B2(new_n801), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n802), .A2(G116), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT46), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n1002), .A2(new_n1003), .B1(new_n805), .B2(G283), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n202), .B2(new_n779), .C1(new_n518), .C2(new_n788), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G317), .B2(new_n786), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n773), .A2(new_n561), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n354), .B1(new_n794), .B2(G107), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT108), .Z(new_n1010));
  NAND4_X1  g0810(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n797), .A2(new_n804), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1001), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT47), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n993), .B1(new_n1014), .B2(new_n762), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1015), .B(new_n768), .C1(new_n961), .C2(new_n769), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n991), .A2(new_n1016), .ZN(G387));
  OAI21_X1  g0817(.A(new_n768), .B1(new_n696), .B2(new_n769), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n561), .A2(new_n805), .B1(new_n773), .B2(G317), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n804), .B2(new_n788), .C1(new_n775), .C2(new_n797), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT48), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n776), .B2(new_n784), .C1(new_n518), .C2(new_n801), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT49), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n786), .A2(G326), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n354), .B1(new_n815), .B2(G116), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n794), .A2(new_n488), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n211), .B2(new_n806), .C1(new_n410), .C2(new_n788), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G150), .B2(new_n786), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n773), .A2(G50), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n779), .A2(new_n202), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n801), .A2(new_n447), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(G159), .C2(new_n798), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1029), .A2(new_n354), .A3(new_n1030), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n761), .B1(new_n1026), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n241), .A2(G45), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT109), .Z(new_n1037));
  XOR2_X1   g0837(.A(new_n707), .B(KEYINPUT110), .Z(new_n1038));
  NOR2_X1   g0838(.A1(new_n313), .A2(G50), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT50), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(G68), .A2(G77), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1038), .A2(new_n1040), .A3(new_n257), .A4(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1037), .A2(new_n753), .A3(new_n1042), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(G107), .B2(new_n207), .C1(new_n707), .C2(new_n756), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1018), .B(new_n1035), .C1(new_n766), .C2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n977), .B2(new_n990), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n978), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n705), .B1(new_n977), .B2(new_n746), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1046), .B1(new_n1047), .B2(new_n1048), .ZN(G393));
  OAI211_X1 g0849(.A(new_n988), .B(new_n705), .C1(new_n987), .C2(new_n1047), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n987), .A2(KEYINPUT111), .B1(G1), .B2(new_n748), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(KEYINPUT111), .B2(new_n987), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n952), .A2(new_n769), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1053), .A2(KEYINPUT112), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n354), .B1(new_n786), .B2(G322), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n773), .A2(G311), .B1(new_n798), .B2(G317), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1055), .B1(KEYINPUT52), .B2(new_n1056), .C1(new_n776), .C2(new_n801), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n1056), .A2(KEYINPUT52), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n806), .A2(new_n518), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n789), .A2(new_n561), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n816), .B(new_n1060), .C1(new_n784), .C2(new_n547), .ZN(new_n1061));
  NOR4_X1   g0861(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .A4(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n794), .A2(G77), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n773), .A2(G159), .B1(new_n798), .B2(G150), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(KEYINPUT51), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n785), .A2(new_n998), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n801), .A2(new_n211), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n805), .A2(new_n443), .B1(G50), .B2(new_n789), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n834), .A2(new_n436), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(new_n1064), .C2(KEYINPUT51), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .A4(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n762), .B1(new_n1062), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1053), .A2(KEYINPUT112), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n753), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n766), .B1(new_n202), .B2(new_n207), .C1(new_n248), .C2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n768), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT113), .Z(new_n1078));
  NAND4_X1  g0878(.A1(new_n1054), .A2(new_n1073), .A3(new_n1074), .A4(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1050), .A2(new_n1052), .A3(new_n1079), .ZN(G390));
  NOR3_X1   g0880(.A1(new_n889), .A2(new_n890), .A3(new_n921), .ZN(new_n1081));
  AOI21_X1  g0881(.A(KEYINPUT39), .B1(new_n905), .B2(new_n906), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n929), .A2(new_n920), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n718), .A2(new_n688), .A3(new_n824), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n825), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n927), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n920), .B1(new_n905), .B2(new_n906), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n744), .A2(G330), .A3(new_n852), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1090), .A2(new_n927), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n1083), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n871), .A2(new_n908), .A3(G330), .A4(new_n861), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n923), .B1(new_n924), .B2(new_n921), .ZN(new_n1096));
  INV_X1    g0896(.A(G125), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n785), .A2(new_n1097), .B1(new_n808), .B2(new_n784), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n802), .A2(G150), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT53), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n773), .A2(G132), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n844), .B2(new_n788), .ZN(new_n1102));
  XOR2_X1   g0902(.A(KEYINPUT54), .B(G143), .Z(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n354), .B1(new_n806), .B2(new_n1104), .ZN(new_n1105));
  NOR4_X1   g0905(.A1(new_n1098), .A2(new_n1100), .A3(new_n1102), .A4(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(G128), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1106), .B1(new_n375), .B2(new_n779), .C1(new_n1107), .C2(new_n797), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1063), .B1(new_n202), .B2(new_n806), .C1(new_n203), .C2(new_n788), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G294), .B2(new_n786), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n773), .A2(G116), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1110), .A2(new_n813), .A3(new_n840), .A4(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n436), .B1(new_n797), .B2(new_n776), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1108), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1096), .A2(new_n763), .B1(new_n762), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n749), .B1(new_n850), .B2(new_n410), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT117), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1095), .A2(new_n990), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT114), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1090), .A2(new_n927), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n908), .A2(G330), .A3(new_n852), .A4(new_n861), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1120), .B1(new_n1121), .B2(new_n927), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1084), .A2(new_n825), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1090), .A2(new_n927), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1093), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n928), .A2(new_n825), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1122), .A2(new_n1123), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n458), .A2(new_n460), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n918), .B(new_n678), .C1(new_n722), .C2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1119), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1121), .A2(new_n927), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1131), .A2(new_n825), .A3(new_n1084), .A4(new_n1091), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1134), .A2(new_n936), .A3(KEYINPUT114), .A4(new_n918), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n1130), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1083), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1126), .A2(new_n1086), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n920), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1140), .A2(new_n1096), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1137), .B1(new_n1141), .B2(new_n1093), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1136), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT115), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1136), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1130), .A2(new_n1135), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT115), .B1(new_n1095), .B2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n705), .B(new_n1143), .C1(new_n1145), .C2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT116), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1144), .B1(new_n1136), .B2(new_n1142), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1095), .A2(KEYINPUT115), .A3(new_n1146), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n706), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(KEYINPUT116), .B1(new_n1153), .B2(new_n1143), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1118), .B1(new_n1150), .B2(new_n1154), .ZN(G378));
  INV_X1    g0955(.A(KEYINPUT120), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n433), .A2(new_n435), .ZN(new_n1157));
  XOR2_X1   g0957(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1158));
  XOR2_X1   g0958(.A(new_n1157), .B(new_n1158), .Z(new_n1159));
  NAND2_X1  g0959(.A1(new_n408), .A2(new_n876), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1159), .B(new_n1160), .Z(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n911), .B2(G330), .ZN(new_n1162));
  AND4_X1   g0962(.A1(G330), .A2(new_n914), .A3(new_n916), .A4(new_n1161), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n931), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1161), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n917), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n925), .A2(new_n926), .A3(new_n930), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n914), .A2(new_n1161), .A3(new_n916), .A4(G330), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1156), .B1(new_n1164), .B2(new_n1169), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1169), .A2(new_n1156), .ZN(new_n1171));
  OAI21_X1  g0971(.A(KEYINPUT121), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1167), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1174));
  OAI21_X1  g0974(.A(KEYINPUT120), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT121), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1169), .A2(new_n1156), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1172), .A2(new_n1178), .A3(new_n990), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n794), .A2(G68), .B1(new_n488), .B2(new_n805), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1180), .B1(new_n203), .B2(new_n774), .C1(new_n776), .C2(new_n785), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1032), .B(new_n1181), .C1(G97), .C2(new_n789), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n779), .A2(new_n220), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT118), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1185), .A2(G41), .A3(new_n354), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1182), .B(new_n1186), .C1(new_n547), .C2(new_n797), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT58), .Z(new_n1188));
  OAI21_X1  g0988(.A(new_n375), .B1(new_n268), .B2(G41), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n774), .A2(new_n1107), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n805), .A2(G137), .B1(G132), .B2(new_n789), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT119), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n1097), .B2(new_n797), .C1(new_n801), .C2(new_n1104), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1190), .B(new_n1193), .C1(G150), .C2(new_n794), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT59), .ZN(new_n1195));
  AOI21_X1  g0995(.A(G33), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G41), .B1(new_n786), .B2(G124), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(new_n808), .C2(new_n779), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1189), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n762), .B1(new_n1188), .B2(new_n1200), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1201), .A2(new_n768), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(G50), .B2(new_n851), .C1(new_n1165), .C2(new_n764), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1179), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT57), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1172), .A2(new_n1178), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1129), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1205), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n936), .B(new_n918), .C1(new_n1145), .C2(new_n1147), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1205), .B1(new_n1164), .B2(new_n1169), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n706), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1204), .B1(new_n1208), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(G375));
  AOI21_X1  g1013(.A(new_n1146), .B1(new_n1129), .B2(new_n1127), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n970), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1027), .B1(new_n518), .B2(new_n797), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n354), .B(new_n1216), .C1(G303), .C2(new_n786), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n788), .A2(new_n547), .B1(new_n779), .B2(new_n447), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G97), .B2(new_n802), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n203), .B2(new_n806), .C1(new_n776), .C2(new_n774), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1104), .A2(new_n788), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1185), .A2(KEYINPUT122), .A3(new_n436), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G132), .B2(new_n798), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n773), .A2(G137), .ZN(new_n1225));
  OAI21_X1  g1025(.A(KEYINPUT122), .B1(new_n1185), .B2(new_n436), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n785), .A2(new_n1107), .B1(new_n375), .B2(new_n784), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n806), .A2(new_n403), .B1(new_n801), .B2(new_n808), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1221), .B1(new_n1222), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n762), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1232), .B(new_n768), .C1(new_n764), .C2(new_n1086), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n211), .B2(new_n850), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n1134), .B2(new_n990), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1215), .A2(new_n1235), .ZN(G381));
  NAND2_X1  g1036(.A1(new_n1148), .A2(new_n1118), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(G375), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(G384), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(G381), .A2(G396), .A3(G393), .ZN(new_n1240));
  INV_X1    g1040(.A(G390), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(new_n991), .A3(new_n1016), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .A4(new_n1243), .ZN(G407));
  INV_X1    g1044(.A(G213), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n1238), .B2(new_n686), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(G407), .ZN(G409));
  NAND2_X1  g1047(.A1(G387), .A2(G390), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1242), .ZN(new_n1249));
  XOR2_X1   g1049(.A(G393), .B(G396), .Z(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1250), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1248), .A2(new_n1242), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT60), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1129), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1255), .B1(new_n1256), .B2(new_n1134), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n705), .B(new_n1257), .C1(new_n1214), .C2(new_n1255), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1235), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1239), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(G384), .A3(new_n1235), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1245), .A2(G343), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(G2897), .ZN(new_n1264));
  XOR2_X1   g1064(.A(new_n1264), .B(KEYINPUT124), .Z(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1262), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1260), .A2(new_n1261), .A3(new_n1265), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1269), .A2(KEYINPUT125), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT125), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1208), .A2(new_n1211), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1204), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(G378), .A3(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1209), .A2(new_n970), .A3(new_n1172), .A4(new_n1178), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n990), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT123), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1278), .A2(new_n1279), .A3(new_n1203), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1279), .B1(new_n1278), .B2(new_n1203), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1237), .B1(new_n1277), .B2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1263), .B1(new_n1276), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1254), .B1(new_n1273), .B2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT61), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT63), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1289), .B1(new_n1286), .B2(new_n1262), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1262), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1285), .A2(KEYINPUT63), .A3(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1287), .A2(new_n1288), .A3(new_n1290), .A4(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1288), .B1(new_n1285), .B2(new_n1269), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(new_n1285), .B2(new_n1291), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1283), .B1(new_n1212), .B2(G378), .ZN(new_n1298));
  NOR4_X1   g1098(.A1(new_n1298), .A2(new_n1263), .A3(new_n1262), .A4(new_n1295), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1294), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1254), .B(KEYINPUT127), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1293), .B1(new_n1302), .B2(new_n1303), .ZN(G405));
  OAI21_X1  g1104(.A(new_n1276), .B1(new_n1212), .B2(new_n1237), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1305), .B(new_n1291), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1306), .B(new_n1254), .ZN(G402));
endmodule


