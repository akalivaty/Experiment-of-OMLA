//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(KEYINPUT64), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n208), .B1(new_n209), .B2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G13), .ZN(new_n211));
  NAND4_X1  g0011(.A1(new_n211), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n202), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n217), .A2(G20), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G87), .A2(G250), .ZN(new_n222));
  INV_X1    g0022(.A(G58), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(G107), .B2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT65), .B(G68), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G238), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n230));
  NAND4_X1  g0030(.A1(new_n226), .A2(new_n228), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(new_n209), .ZN(new_n232));
  OR2_X1    g0032(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT66), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n221), .B(new_n234), .C1(KEYINPUT1), .C2(new_n232), .ZN(G361));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT69), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n248), .B(new_n252), .ZN(G351));
  OR2_X1    g0053(.A1(KEYINPUT74), .A2(KEYINPUT10), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT74), .A2(KEYINPUT10), .ZN(new_n255));
  OAI21_X1  g0055(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n256));
  INV_X1    g0056(.A(G150), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G20), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G33), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT8), .B(G58), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n256), .B1(new_n257), .B2(new_n259), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n218), .ZN(new_n265));
  INV_X1    g0065(.A(G50), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n211), .A2(new_n260), .A3(G1), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n263), .A2(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G20), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n267), .A2(new_n265), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT71), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR3_X1   g0073(.A1(new_n267), .A2(new_n265), .A3(KEYINPUT71), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n268), .B1(new_n275), .B2(new_n266), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT9), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n276), .B1(KEYINPUT73), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(KEYINPUT73), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  INV_X1    g0081(.A(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(G222), .A3(new_n286), .ZN(new_n287));
  XOR2_X1   g0087(.A(new_n287), .B(KEYINPUT70), .Z(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G223), .ZN(new_n290));
  INV_X1    g0090(.A(G77), .ZN(new_n291));
  OAI22_X1  g0091(.A1(new_n289), .A2(new_n290), .B1(new_n291), .B2(new_n285), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G41), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n219), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n269), .B1(G41), .B2(G45), .ZN(new_n297));
  INV_X1    g0097(.A(G274), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n295), .A2(new_n297), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n299), .B1(new_n301), .B2(G226), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(G200), .B1(new_n296), .B2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(G190), .B(new_n302), .C1(new_n293), .C2(new_n295), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n254), .B(new_n255), .C1(new_n280), .C2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n306), .ZN(new_n308));
  INV_X1    g0108(.A(new_n279), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n278), .B(new_n309), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n308), .A2(new_n310), .A3(KEYINPUT74), .A4(KEYINPUT10), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(new_n296), .B2(new_n303), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n314), .B(new_n302), .C1(new_n293), .C2(new_n295), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(new_n276), .A3(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n307), .A2(new_n311), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n290), .A2(new_n286), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n285), .B(new_n318), .C1(G226), .C2(new_n286), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G33), .A2(G87), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n295), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n299), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n300), .B2(new_n224), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n321), .A2(new_n323), .A3(new_n314), .ZN(new_n324));
  INV_X1    g0124(.A(new_n321), .ZN(new_n325));
  INV_X1    g0125(.A(new_n323), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n324), .B1(G169), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n265), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n201), .B1(new_n227), .B2(G58), .ZN(new_n330));
  INV_X1    g0130(.A(G159), .ZN(new_n331));
  OAI22_X1  g0131(.A1(new_n330), .A2(new_n260), .B1(new_n331), .B2(new_n259), .ZN(new_n332));
  INV_X1    g0132(.A(G68), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n283), .A2(new_n260), .A3(new_n284), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT7), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n283), .A2(KEYINPUT7), .A3(new_n260), .A4(new_n284), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n333), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n329), .B1(new_n339), .B2(KEYINPUT16), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT79), .ZN(new_n341));
  AND2_X1   g0141(.A1(KEYINPUT3), .A2(G33), .ZN(new_n342));
  NOR2_X1   g0142(.A1(KEYINPUT3), .A2(G33), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n342), .A2(new_n343), .A3(G20), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n341), .B1(new_n344), .B2(KEYINPUT7), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n334), .A2(KEYINPUT79), .A3(new_n335), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT80), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n337), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n337), .A2(new_n347), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n345), .B(new_n346), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n332), .B1(new_n350), .B2(new_n227), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n340), .B1(new_n351), .B2(KEYINPUT16), .ZN(new_n352));
  INV_X1    g0152(.A(new_n262), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n275), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n267), .B2(new_n353), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n328), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n356), .B(KEYINPUT18), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n325), .A2(G190), .A3(new_n326), .ZN(new_n358));
  OAI21_X1  g0158(.A(G200), .B1(new_n321), .B2(new_n323), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n352), .A2(new_n355), .A3(new_n360), .ZN(new_n361));
  XNOR2_X1  g0161(.A(new_n361), .B(KEYINPUT17), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n271), .A2(G68), .A3(new_n270), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT77), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n227), .A2(new_n260), .ZN(new_n366));
  OAI22_X1  g0166(.A1(new_n259), .A2(new_n266), .B1(new_n261), .B2(new_n291), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n265), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT11), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n368), .A2(new_n369), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT12), .B1(new_n267), .B2(new_n333), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n211), .A2(G1), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n373), .A2(KEYINPUT12), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n372), .B1(new_n366), .B2(new_n374), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n365), .A2(new_n370), .A3(new_n371), .A4(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(KEYINPUT78), .A2(KEYINPUT14), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n285), .A2(G232), .A3(G1698), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n285), .A2(G226), .A3(new_n286), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G33), .A2(G97), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT75), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(KEYINPUT75), .A2(G33), .A3(G97), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n378), .A2(new_n379), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G238), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n322), .B1(new_n300), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT13), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n389), .B1(new_n385), .B2(new_n386), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT13), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n312), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(KEYINPUT78), .A2(KEYINPUT14), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n377), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT76), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n391), .A2(new_n399), .A3(KEYINPUT13), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT76), .B1(new_n393), .B2(new_n394), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n400), .A2(new_n401), .A3(G179), .A4(new_n395), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n387), .A2(new_n394), .A3(new_n390), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n394), .B1(new_n387), .B2(new_n390), .ZN(new_n404));
  OAI211_X1 g0204(.A(G169), .B(new_n377), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n376), .B1(new_n398), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n376), .ZN(new_n408));
  OAI21_X1  g0208(.A(G200), .B1(new_n403), .B2(new_n404), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n400), .A2(new_n401), .A3(new_n395), .ZN(new_n410));
  INV_X1    g0210(.A(G190), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n408), .B(new_n409), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G20), .A2(G77), .ZN(new_n414));
  XNOR2_X1  g0214(.A(KEYINPUT15), .B(G87), .ZN(new_n415));
  OAI221_X1 g0215(.A(new_n414), .B1(new_n262), .B2(new_n259), .C1(new_n261), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n265), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT72), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n291), .B1(new_n269), .B2(G20), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n271), .A2(new_n419), .B1(new_n291), .B2(new_n267), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n285), .A2(G232), .A3(new_n286), .ZN(new_n422));
  OAI221_X1 g0222(.A(new_n422), .B1(new_n205), .B2(new_n285), .C1(new_n289), .C2(new_n388), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n386), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n299), .B1(new_n301), .B2(G244), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(new_n314), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n425), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n312), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n421), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(G200), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n424), .B2(new_n425), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n427), .A2(new_n411), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n421), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NOR4_X1   g0236(.A1(new_n317), .A2(new_n363), .A3(new_n413), .A4(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT86), .ZN(new_n438));
  INV_X1    g0238(.A(G45), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(G1), .ZN(new_n440));
  NAND2_X1  g0240(.A1(KEYINPUT5), .A2(G41), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(KEYINPUT5), .A2(G41), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n440), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n444), .A2(G257), .A3(new_n295), .ZN(new_n445));
  OAI211_X1 g0245(.A(G244), .B(new_n286), .C1(new_n342), .C2(new_n343), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT4), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n285), .A2(KEYINPUT4), .A3(G244), .A4(new_n286), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n285), .A2(G250), .A3(G1698), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G283), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n448), .A2(new_n449), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n445), .B1(new_n452), .B2(new_n386), .ZN(new_n453));
  OR2_X1    g0253(.A1(KEYINPUT5), .A2(G41), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n441), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n455), .A2(new_n295), .A3(G274), .A4(new_n440), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n453), .A2(new_n314), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n453), .A2(new_n456), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n312), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n259), .A2(new_n291), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n460), .B1(new_n350), .B2(G107), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT6), .ZN(new_n462));
  XOR2_X1   g0262(.A(KEYINPUT81), .B(G97), .Z(new_n463));
  AOI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(new_n205), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G97), .A2(G107), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n206), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT82), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g0268(.A(KEYINPUT81), .B(G97), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT6), .B1(new_n469), .B2(G107), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT82), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(new_n471), .A3(new_n466), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n468), .A2(new_n472), .A3(G20), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n329), .B1(new_n461), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n267), .A2(new_n204), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n373), .A2(G20), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n269), .A2(G33), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n329), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n475), .B1(new_n479), .B2(new_n204), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n457), .B(new_n459), .C1(new_n474), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n350), .A2(G107), .ZN(new_n482));
  INV_X1    g0282(.A(new_n460), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n473), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n265), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n452), .A2(new_n386), .ZN(new_n486));
  INV_X1    g0286(.A(new_n445), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n486), .A2(new_n411), .A3(new_n456), .A4(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n456), .ZN(new_n489));
  AOI211_X1 g0289(.A(new_n489), .B(new_n445), .C1(new_n452), .C2(new_n386), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n488), .B1(new_n490), .B2(G200), .ZN(new_n491));
  INV_X1    g0291(.A(new_n480), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n485), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n481), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT19), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(new_n469), .B2(new_n261), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n285), .A2(new_n260), .A3(G68), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n382), .A2(KEYINPUT19), .A3(new_n383), .ZN(new_n499));
  NOR2_X1   g0299(.A1(G87), .A2(G107), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n499), .A2(new_n260), .B1(new_n469), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n265), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n415), .A2(new_n267), .ZN(new_n503));
  INV_X1    g0303(.A(new_n415), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n478), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT84), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n502), .A2(KEYINPUT84), .A3(new_n503), .A4(new_n505), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n269), .A2(G45), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G250), .ZN(new_n512));
  OAI22_X1  g0312(.A1(new_n386), .A2(new_n512), .B1(new_n298), .B2(new_n511), .ZN(new_n513));
  OAI211_X1 g0313(.A(G244), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n514));
  OAI211_X1 g0314(.A(G238), .B(new_n286), .C1(new_n342), .C2(new_n343), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G116), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n513), .B1(new_n517), .B2(new_n386), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n518), .A2(G169), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n314), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT83), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n518), .A2(KEYINPUT83), .A3(new_n314), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n510), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT85), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n518), .A2(new_n526), .A3(G190), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n526), .B1(new_n518), .B2(G190), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n518), .A2(new_n431), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(G87), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n502), .B(new_n503), .C1(new_n533), .C2(new_n479), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n530), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n525), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n438), .B1(new_n494), .B2(new_n537), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n534), .A2(new_n528), .A3(new_n529), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n539), .A2(new_n532), .B1(new_n510), .B2(new_n524), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n540), .A2(KEYINPUT86), .A3(new_n481), .A4(new_n493), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n267), .A2(KEYINPUT25), .A3(new_n205), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT25), .B1(new_n267), .B2(new_n205), .ZN(new_n543));
  OAI22_X1  g0343(.A1(new_n479), .A2(new_n205), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n260), .B(G87), .C1(new_n342), .C2(new_n343), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT22), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT22), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n285), .A2(new_n547), .A3(new_n260), .A4(G87), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT24), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n260), .A2(G33), .A3(G116), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT88), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT23), .ZN(new_n553));
  AOI21_X1  g0353(.A(KEYINPUT87), .B1(new_n205), .B2(G20), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT23), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT88), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n551), .B(new_n553), .C1(new_n554), .C2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT87), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT23), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n559), .A2(KEYINPUT88), .B1(G20), .B2(new_n205), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n549), .A2(new_n550), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n550), .B1(new_n549), .B2(new_n561), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n265), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT89), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT89), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n566), .B(new_n265), .C1(new_n562), .C2(new_n563), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n544), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n444), .A2(G264), .A3(new_n295), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n569), .A2(new_n456), .ZN(new_n570));
  OAI211_X1 g0370(.A(G257), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n571));
  OAI211_X1 g0371(.A(G250), .B(new_n286), .C1(new_n342), .C2(new_n343), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G33), .A2(G294), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n386), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT90), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(new_n577), .A3(G169), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n314), .B2(new_n576), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n577), .B1(new_n576), .B2(G169), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n568), .A2(new_n581), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n570), .A2(new_n411), .A3(new_n575), .ZN(new_n583));
  AOI21_X1  g0383(.A(G200), .B1(new_n570), .B2(new_n575), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI211_X1 g0385(.A(new_n544), .B(new_n585), .C1(new_n565), .C2(new_n567), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n386), .B1(new_n440), .B2(new_n455), .ZN(new_n587));
  INV_X1    g0387(.A(new_n444), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n386), .A2(new_n298), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n587), .A2(G270), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(G264), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n591));
  OAI211_X1 g0391(.A(G257), .B(new_n286), .C1(new_n342), .C2(new_n343), .ZN(new_n592));
  INV_X1    g0392(.A(G303), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n591), .B(new_n592), .C1(new_n593), .C2(new_n285), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n386), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G190), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n260), .B(new_n451), .C1(new_n469), .C2(G33), .ZN(new_n599));
  INV_X1    g0399(.A(G116), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n264), .A2(new_n218), .B1(G20), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(KEYINPUT20), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT20), .B1(new_n599), .B2(new_n601), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n476), .A2(G116), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n478), .B2(G116), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n596), .A2(G200), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n598), .A2(new_n605), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n607), .B1(new_n603), .B2(new_n604), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n312), .B1(new_n590), .B2(new_n595), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT21), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n610), .A2(KEYINPUT21), .A3(new_n611), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n597), .A2(new_n610), .A3(G179), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n609), .A2(new_n614), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n582), .A2(new_n586), .A3(new_n617), .ZN(new_n618));
  AND4_X1   g0418(.A1(new_n437), .A2(new_n538), .A3(new_n541), .A4(new_n618), .ZN(G372));
  INV_X1    g0419(.A(new_n316), .ZN(new_n620));
  INV_X1    g0420(.A(new_n407), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n412), .B2(new_n430), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n622), .A2(KEYINPUT95), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n362), .B1(new_n622), .B2(KEYINPUT95), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n357), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n307), .A2(new_n311), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n620), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT92), .ZN(new_n628));
  INV_X1    g0428(.A(new_n544), .ZN(new_n629));
  INV_X1    g0429(.A(new_n585), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n549), .A2(new_n561), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT24), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n549), .A2(new_n550), .A3(new_n561), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n566), .B1(new_n634), .B2(new_n265), .ZN(new_n635));
  INV_X1    g0435(.A(new_n567), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n629), .B(new_n630), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n637), .A2(new_n481), .A3(new_n493), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n531), .A2(KEYINPUT91), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n531), .A2(KEYINPUT91), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n530), .A2(new_n639), .A3(new_n535), .A4(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n519), .B1(new_n314), .B2(new_n518), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n510), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n628), .B1(new_n638), .B2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n481), .A2(new_n493), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n639), .A2(new_n640), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n647), .A2(new_n539), .B1(new_n510), .B2(new_n642), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n646), .A2(KEYINPUT92), .A3(new_n637), .A4(new_n648), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(new_n568), .B2(new_n581), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT93), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n579), .A2(new_n580), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n629), .B1(new_n635), .B2(new_n636), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT93), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n645), .A2(new_n649), .A3(new_n652), .A4(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT26), .B1(new_n537), .B2(new_n481), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n457), .B1(new_n490), .B2(G169), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n485), .B2(new_n492), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n662), .A2(new_n663), .A3(new_n643), .A4(new_n641), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT94), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n660), .A2(new_n664), .A3(new_n665), .A4(new_n643), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n660), .A2(new_n664), .A3(new_n643), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT94), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n659), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n437), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n627), .A2(new_n670), .ZN(G369));
  NAND2_X1  g0471(.A1(new_n654), .A2(new_n655), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n373), .A2(new_n260), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n672), .A2(new_n637), .A3(new_n653), .A4(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n582), .A2(new_n679), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n672), .A2(new_n637), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n568), .A2(new_n679), .ZN(new_n685));
  OAI22_X1  g0485(.A1(new_n684), .A2(new_n685), .B1(new_n672), .B2(new_n679), .ZN(new_n686));
  INV_X1    g0486(.A(G330), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n610), .A2(new_n678), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n617), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n653), .A2(new_n688), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n687), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n686), .A2(new_n691), .A3(KEYINPUT96), .ZN(new_n692));
  AOI21_X1  g0492(.A(KEYINPUT96), .B1(new_n686), .B2(new_n691), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n683), .B1(new_n692), .B2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n213), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n469), .A2(new_n600), .A3(new_n500), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n696), .A2(new_n269), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n698), .B1(new_n217), .B2(new_n696), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT28), .Z(new_n700));
  NAND4_X1  g0500(.A1(new_n618), .A2(new_n538), .A3(new_n541), .A4(new_n679), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT31), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n518), .A2(G179), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(new_n576), .A3(new_n596), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n490), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT97), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n569), .A2(new_n456), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n386), .B2(new_n574), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n453), .A2(new_n708), .A3(new_n518), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n590), .A2(new_n595), .A3(G179), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n706), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n705), .B1(new_n711), .B2(KEYINPUT30), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n706), .B(new_n713), .C1(new_n709), .C2(new_n710), .ZN(new_n714));
  AOI211_X1 g0514(.A(new_n702), .B(new_n679), .C1(new_n712), .C2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n711), .A2(KEYINPUT30), .ZN(new_n716));
  INV_X1    g0516(.A(new_n705), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(new_n714), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(KEYINPUT31), .B1(new_n718), .B2(new_n678), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n687), .B1(new_n701), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n669), .A2(new_n679), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT98), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT29), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT98), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n669), .A2(new_n725), .A3(new_n679), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n638), .A2(new_n644), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT99), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(new_n729), .A3(new_n651), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n648), .A2(new_n481), .A3(new_n493), .A4(new_n637), .ZN(new_n731));
  OAI21_X1  g0531(.A(KEYINPUT99), .B1(new_n731), .B2(new_n656), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT26), .B1(new_n644), .B2(new_n481), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n540), .A2(new_n662), .A3(new_n663), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n734), .A2(new_n643), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n678), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT29), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n721), .B1(new_n727), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n700), .B1(new_n739), .B2(G1), .ZN(G364));
  NOR2_X1   g0540(.A1(new_n211), .A2(G20), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n269), .B1(new_n741), .B2(G45), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n696), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n691), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n689), .A2(new_n690), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n745), .B1(G330), .B2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n744), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n213), .A2(G355), .A3(new_n285), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n252), .A2(new_n439), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n695), .A2(new_n285), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(G45), .B2(new_n216), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n749), .B1(G116), .B2(new_n213), .C1(new_n750), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n218), .B1(G20), .B2(new_n312), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n748), .B1(new_n753), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT100), .ZN(new_n760));
  INV_X1    g0560(.A(new_n756), .ZN(new_n761));
  INV_X1    g0561(.A(new_n757), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n260), .A2(new_n314), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n763), .A2(KEYINPUT101), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(KEYINPUT101), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n764), .A2(new_n431), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G190), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n411), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G311), .A2(new_n767), .B1(new_n768), .B2(G322), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n763), .A2(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G190), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OR2_X1    g0572(.A1(KEYINPUT33), .A2(G317), .ZN(new_n773));
  NAND2_X1  g0573(.A1(KEYINPUT33), .A2(G317), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n770), .A2(new_n411), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G326), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G179), .A2(G200), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n260), .B1(new_n779), .B2(G190), .ZN(new_n780));
  INV_X1    g0580(.A(G294), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n777), .A2(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n775), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n431), .A2(G179), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n784), .A2(G20), .A3(new_n411), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n285), .B1(new_n786), .B2(G283), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n784), .A2(G20), .A3(G190), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n779), .A2(G20), .A3(new_n411), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n789), .A2(G303), .B1(new_n791), .B2(G329), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n769), .A2(new_n783), .A3(new_n787), .A4(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(KEYINPUT103), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n793), .A2(KEYINPUT103), .ZN(new_n795));
  INV_X1    g0595(.A(new_n780), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G97), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n790), .A2(new_n331), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT102), .B(KEYINPUT32), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n797), .B1(new_n798), .B2(new_n799), .C1(new_n772), .C2(new_n333), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n777), .B2(new_n266), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n785), .A2(new_n205), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n285), .B1(new_n788), .B2(new_n533), .ZN(new_n804));
  NOR4_X1   g0604(.A1(new_n800), .A2(new_n802), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G58), .A2(new_n768), .B1(new_n767), .B2(G77), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n794), .B(new_n795), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n760), .B1(new_n746), .B2(new_n761), .C1(new_n762), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n747), .A2(new_n808), .ZN(G396));
  AOI21_X1  g0609(.A(new_n679), .B1(new_n418), .B2(new_n420), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n429), .B1(new_n434), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n430), .A2(new_n679), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n723), .A2(new_n726), .A3(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n813), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n669), .A2(new_n679), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n721), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n744), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n818), .B2(new_n817), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n757), .A2(new_n754), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT104), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n748), .B1(new_n823), .B2(new_n291), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G137), .A2(new_n776), .B1(new_n771), .B2(G150), .ZN(new_n825));
  INV_X1    g0625(.A(new_n767), .ZN(new_n826));
  INV_X1    g0626(.A(G143), .ZN(new_n827));
  INV_X1    g0627(.A(new_n768), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n825), .B1(new_n826), .B2(new_n331), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT34), .ZN(new_n830));
  INV_X1    g0630(.A(G132), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n285), .B1(new_n790), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n786), .A2(G68), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n266), .B2(new_n788), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT106), .Z(new_n835));
  AOI211_X1 g0635(.A(new_n832), .B(new_n835), .C1(G58), .C2(new_n796), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n797), .B1(new_n828), .B2(new_n781), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT105), .Z(new_n838));
  INV_X1    g0638(.A(G283), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n772), .A2(new_n839), .B1(new_n777), .B2(new_n593), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n285), .B1(new_n791), .B2(G311), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n841), .B1(new_n533), .B2(new_n785), .C1(new_n205), .C2(new_n788), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n840), .B(new_n842), .C1(G116), .C2(new_n767), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n830), .A2(new_n836), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n824), .B1(new_n762), .B2(new_n844), .C1(new_n815), .C2(new_n755), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n820), .A2(new_n845), .ZN(G384));
  NOR3_X1   g0646(.A1(new_n218), .A2(new_n260), .A3(new_n600), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n468), .A2(new_n472), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT35), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n849), .B2(new_n848), .ZN(new_n851));
  XNOR2_X1  g0651(.A(KEYINPUT107), .B(KEYINPUT36), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n227), .A2(G58), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n217), .A2(new_n854), .A3(G77), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n333), .A2(G50), .ZN(new_n856));
  OAI211_X1 g0656(.A(G1), .B(new_n211), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT108), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n727), .A2(new_n437), .A3(new_n738), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n627), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n376), .A2(new_n678), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n407), .A2(new_n412), .A3(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n376), .B(new_n678), .C1(new_n398), .C2(new_n406), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n816), .B2(new_n812), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n854), .A2(new_n202), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n868), .A2(G20), .B1(G159), .B2(new_n258), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n336), .A2(new_n337), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(G68), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT16), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n265), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n339), .A2(KEYINPUT16), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n355), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n328), .ZN(new_n877));
  INV_X1    g0677(.A(new_n676), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n867), .B1(new_n879), .B2(new_n361), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n350), .A2(new_n227), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT16), .B1(new_n882), .B2(new_n869), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n355), .B1(new_n883), .B2(new_n874), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n877), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n676), .B(KEYINPUT109), .Z(new_n886));
  NAND2_X1  g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n885), .A2(new_n887), .A3(new_n867), .A4(new_n361), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT110), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n881), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n876), .A2(new_n878), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n357), .B2(new_n362), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n892), .A2(new_n895), .A3(KEYINPUT38), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n352), .A2(new_n355), .A3(new_n360), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n898), .A2(new_n356), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n899), .A2(KEYINPUT110), .A3(new_n867), .A4(new_n887), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n888), .A2(new_n889), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n880), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n897), .B1(new_n902), .B2(new_n894), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n896), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n866), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n621), .A2(new_n679), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n896), .A2(new_n903), .A3(KEYINPUT39), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n899), .A2(new_n887), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n890), .B2(new_n891), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n887), .B1(new_n357), .B2(new_n362), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT38), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n902), .A2(new_n894), .A3(new_n897), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n907), .B(new_n908), .C1(new_n916), .C2(KEYINPUT39), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n357), .A2(new_n886), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n905), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n860), .B(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n701), .A2(new_n720), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT40), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n813), .B1(new_n862), .B2(new_n863), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n904), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n922), .A2(new_n924), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n900), .A2(new_n901), .B1(new_n909), .B2(KEYINPUT37), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n897), .B1(new_n928), .B2(new_n912), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n927), .B1(new_n896), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n926), .B1(new_n930), .B2(new_n923), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n437), .A2(new_n922), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n687), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n932), .B2(new_n931), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n921), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n269), .B2(new_n741), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n921), .A2(new_n934), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n853), .B(new_n858), .C1(new_n936), .C2(new_n937), .ZN(G367));
  INV_X1    g0738(.A(new_n739), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n727), .A2(new_n738), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT44), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n662), .A2(new_n678), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n678), .B1(new_n474), .B2(new_n480), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n481), .A2(new_n493), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n941), .B1(new_n683), .B2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n945), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n682), .A2(KEYINPUT44), .A3(new_n947), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n680), .A2(new_n945), .A3(KEYINPUT45), .A4(new_n681), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT45), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n682), .B2(new_n947), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n946), .A2(new_n948), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n692), .A2(new_n693), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n650), .A2(new_n678), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n686), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n691), .ZN(new_n957));
  AND3_X1   g0757(.A1(new_n956), .A2(new_n957), .A3(new_n680), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n957), .B1(new_n956), .B2(new_n680), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n940), .A2(new_n954), .A3(new_n818), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(KEYINPUT112), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT112), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n739), .A2(new_n963), .A3(new_n954), .A4(new_n960), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n939), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(KEYINPUT111), .B(KEYINPUT41), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n696), .B(new_n966), .Z(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n742), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n947), .A2(new_n680), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT42), .Z(new_n971));
  NAND3_X1  g0771(.A1(new_n646), .A2(new_n582), .A3(new_n943), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n678), .B1(new_n972), .B2(new_n481), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT43), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n534), .A2(new_n678), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n643), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(new_n648), .B2(new_n975), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n971), .A2(new_n973), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n974), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n978), .B(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n953), .A2(new_n945), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n969), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n751), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n239), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n758), .B1(new_n213), .B2(new_n415), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n744), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n780), .A2(new_n333), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n777), .A2(new_n827), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n988), .B(new_n989), .C1(G159), .C2(new_n771), .ZN(new_n990));
  INV_X1    g0790(.A(new_n285), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n291), .A2(new_n785), .B1(new_n788), .B2(new_n223), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n991), .B(new_n992), .C1(G137), .C2(new_n791), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G50), .A2(new_n767), .B1(new_n768), .B2(G150), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n990), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n788), .A2(new_n600), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT46), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G294), .B2(new_n771), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n780), .A2(new_n205), .ZN(new_n999));
  INV_X1    g0799(.A(G317), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n991), .B1(new_n790), .B2(new_n1000), .C1(new_n785), .C2(new_n469), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n999), .B(new_n1001), .C1(G311), .C2(new_n776), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G283), .A2(new_n767), .B1(new_n768), .B2(G303), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n998), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n995), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT47), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n987), .B1(new_n1006), .B2(new_n757), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n977), .A2(new_n756), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n983), .A2(new_n1009), .ZN(G387));
  NOR3_X1   g0810(.A1(new_n243), .A2(new_n439), .A3(new_n285), .ZN(new_n1011));
  OR3_X1    g0811(.A1(new_n262), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1012));
  OAI21_X1  g0812(.A(KEYINPUT50), .B1(new_n262), .B2(G50), .ZN(new_n1013));
  AOI21_X1  g0813(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n697), .B1(new_n1015), .B2(new_n991), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n213), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1017), .B(new_n758), .C1(new_n205), .C2(new_n213), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n744), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G50), .A2(new_n768), .B1(new_n767), .B2(G68), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n796), .A2(new_n504), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n777), .B2(new_n331), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n353), .B2(new_n771), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n285), .B1(new_n790), .B2(new_n257), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n788), .A2(new_n291), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(G97), .C2(new_n786), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1020), .A2(new_n1023), .A3(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G311), .A2(new_n771), .B1(new_n776), .B2(G322), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n826), .B2(new_n593), .C1(new_n1000), .C2(new_n828), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT48), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n789), .A2(G294), .B1(new_n796), .B2(G283), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT49), .Z(new_n1035));
  OAI221_X1 g0835(.A(new_n991), .B1(new_n790), .B2(new_n778), .C1(new_n785), .C2(new_n600), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1027), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1019), .B1(new_n1037), .B2(new_n757), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n686), .A2(new_n761), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n960), .A2(new_n743), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n960), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n696), .B1(new_n939), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n739), .A2(new_n960), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1040), .B1(new_n1042), .B2(new_n1043), .ZN(G393));
  NAND2_X1  g0844(.A1(new_n954), .A2(new_n743), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n248), .A2(new_n984), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n758), .B1(new_n213), .B2(new_n469), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n744), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n780), .A2(new_n291), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n789), .A2(new_n227), .B1(new_n791), .B2(G143), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1050), .B(new_n285), .C1(new_n533), .C2(new_n785), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n1049), .B(new_n1051), .C1(G50), .C2(new_n771), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n262), .B2(new_n826), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n768), .A2(G159), .B1(G150), .B2(new_n776), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT51), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n768), .A2(G311), .B1(G317), .B2(new_n776), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT52), .ZN(new_n1057));
  INV_X1    g0857(.A(G322), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n788), .A2(new_n839), .B1(new_n790), .B2(new_n1058), .ZN(new_n1059));
  NOR3_X1   g0859(.A1(new_n1059), .A2(new_n803), .A3(new_n285), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n771), .A2(G303), .B1(G116), .B2(new_n796), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(new_n826), .C2(new_n781), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n1053), .A2(new_n1055), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1048), .B1(new_n1063), .B2(new_n757), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n945), .B2(new_n761), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1045), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n962), .A2(new_n964), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n954), .B1(new_n739), .B2(new_n960), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n696), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1066), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(G390));
  NAND2_X1  g0872(.A1(new_n437), .A2(new_n721), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n859), .A2(new_n627), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n907), .B1(new_n896), .B2(new_n929), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n737), .A2(new_n811), .B1(new_n430), .B2(new_n679), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1075), .B1(new_n1076), .B2(new_n865), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n816), .A2(new_n812), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n907), .B1(new_n1078), .B2(new_n864), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n896), .A2(KEYINPUT39), .A3(new_n903), .ZN(new_n1080));
  AOI21_X1  g0880(.A(KEYINPUT39), .B1(new_n896), .B2(new_n929), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1077), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n721), .A2(new_n924), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n866), .A2(new_n907), .B1(new_n1081), .B2(new_n1080), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1087), .A2(new_n1077), .A3(new_n1084), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n687), .B(new_n813), .C1(new_n701), .C2(new_n720), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1084), .B1(new_n1089), .B2(new_n864), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1078), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n922), .A2(G330), .A3(new_n815), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n865), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n733), .A2(new_n736), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1094), .A2(new_n679), .A3(new_n811), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1093), .A2(new_n1095), .A3(new_n812), .A4(new_n1084), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1074), .A2(new_n1086), .A3(new_n1088), .A4(new_n1097), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n859), .A2(new_n1097), .A3(new_n627), .A4(new_n1073), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1087), .A2(new_n1077), .A3(new_n1084), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1084), .B1(new_n1087), .B2(new_n1077), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1098), .A2(new_n696), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT116), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1086), .A2(new_n743), .A3(new_n1088), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT113), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1086), .A2(KEYINPUT113), .A3(new_n743), .A4(new_n1088), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n754), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n991), .B1(new_n791), .B2(G125), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n266), .B2(new_n785), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(KEYINPUT114), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(KEYINPUT54), .B(G143), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1113), .B1(new_n826), .B2(new_n1114), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n828), .A2(new_n831), .B1(new_n1112), .B2(KEYINPUT114), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n788), .A2(new_n257), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT53), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(G128), .A2(new_n776), .B1(new_n771), .B2(G137), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1118), .B(new_n1119), .C1(new_n331), .C2(new_n780), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n1115), .A2(new_n1116), .A3(new_n1120), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n600), .A2(new_n828), .B1(new_n826), .B2(new_n469), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G107), .A2(new_n771), .B1(new_n776), .B2(G283), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1049), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n791), .A2(G294), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1123), .A2(new_n833), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n991), .B1(new_n788), .B2(new_n533), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT115), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n1122), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n757), .B1(new_n1121), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n748), .B1(new_n823), .B2(new_n262), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1110), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1104), .B1(new_n1109), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1132), .ZN(new_n1134));
  AOI211_X1 g0934(.A(KEYINPUT116), .B(new_n1134), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1103), .B1(new_n1133), .B2(new_n1135), .ZN(G378));
  INV_X1    g0936(.A(KEYINPUT119), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n1100), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n859), .A2(new_n627), .A3(new_n1073), .ZN(new_n1139));
  OAI21_X1  g0939(.A(KEYINPUT57), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n276), .A2(new_n878), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n626), .A2(new_n316), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n317), .A2(new_n276), .A3(new_n878), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1142), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n864), .A2(new_n815), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n701), .B2(new_n720), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n914), .B2(new_n915), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1153), .A2(KEYINPUT40), .B1(new_n904), .B2(new_n925), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1150), .B1(new_n1154), .B2(new_n687), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n896), .A2(new_n929), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n923), .B1(new_n1156), .B2(new_n1152), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n896), .B2(new_n903), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1149), .B(G330), .C1(new_n1157), .C2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1155), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(KEYINPUT118), .B1(new_n1161), .B2(new_n920), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1160), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1149), .B1(new_n931), .B2(G330), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n920), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n918), .B1(new_n1082), .B2(new_n907), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1155), .A2(new_n905), .A3(new_n1166), .A4(new_n1160), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1162), .B1(new_n1168), .B2(KEYINPUT118), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1137), .B1(new_n1140), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1168), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1069), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1163), .A2(new_n1164), .A3(new_n920), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1155), .A2(new_n1160), .B1(new_n1166), .B2(new_n905), .ZN(new_n1175));
  OAI21_X1  g0975(.A(KEYINPUT118), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1162), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1172), .B1(new_n1098), .B2(new_n1074), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1178), .A2(KEYINPUT119), .A3(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1170), .A2(new_n1173), .A3(new_n1180), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(G128), .A2(new_n768), .B1(new_n767), .B2(G137), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NOR3_X1   g0983(.A1(new_n788), .A2(new_n1114), .A3(KEYINPUT117), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(G125), .B2(new_n776), .ZN(new_n1185));
  OAI21_X1  g0985(.A(KEYINPUT117), .B1(new_n788), .B2(new_n1114), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n771), .A2(G132), .B1(G150), .B2(new_n796), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  OR3_X1    g0988(.A1(new_n1183), .A2(KEYINPUT59), .A3(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(KEYINPUT59), .B1(new_n1183), .B2(new_n1188), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n786), .A2(G159), .ZN(new_n1191));
  AOI211_X1 g0991(.A(G33), .B(G41), .C1(new_n791), .C2(G124), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n777), .A2(new_n600), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n988), .B(new_n1194), .C1(G97), .C2(new_n771), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n785), .A2(new_n223), .B1(new_n839), .B2(new_n790), .ZN(new_n1196));
  NOR4_X1   g0996(.A1(new_n1196), .A2(new_n1025), .A3(G41), .A4(new_n285), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(G107), .A2(new_n768), .B1(new_n767), .B2(new_n504), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT58), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n266), .B1(new_n342), .B2(G41), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1193), .A2(new_n1201), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n757), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n748), .B1(new_n266), .B2(new_n821), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1205), .B(new_n1206), .C1(new_n1149), .C2(new_n755), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n1168), .B2(new_n743), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1181), .A2(new_n1209), .ZN(G375));
  INV_X1    g1010(.A(new_n1097), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1139), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1212), .A2(new_n967), .A3(new_n1099), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n789), .A2(G159), .B1(new_n791), .B2(G128), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n991), .B1(new_n786), .B2(G58), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(new_n266), .C2(new_n780), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n831), .A2(new_n777), .B1(new_n772), .B2(new_n1114), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G137), .B2(new_n768), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT121), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1216), .B(new_n1219), .C1(G150), .C2(new_n767), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n205), .A2(new_n826), .B1(new_n828), .B2(new_n839), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G116), .A2(new_n771), .B1(new_n776), .B2(G294), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n791), .A2(G303), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n789), .A2(G97), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1222), .A2(new_n1021), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n285), .B1(new_n786), .B2(G77), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT120), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1221), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n757), .B1(new_n1220), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n748), .B1(new_n823), .B2(new_n333), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n865), .B2(new_n754), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1097), .B2(new_n743), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1213), .A2(new_n1233), .ZN(G381));
  OR3_X1    g1034(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1235), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(KEYINPUT122), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1109), .A2(new_n1103), .A3(new_n1132), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1181), .A2(new_n1209), .A3(new_n1238), .ZN(new_n1239));
  OR2_X1    g1039(.A1(new_n1237), .A2(new_n1239), .ZN(G407));
  OAI211_X1 g1040(.A(G407), .B(G213), .C1(G343), .C2(new_n1239), .ZN(G409));
  NAND3_X1  g1041(.A1(G378), .A2(new_n1181), .A3(new_n1209), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1207), .B1(new_n1169), .B2(new_n742), .C1(new_n968), .C2(new_n1171), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1238), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n677), .A2(G213), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1099), .A2(KEYINPUT60), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1212), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1139), .A2(KEYINPUT60), .A3(new_n1211), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1249), .A2(new_n696), .A3(new_n1250), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1251), .A2(G384), .A3(new_n1233), .ZN(new_n1252));
  AOI21_X1  g1052(.A(G384), .B1(new_n1251), .B2(new_n1233), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n677), .A2(G213), .A3(G2897), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1254), .A2(KEYINPUT123), .A3(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1254), .A2(KEYINPUT123), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1255), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1253), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1251), .A2(G384), .A3(new_n1233), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT123), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1259), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1256), .B1(new_n1258), .B2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT61), .B1(new_n1247), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT125), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT62), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1245), .A2(new_n1246), .A3(new_n1269), .A4(new_n1254), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1242), .A2(new_n1244), .B1(G213), .B2(new_n677), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1271), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1273), .A2(new_n1274), .A3(new_n1269), .A4(new_n1254), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1266), .A2(new_n1272), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G387), .A2(new_n1071), .ZN(new_n1277));
  XOR2_X1   g1077(.A(G393), .B(G396), .Z(new_n1278));
  NAND3_X1  g1078(.A1(new_n983), .A2(new_n1009), .A3(G390), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1278), .ZN(new_n1281));
  AOI21_X1  g1081(.A(G390), .B1(new_n983), .B2(new_n1009), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1009), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n1283), .B(new_n1071), .C1(new_n969), .C2(new_n982), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1281), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1280), .A2(new_n1285), .A3(KEYINPUT126), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT126), .B1(new_n1280), .B2(new_n1285), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1276), .A2(new_n1288), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1280), .A2(new_n1285), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT61), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1262), .A2(new_n1263), .A3(new_n1259), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1255), .B1(new_n1254), .B2(KEYINPUT123), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1292), .B1(new_n1293), .B2(new_n1257), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1290), .B(new_n1291), .C1(new_n1273), .C2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT63), .B1(new_n1273), .B2(new_n1254), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1245), .A2(KEYINPUT63), .A3(new_n1246), .A4(new_n1254), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(KEYINPUT124), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT124), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1273), .A2(new_n1300), .A3(KEYINPUT63), .A4(new_n1254), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1297), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1289), .A2(new_n1303), .ZN(G405));
  INV_X1    g1104(.A(KEYINPUT127), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G375), .A2(new_n1238), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1242), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1254), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1306), .A2(new_n1242), .A3(new_n1262), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1280), .A2(new_n1285), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT126), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1280), .A2(new_n1285), .A3(KEYINPUT126), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1305), .B1(new_n1310), .B2(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1288), .A2(KEYINPUT127), .A3(new_n1308), .A4(new_n1309), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1310), .A2(new_n1315), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1316), .A2(new_n1317), .A3(new_n1318), .ZN(G402));
endmodule


