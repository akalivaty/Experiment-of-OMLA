//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1228, new_n1229, new_n1230;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  OR2_X1    g0006(.A1(new_n206), .A2(KEYINPUT64), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(KEYINPUT64), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI211_X1 g0022(.A(new_n216), .B(new_n222), .C1(G116), .C2(G270), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(new_n208), .B2(new_n207), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n201), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n212), .B(new_n225), .C1(new_n228), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(new_n219), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT2), .ZN(new_n235));
  INV_X1    g0035(.A(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G264), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n239), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n218), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT65), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n202), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G107), .ZN(new_n247));
  INV_X1    g0047(.A(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n245), .B(new_n249), .ZN(G351));
  AOI21_X1  g0050(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G232), .A3(G1698), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n257), .B1(new_n259), .B2(new_n236), .ZN(new_n260));
  INV_X1    g0060(.A(G97), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n253), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n251), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  INV_X1    g0064(.A(G45), .ZN(new_n265));
  AOI21_X1  g0065(.A(G1), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G274), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n251), .A2(new_n266), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G238), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n263), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT13), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT73), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT13), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n263), .A2(new_n273), .A3(new_n267), .A4(new_n269), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n271), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n270), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G169), .ZN(new_n278));
  OAI21_X1  g0078(.A(KEYINPUT14), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n271), .A2(G179), .A3(new_n274), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT14), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n275), .A2(new_n281), .A3(G169), .A4(new_n276), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G1), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT70), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n284), .A2(KEYINPUT70), .A3(G13), .A4(G20), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n290), .A2(KEYINPUT74), .A3(KEYINPUT12), .A4(new_n214), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT74), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT12), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n290), .A2(new_n214), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n294), .B1(new_n292), .B2(new_n293), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n226), .B1(new_n206), .B2(new_n253), .ZN(new_n296));
  AOI211_X1 g0096(.A(new_n296), .B(new_n290), .C1(new_n284), .C2(G20), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n291), .B(new_n295), .C1(new_n298), .C2(new_n214), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n253), .A2(G20), .ZN(new_n300));
  NOR2_X1   g0100(.A1(G20), .A2(G33), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n300), .A2(G77), .B1(new_n301), .B2(G50), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(new_n227), .B2(G68), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n296), .ZN(new_n304));
  XOR2_X1   g0104(.A(new_n304), .B(KEYINPUT11), .Z(new_n305));
  NOR2_X1   g0105(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n283), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  OR2_X1    g0109(.A1(KEYINPUT66), .A2(G226), .ZN(new_n310));
  NAND2_X1  g0110(.A1(KEYINPUT66), .A2(G226), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n268), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G222), .ZN(new_n313));
  INV_X1    g0113(.A(G77), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n259), .A2(new_n313), .B1(new_n314), .B2(new_n256), .ZN(new_n315));
  AND2_X1   g0115(.A1(KEYINPUT3), .A2(G33), .ZN(new_n316));
  NOR2_X1   g0116(.A1(KEYINPUT3), .A2(G33), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(new_n258), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n315), .B1(G223), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n251), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n267), .B(new_n312), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(G179), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n218), .A2(KEYINPUT67), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT68), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G58), .ZN(new_n326));
  OAI211_X1 g0126(.A(KEYINPUT8), .B(new_n324), .C1(new_n326), .C2(KEYINPUT67), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n326), .A2(KEYINPUT8), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n329), .A2(new_n300), .B1(G150), .B2(new_n301), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n330), .A2(KEYINPUT69), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n203), .A2(G20), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(KEYINPUT69), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n334), .A2(new_n296), .B1(new_n202), .B2(new_n290), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n297), .A2(G50), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI211_X1 g0137(.A(new_n323), .B(new_n337), .C1(new_n278), .C2(new_n322), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n335), .A2(new_n336), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT9), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G190), .ZN(new_n342));
  OR2_X1    g0142(.A1(new_n322), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n335), .A2(KEYINPUT9), .A3(new_n336), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n322), .A2(G200), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n341), .A2(new_n343), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT10), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n344), .A2(new_n345), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT10), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n348), .A2(new_n349), .A3(new_n343), .A4(new_n341), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n338), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n267), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(new_n268), .B2(G244), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n256), .A2(G232), .A3(new_n258), .ZN(new_n354));
  INV_X1    g0154(.A(G107), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n256), .A2(G1698), .ZN(new_n356));
  OAI221_X1 g0156(.A(new_n354), .B1(new_n355), .B2(new_n256), .C1(new_n356), .C2(new_n215), .ZN(new_n357));
  XOR2_X1   g0157(.A(new_n357), .B(KEYINPUT71), .Z(new_n358));
  OAI21_X1  g0158(.A(new_n353), .B1(new_n358), .B2(new_n321), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n359), .A2(G179), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n278), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n290), .A2(new_n314), .ZN(new_n362));
  XOR2_X1   g0162(.A(KEYINPUT15), .B(G87), .Z(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n300), .ZN(new_n365));
  INV_X1    g0165(.A(new_n301), .ZN(new_n366));
  XNOR2_X1  g0166(.A(KEYINPUT8), .B(G58), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n364), .A2(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n227), .A2(new_n314), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n296), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n362), .B(new_n370), .C1(new_n298), .C2(new_n314), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n360), .A2(new_n361), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n371), .B1(new_n359), .B2(G200), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n342), .B2(new_n359), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n351), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT72), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n351), .A2(KEYINPUT72), .A3(new_n372), .A4(new_n374), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n309), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n271), .A2(G190), .A3(new_n274), .ZN(new_n380));
  INV_X1    g0180(.A(G200), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n306), .B(new_n380), .C1(new_n277), .C2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT18), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n329), .A2(new_n289), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n297), .B2(new_n329), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT7), .B1(new_n318), .B2(new_n227), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n254), .A2(KEYINPUT7), .A3(new_n227), .A4(new_n255), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(G68), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT75), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT67), .B(G58), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n229), .B1(new_n392), .B2(new_n214), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n393), .A2(G20), .B1(G159), .B2(new_n301), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n254), .A2(new_n227), .A3(new_n255), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT7), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n388), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT75), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n399), .A3(G68), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n391), .A2(KEYINPUT16), .A3(new_n394), .A4(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT76), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n401), .B(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n394), .A2(new_n390), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT16), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n403), .A2(KEYINPUT77), .A3(new_n296), .A4(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n399), .B1(new_n398), .B2(G68), .ZN(new_n408));
  AOI211_X1 g0208(.A(KEYINPUT75), .B(new_n214), .C1(new_n397), .C2(new_n388), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n410), .A2(new_n402), .A3(KEYINPUT16), .A4(new_n394), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n401), .A2(KEYINPUT76), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n411), .A2(new_n412), .A3(new_n296), .A4(new_n406), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT77), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n386), .B1(new_n407), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n318), .A2(G1698), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G223), .ZN(new_n418));
  OAI221_X1 g0218(.A(new_n418), .B1(new_n253), .B2(new_n220), .C1(new_n236), .C2(new_n356), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n352), .B1(new_n419), .B2(new_n251), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n268), .A2(G232), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G179), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(G169), .B2(new_n422), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n383), .B1(new_n416), .B2(new_n425), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n413), .A2(new_n414), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n413), .A2(new_n414), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n385), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n422), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(G179), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n278), .B2(new_n430), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n429), .A2(KEYINPUT18), .A3(new_n432), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n420), .A2(new_n342), .A3(new_n421), .ZN(new_n434));
  AOI21_X1  g0234(.A(G200), .B1(new_n420), .B2(new_n421), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n385), .B(new_n437), .C1(new_n427), .C2(new_n428), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT17), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT17), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n416), .A2(new_n440), .A3(new_n437), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n426), .A2(new_n433), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n382), .B1(new_n442), .B2(KEYINPUT78), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n443), .B1(KEYINPUT78), .B2(new_n442), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n379), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n296), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n289), .B(new_n447), .C1(G1), .C2(new_n253), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n448), .B(KEYINPUT80), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G107), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n289), .A2(G107), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT25), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n256), .A2(KEYINPUT89), .A3(new_n227), .A4(G87), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n453), .B(KEYINPUT22), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n227), .A2(G107), .ZN(new_n455));
  XNOR2_X1  g0255(.A(new_n455), .B(KEYINPUT23), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n454), .B(new_n456), .C1(new_n248), .C2(new_n365), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT24), .ZN(new_n458));
  XNOR2_X1  g0258(.A(new_n457), .B(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n450), .B(new_n452), .C1(new_n459), .C2(new_n447), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n265), .A2(G1), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT81), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n461), .B(new_n462), .C1(KEYINPUT5), .C2(new_n264), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n284), .B(G45), .C1(new_n264), .C2(KEYINPUT5), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT81), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n264), .A2(KEYINPUT5), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n467), .A2(new_n321), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G264), .ZN(new_n469));
  INV_X1    g0269(.A(G257), .ZN(new_n470));
  OAI22_X1  g0270(.A1(new_n221), .A2(new_n259), .B1(new_n356), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(G294), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n253), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n251), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n463), .A2(new_n465), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n475), .A2(G274), .A3(new_n321), .A4(new_n466), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n469), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n278), .ZN(new_n478));
  INV_X1    g0278(.A(new_n477), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n423), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n460), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n256), .A2(new_n227), .A3(G68), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n365), .A2(new_n261), .ZN(new_n483));
  XNOR2_X1  g0283(.A(KEYINPUT83), .B(G87), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n484), .A2(G97), .A3(G107), .ZN(new_n485));
  AOI21_X1  g0285(.A(G20), .B1(new_n262), .B2(KEYINPUT19), .ZN(new_n486));
  OAI221_X1 g0286(.A(new_n482), .B1(new_n483), .B2(KEYINPUT19), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n487), .A2(new_n296), .B1(new_n290), .B2(new_n364), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT80), .ZN(new_n489));
  XNOR2_X1  g0289(.A(new_n448), .B(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n488), .B1(new_n490), .B2(new_n364), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT84), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OR3_X1    g0293(.A1(new_n251), .A2(new_n221), .A3(new_n461), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n461), .A2(G274), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT82), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n461), .A2(KEYINPUT82), .A3(G274), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n256), .A2(G238), .A3(new_n258), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n256), .A2(G244), .A3(G1698), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G116), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n500), .B1(new_n251), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n278), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n423), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n488), .B(KEYINPUT84), .C1(new_n490), .C2(new_n364), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n493), .A2(new_n507), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n488), .B1(new_n490), .B2(new_n220), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(G190), .B2(new_n505), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n381), .B2(new_n505), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n481), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n479), .A2(new_n381), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n477), .A2(new_n342), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n460), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  XNOR2_X1  g0317(.A(G97), .B(G107), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT6), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(G97), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(KEYINPUT79), .ZN(new_n522));
  MUX2_X1   g0322(.A(new_n518), .B(new_n521), .S(new_n522), .Z(new_n523));
  AOI22_X1  g0323(.A1(new_n523), .A2(G20), .B1(G107), .B2(new_n398), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n314), .B2(new_n366), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n525), .A2(new_n296), .B1(G97), .B2(new_n449), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n290), .A2(new_n261), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT4), .ZN(new_n529));
  INV_X1    g0329(.A(G244), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n529), .B1(new_n259), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n417), .A2(KEYINPUT4), .A3(G244), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n319), .A2(G250), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G283), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n531), .A2(new_n532), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n251), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n468), .A2(G257), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n536), .A2(new_n537), .A3(new_n476), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G179), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n536), .A2(new_n537), .A3(new_n476), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G169), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n528), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n540), .A2(G200), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n342), .B2(new_n540), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n543), .B1(new_n545), .B2(new_n528), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n517), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n534), .B(new_n227), .C1(G33), .C2(new_n261), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n548), .B(new_n296), .C1(new_n227), .C2(G116), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT20), .ZN(new_n550));
  OR3_X1    g0350(.A1(new_n549), .A2(KEYINPUT86), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(KEYINPUT86), .B1(new_n549), .B2(new_n550), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n550), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n290), .A2(new_n248), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n554), .B(new_n555), .C1(new_n248), .C2(new_n448), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n256), .A2(G264), .A3(G1698), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n318), .A2(G303), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n557), .B(new_n558), .C1(new_n259), .C2(new_n470), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n251), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n467), .A2(G270), .A3(new_n321), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n476), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT85), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT85), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n560), .A2(new_n476), .A3(new_n564), .A4(new_n561), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n556), .B1(new_n566), .B2(G200), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n342), .B2(new_n566), .ZN(new_n568));
  XNOR2_X1  g0368(.A(new_n568), .B(KEYINPUT88), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n278), .B1(new_n563), .B2(new_n565), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n570), .A2(KEYINPUT21), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n562), .A2(new_n423), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n556), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n570), .A2(new_n556), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT21), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT87), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT87), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n574), .A2(new_n578), .A3(new_n575), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n573), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n569), .A2(new_n580), .ZN(new_n581));
  AND4_X1   g0381(.A1(new_n446), .A2(new_n514), .A3(new_n547), .A4(new_n581), .ZN(G372));
  NAND4_X1  g0382(.A1(new_n481), .A2(new_n579), .A3(new_n573), .A4(new_n577), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n504), .A2(new_n251), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT90), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n504), .A2(KEYINPUT90), .A3(new_n251), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n500), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n512), .B1(new_n381), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n500), .ZN(new_n590));
  INV_X1    g0390(.A(new_n587), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT90), .B1(new_n504), .B2(new_n251), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n278), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n493), .A2(new_n508), .A3(new_n509), .A4(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n547), .A2(new_n583), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n542), .A2(KEYINPUT91), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT91), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n539), .A2(new_n599), .A3(new_n541), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n601), .A2(new_n528), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT26), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n603), .A3(new_n596), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n513), .A2(new_n510), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT26), .B1(new_n605), .B2(new_n543), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n597), .A2(new_n604), .A3(new_n595), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n446), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT92), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT18), .B1(new_n429), .B2(new_n432), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n416), .A2(new_n383), .A3(new_n425), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n426), .A2(new_n433), .A3(KEYINPUT92), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n439), .A2(new_n441), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n372), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n309), .B1(new_n617), .B2(new_n382), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n614), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n347), .A2(new_n350), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n338), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n608), .A2(new_n621), .ZN(G369));
  INV_X1    g0422(.A(G13), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n623), .A2(G20), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n284), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n625), .A2(KEYINPUT27), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(KEYINPUT27), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(G213), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(G343), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n556), .A2(new_n630), .ZN(new_n631));
  MUX2_X1   g0431(.A(new_n580), .B(new_n581), .S(new_n631), .Z(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(G330), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n460), .A2(new_n630), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n481), .B1(new_n517), .B2(new_n635), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n481), .A2(new_n630), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n630), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n580), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(new_n637), .A3(new_n636), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n637), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n639), .A2(new_n644), .ZN(G399));
  INV_X1    g0445(.A(new_n210), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(G41), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n485), .A2(new_n248), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n647), .A2(new_n284), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n231), .B2(new_n647), .ZN(new_n650));
  XOR2_X1   g0450(.A(new_n650), .B(KEYINPUT28), .Z(new_n651));
  AOI21_X1  g0451(.A(G179), .B1(new_n593), .B2(KEYINPUT93), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT93), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n588), .A2(new_n653), .ZN(new_n654));
  AND4_X1   g0454(.A1(KEYINPUT94), .A2(new_n652), .A3(new_n566), .A4(new_n654), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n563), .A2(new_n565), .B1(new_n588), .B2(new_n653), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT94), .B1(new_n656), .B2(new_n652), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n477), .B(new_n540), .C1(new_n655), .C2(new_n657), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n505), .A2(new_n474), .A3(new_n469), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n538), .A2(new_n659), .A3(new_n572), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT30), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  AND4_X1   g0462(.A1(KEYINPUT95), .A2(new_n662), .A3(KEYINPUT31), .A4(new_n630), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n640), .B1(new_n658), .B2(new_n661), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT95), .B1(new_n664), .B2(KEYINPUT31), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n662), .A2(new_n630), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT31), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(KEYINPUT96), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n662), .A2(KEYINPUT31), .A3(new_n630), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT95), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n664), .A2(KEYINPUT95), .A3(KEYINPUT31), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n673), .A2(new_n669), .A3(KEYINPUT96), .A4(new_n674), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n581), .A2(new_n514), .A3(new_n547), .A4(new_n640), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(G330), .B1(new_n670), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n607), .A2(new_n640), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(KEYINPUT29), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT29), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n605), .A2(KEYINPUT26), .A3(new_n543), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n596), .A2(new_n528), .A3(new_n601), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n682), .B1(new_n683), .B2(KEYINPUT26), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n684), .A2(new_n597), .A3(new_n595), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n681), .B1(new_n685), .B2(new_n640), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n678), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT97), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n688), .B(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n651), .B1(new_n690), .B2(G1), .ZN(G364));
  INV_X1    g0491(.A(new_n647), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n284), .B1(new_n624), .B2(G45), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT98), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n634), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(G330), .B2(new_n632), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n226), .B1(G20), .B2(new_n278), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n227), .A2(G179), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(new_n342), .A3(G200), .ZN(new_n700));
  INV_X1    g0500(.A(G283), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n318), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n227), .A2(new_n423), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G200), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT102), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G190), .ZN(new_n706));
  XNOR2_X1  g0506(.A(KEYINPUT33), .B(G317), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n702), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NOR4_X1   g0508(.A1(new_n227), .A2(new_n423), .A3(new_n342), .A4(G200), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT100), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n709), .A2(KEYINPUT100), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G322), .ZN(new_n715));
  NOR2_X1   g0515(.A1(G190), .A2(G200), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n699), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT104), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n703), .A2(KEYINPUT101), .A3(new_n716), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT101), .B1(new_n703), .B2(new_n716), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n719), .A2(G329), .B1(new_n724), .B2(G311), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n708), .A2(new_n715), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n705), .A2(new_n342), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n342), .A2(G179), .A3(G200), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n227), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n727), .A2(G326), .B1(G294), .B2(new_n730), .ZN(new_n731));
  XOR2_X1   g0531(.A(new_n731), .B(KEYINPUT103), .Z(new_n732));
  NAND3_X1  g0532(.A1(new_n699), .A2(G190), .A3(G200), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI211_X1 g0534(.A(new_n726), .B(new_n732), .C1(G303), .C2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n318), .B1(new_n724), .B2(G77), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n484), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n736), .B(new_n737), .C1(new_n713), .C2(new_n392), .ZN(new_n738));
  INV_X1    g0538(.A(new_n717), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G159), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n740), .A2(KEYINPUT32), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n700), .A2(new_n355), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n742), .B1(new_n740), .B2(KEYINPUT32), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n727), .ZN(new_n745));
  INV_X1    g0545(.A(new_n706), .ZN(new_n746));
  OAI221_X1 g0546(.A(new_n744), .B1(new_n745), .B2(new_n202), .C1(new_n214), .C2(new_n746), .ZN(new_n747));
  AOI211_X1 g0547(.A(new_n738), .B(new_n747), .C1(G97), .C2(new_n730), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n698), .B1(new_n735), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n749), .B1(new_n632), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n231), .A2(new_n265), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n318), .B(new_n755), .C1(new_n245), .C2(new_n265), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n256), .A2(G355), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n756), .A2(new_n210), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n752), .A2(new_n698), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n758), .B(new_n759), .C1(new_n248), .C2(new_n210), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(new_n695), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT99), .Z(new_n762));
  OAI21_X1  g0562(.A(new_n697), .B1(new_n754), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT105), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(G396));
  NAND2_X1  g0565(.A1(new_n371), .A2(new_n630), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n374), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n617), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n372), .A2(new_n630), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n679), .B(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(new_n678), .ZN(new_n772));
  INV_X1    g0572(.A(new_n695), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G137), .A2(new_n727), .B1(new_n706), .B2(G150), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT106), .Z(new_n776));
  INV_X1    g0576(.A(G143), .ZN(new_n777));
  INV_X1    g0577(.A(G159), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n776), .B1(new_n777), .B2(new_n713), .C1(new_n778), .C2(new_n723), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT34), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n256), .B1(new_n733), .B2(new_n202), .C1(new_n729), .C2(new_n392), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(new_n719), .B2(G132), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n780), .B(new_n782), .C1(new_n214), .C2(new_n700), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n700), .A2(new_n220), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n713), .A2(new_n472), .B1(new_n248), .B2(new_n723), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(G311), .B2(new_n719), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n256), .B1(new_n730), .B2(G97), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(new_n355), .B2(new_n733), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(new_n706), .B2(G283), .ZN(new_n789));
  INV_X1    g0589(.A(G303), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n786), .B(new_n789), .C1(new_n790), .C2(new_n745), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n783), .B1(new_n784), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n773), .B1(new_n792), .B2(new_n698), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n698), .A2(new_n750), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n793), .B1(G77), .B2(new_n795), .C1(new_n770), .C2(new_n751), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n774), .A2(new_n796), .ZN(G384));
  XNOR2_X1  g0597(.A(new_n413), .B(KEYINPUT77), .ZN(new_n798));
  INV_X1    g0598(.A(new_n628), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n798), .A2(new_n386), .B1(new_n432), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT37), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n800), .A2(new_n801), .A3(new_n438), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n431), .B(new_n628), .C1(new_n430), .C2(new_n278), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n410), .A2(new_n394), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n405), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n403), .A2(new_n296), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n385), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n438), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(KEYINPUT37), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n802), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n807), .A2(new_n799), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n811), .B(KEYINPUT38), .C1(new_n442), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n407), .A2(new_n415), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n814), .A2(new_n385), .B1(new_n425), .B2(new_n628), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n386), .B(new_n436), .C1(new_n407), .C2(new_n415), .ZN(new_n816));
  OAI21_X1  g0616(.A(KEYINPUT37), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n817), .A2(new_n802), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n612), .A2(new_n615), .A3(new_n613), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n429), .A2(new_n799), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n818), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n813), .B1(new_n822), .B2(KEYINPUT38), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n676), .A2(new_n669), .A3(new_n671), .ZN(new_n824));
  AND3_X1   g0624(.A1(new_n283), .A2(KEYINPUT107), .A3(new_n307), .ZN(new_n825));
  AOI21_X1  g0625(.A(KEYINPUT107), .B1(new_n283), .B2(new_n307), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n382), .B1(new_n306), .B2(new_n640), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n309), .A2(new_n630), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AND3_X1   g0629(.A1(new_n824), .A2(new_n829), .A3(new_n770), .ZN(new_n830));
  AND3_X1   g0630(.A1(new_n823), .A2(new_n830), .A3(KEYINPUT40), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT38), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n426), .A2(new_n433), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n812), .B1(new_n833), .B2(new_n615), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n801), .B1(new_n438), .B2(new_n808), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n815), .A2(new_n816), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n835), .B1(new_n836), .B2(new_n801), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n832), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT108), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n838), .A2(new_n839), .A3(new_n813), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n834), .A2(new_n837), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n841), .A2(KEYINPUT108), .A3(KEYINPUT38), .ZN(new_n842));
  AND3_X1   g0642(.A1(new_n840), .A2(KEYINPUT109), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(KEYINPUT109), .B1(new_n840), .B2(new_n842), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n830), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT40), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n831), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n379), .A2(new_n444), .A3(new_n824), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(G330), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n679), .A2(new_n768), .B1(new_n372), .B2(new_n630), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n851), .A2(new_n829), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n843), .B2(new_n844), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n840), .A2(new_n842), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT39), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n823), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n825), .A2(new_n826), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n640), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n855), .A2(new_n857), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n614), .A2(new_n799), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n853), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n379), .B(new_n444), .C1(new_n680), .C2(new_n686), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n621), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n864), .B(new_n866), .Z(new_n867));
  XNOR2_X1  g0667(.A(new_n850), .B(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n284), .B2(new_n624), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n248), .B1(new_n523), .B2(KEYINPUT35), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n870), .B(new_n228), .C1(KEYINPUT35), .C2(new_n523), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT36), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n231), .B1(new_n392), .B2(new_n214), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n873), .A2(new_n314), .B1(G50), .B2(new_n214), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n874), .A2(G1), .A3(new_n623), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n869), .A2(new_n872), .A3(new_n875), .ZN(G367));
  NAND2_X1  g0676(.A1(new_n602), .A2(new_n630), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n640), .B1(new_n526), .B2(new_n527), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n546), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n639), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n511), .A2(new_n630), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n596), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n595), .B2(new_n884), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT43), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n881), .A2(new_n642), .ZN(new_n888));
  XNOR2_X1  g0688(.A(KEYINPUT111), .B(KEYINPUT42), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n888), .B(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n543), .B1(new_n881), .B2(new_n481), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT110), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n890), .B1(new_n892), .B2(new_n630), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n883), .A2(new_n887), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n883), .B1(new_n893), .B2(new_n887), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n886), .A2(KEYINPUT43), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  OR3_X1    g0697(.A1(new_n894), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n897), .B1(new_n894), .B2(new_n895), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n647), .B(KEYINPUT41), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n643), .A2(new_n881), .ZN(new_n902));
  XOR2_X1   g0702(.A(KEYINPUT112), .B(KEYINPUT44), .Z(new_n903));
  XNOR2_X1  g0703(.A(new_n902), .B(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n643), .A2(new_n881), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT45), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n904), .A2(new_n639), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n639), .B1(new_n906), .B2(new_n904), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT113), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n908), .A2(KEYINPUT113), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n638), .B(new_n641), .Z(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n634), .B2(KEYINPUT114), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT114), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n633), .B(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n912), .B1(new_n914), .B2(new_n911), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n909), .A2(new_n910), .A3(new_n690), .A4(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n901), .B1(new_n916), .B2(new_n690), .ZN(new_n917));
  INV_X1    g0717(.A(new_n693), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n898), .B(new_n899), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(G317), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n318), .B1(new_n717), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n700), .A2(new_n261), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(G107), .B2(new_n730), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n746), .B2(new_n472), .ZN(new_n924));
  AOI211_X1 g0724(.A(new_n921), .B(new_n924), .C1(G311), .C2(new_n727), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT46), .B1(new_n734), .B2(G116), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n734), .A2(KEYINPUT46), .A3(G116), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n926), .B(new_n927), .C1(new_n724), .C2(G283), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n925), .B(new_n928), .C1(new_n790), .C2(new_n713), .ZN(new_n929));
  INV_X1    g0729(.A(G137), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n717), .A2(new_n930), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n714), .A2(G150), .B1(new_n724), .B2(G50), .ZN(new_n932));
  AOI22_X1  g0732(.A1(G143), .A2(new_n727), .B1(new_n706), .B2(G159), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n256), .B1(new_n733), .B2(new_n392), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n729), .A2(new_n214), .ZN(new_n935));
  INV_X1    g0735(.A(new_n700), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n934), .B(new_n935), .C1(G77), .C2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n932), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n929), .B1(new_n931), .B2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT47), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n773), .B1(new_n940), .B2(new_n698), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n210), .A2(new_n318), .ZN(new_n942));
  OAI221_X1 g0742(.A(new_n759), .B1(new_n210), .B2(new_n364), .C1(new_n240), .C2(new_n942), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n941), .B(new_n943), .C1(new_n753), .C2(new_n886), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n919), .A2(new_n944), .ZN(G387));
  OR2_X1    g0745(.A1(new_n690), .A2(new_n915), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n690), .A2(new_n915), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n946), .A2(new_n647), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n915), .A2(new_n918), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n714), .A2(G317), .B1(new_n706), .B2(G311), .ZN(new_n950));
  XOR2_X1   g0750(.A(KEYINPUT115), .B(G322), .Z(new_n951));
  OAI221_X1 g0751(.A(new_n950), .B1(new_n790), .B2(new_n723), .C1(new_n745), .C2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT48), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n953), .B1(new_n701), .B2(new_n729), .C1(new_n472), .C2(new_n733), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT49), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n739), .A2(G326), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n256), .B1(new_n936), .B2(G116), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n745), .A2(new_n778), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n364), .A2(new_n729), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n734), .A2(G77), .ZN(new_n962));
  INV_X1    g0762(.A(G150), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n961), .B(new_n962), .C1(new_n963), .C2(new_n717), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n964), .A2(new_n318), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n714), .A2(G50), .B1(G68), .B2(new_n724), .ZN(new_n966));
  INV_X1    g0766(.A(new_n922), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n706), .A2(new_n329), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n965), .A2(new_n966), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n958), .B1(new_n959), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n773), .B1(new_n970), .B2(new_n698), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n646), .A2(G107), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n367), .A2(G50), .ZN(new_n973));
  AOI21_X1  g0773(.A(G45), .B1(new_n973), .B2(KEYINPUT50), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n974), .B1(KEYINPUT50), .B2(new_n973), .C1(new_n214), .C2(new_n314), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n648), .B1(new_n975), .B2(new_n318), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n237), .A2(new_n256), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n976), .B1(new_n977), .B2(G45), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n759), .B(new_n972), .C1(new_n978), .C2(new_n646), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n971), .B(new_n979), .C1(new_n638), .C2(new_n753), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n949), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n948), .A2(new_n981), .ZN(G393));
  NAND2_X1  g0782(.A1(new_n881), .A2(new_n752), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n759), .B1(new_n261), .B2(new_n210), .C1(new_n249), .C2(new_n942), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n714), .A2(G311), .B1(new_n727), .B2(G317), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT52), .Z(new_n986));
  OAI22_X1  g0786(.A1(new_n729), .A2(new_n248), .B1(new_n733), .B2(new_n701), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n742), .B(new_n987), .C1(new_n706), .C2(G303), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n318), .B1(new_n951), .B2(new_n717), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(new_n724), .B2(G294), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n745), .A2(new_n963), .B1(new_n713), .B2(new_n778), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT51), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n992), .A2(new_n993), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n723), .A2(new_n367), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n730), .A2(G77), .B1(new_n734), .B2(G68), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n777), .B2(new_n717), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n996), .B(new_n998), .C1(G50), .C2(new_n706), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n994), .A2(new_n256), .A3(new_n995), .A4(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n991), .B1(new_n784), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n773), .B1(new_n1001), .B2(new_n698), .ZN(new_n1002));
  AND3_X1   g0802(.A1(new_n983), .A2(new_n984), .A3(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n907), .A2(new_n908), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1003), .B1(new_n1004), .B2(new_n918), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n916), .A2(new_n647), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1004), .B1(new_n690), .B2(new_n915), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(G390));
  NAND2_X1  g0808(.A1(new_n770), .A2(G330), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n829), .B(new_n1010), .C1(new_n670), .C2(new_n677), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n685), .A2(new_n640), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1012), .A2(new_n768), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1013), .A2(new_n769), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1010), .A2(new_n824), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n829), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1011), .A2(new_n1014), .A3(new_n1017), .ZN(new_n1018));
  AND3_X1   g0818(.A1(new_n1010), .A2(new_n824), .A3(new_n829), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1010), .B1(new_n670), .B2(new_n677), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1019), .B1(new_n1020), .B2(new_n1016), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n851), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1018), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(G330), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n848), .A2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n866), .A2(new_n1025), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n855), .A2(new_n857), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n851), .A2(new_n829), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n859), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n829), .B1(new_n1013), .B2(new_n769), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1032), .A2(new_n859), .A3(new_n823), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1019), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n855), .A2(new_n857), .B1(new_n1029), .B2(new_n859), .ZN(new_n1035));
  AND3_X1   g0835(.A1(new_n1032), .A2(new_n859), .A3(new_n823), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n1035), .A2(new_n1036), .A3(new_n1011), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1027), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1011), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1031), .A2(new_n1033), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n1035), .A2(new_n1036), .B1(new_n1016), .B2(new_n1015), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1038), .A2(new_n647), .A3(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n795), .A2(new_n329), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n318), .B1(new_n730), .B2(G159), .ZN(new_n1046));
  INV_X1    g0846(.A(G128), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1046), .B1(new_n202), .B2(new_n700), .C1(new_n745), .C2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G137), .B2(new_n706), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n733), .A2(new_n963), .ZN(new_n1050));
  XOR2_X1   g0850(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1051));
  XNOR2_X1  g0851(.A(new_n1050), .B(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n719), .A2(G125), .ZN(new_n1053));
  XOR2_X1   g0853(.A(KEYINPUT54), .B(G143), .Z(new_n1054));
  AOI22_X1  g0854(.A1(new_n714), .A2(G132), .B1(new_n724), .B2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1049), .A2(new_n1052), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT117), .Z(new_n1057));
  OAI22_X1  g0857(.A1(new_n713), .A2(new_n248), .B1(new_n314), .B2(new_n729), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n318), .B1(new_n220), .B2(new_n733), .C1(new_n745), .C2(new_n701), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n746), .A2(new_n355), .B1(new_n261), .B2(new_n723), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1058), .B(new_n1059), .C1(KEYINPUT118), .C2(new_n1060), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n718), .A2(new_n472), .B1(new_n214), .B2(new_n700), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT119), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1061), .B(new_n1063), .C1(KEYINPUT118), .C2(new_n1060), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n1057), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n698), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n695), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1045), .B(new_n1067), .C1(new_n1028), .C2(new_n750), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1068), .B1(new_n1069), .B2(new_n918), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1044), .A2(new_n1070), .ZN(G378));
  XNOR2_X1  g0871(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n351), .B(KEYINPUT55), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n337), .A2(new_n628), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1073), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1079), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(new_n1072), .A3(new_n1077), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n864), .A2(new_n1084), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1024), .B(new_n831), .C1(new_n845), .C2(new_n846), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n853), .A2(new_n1083), .A3(new_n861), .A4(new_n863), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1085), .A2(new_n1087), .B1(G330), .B2(new_n847), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n918), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(G41), .B1(new_n936), .B2(G159), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n714), .A2(G128), .B1(G150), .B2(new_n730), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G125), .A2(new_n727), .B1(new_n706), .B2(G132), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n734), .A2(new_n1054), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n724), .A2(G137), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT59), .Z(new_n1097));
  AOI21_X1  g0897(.A(G33), .B1(new_n739), .B2(G124), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(G50), .B1(new_n255), .B2(new_n264), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n727), .A2(G116), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n935), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n700), .A2(new_n392), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1101), .A2(new_n1102), .A3(new_n962), .A4(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G97), .B2(new_n706), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n713), .A2(new_n355), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n718), .A2(new_n701), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n723), .A2(new_n364), .ZN(new_n1108));
  NOR4_X1   g0908(.A1(new_n1106), .A2(new_n256), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1105), .A2(new_n264), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT58), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1100), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1091), .A2(new_n1099), .B1(new_n1113), .B2(KEYINPUT120), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1114), .B1(KEYINPUT120), .B2(new_n1113), .C1(new_n1111), .C2(new_n1110), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n773), .B1(new_n1115), .B2(new_n698), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1116), .B1(G50), .B2(new_n795), .C1(new_n1083), .C2(new_n751), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT122), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1090), .A2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n865), .B(new_n621), .C1(new_n1024), .C2(new_n848), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1041), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1088), .A2(new_n1089), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT57), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n692), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OAI221_X1 g0925(.A(KEYINPUT57), .B1(new_n1122), .B2(new_n1121), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1120), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(G375));
  OR2_X1    g0928(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1129), .A2(new_n1121), .A3(new_n1018), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1130), .A2(new_n900), .A3(new_n1041), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n829), .A2(new_n751), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n795), .A2(G68), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n719), .A2(G303), .B1(new_n724), .B2(G107), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n256), .B1(new_n734), .B2(G97), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1134), .B(new_n1135), .C1(new_n314), .C2(new_n700), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G116), .B2(new_n706), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n961), .B1(new_n713), .B2(new_n701), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT123), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1137), .B(new_n1139), .C1(new_n472), .C2(new_n745), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1103), .B(new_n256), .C1(new_n778), .C2(new_n733), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n727), .A2(G132), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(new_n706), .C2(new_n1054), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n713), .A2(new_n930), .B1(new_n718), .B2(new_n1047), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(G150), .B2(new_n724), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1143), .B(new_n1145), .C1(new_n202), .C2(new_n729), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1066), .B1(new_n1140), .B2(new_n1146), .ZN(new_n1147));
  NOR4_X1   g0947(.A1(new_n1132), .A2(new_n773), .A3(new_n1133), .A4(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n1023), .B2(new_n918), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1131), .A2(new_n1149), .ZN(G381));
  NAND4_X1  g0950(.A1(new_n1090), .A2(new_n1119), .A3(new_n1070), .A4(new_n1044), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(G393), .A2(G396), .ZN(new_n1154));
  INV_X1    g0954(.A(G390), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1154), .A2(new_n1155), .A3(new_n919), .A4(new_n944), .ZN(new_n1156));
  OR4_X1    g0956(.A1(G384), .A2(new_n1153), .A3(new_n1156), .A4(G381), .ZN(G407));
  OAI211_X1 g0957(.A(G407), .B(G213), .C1(G343), .C2(new_n1153), .ZN(G409));
  NAND3_X1  g0958(.A1(new_n919), .A2(new_n944), .A3(G390), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(G390), .B1(new_n919), .B2(new_n944), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n764), .B1(new_n948), .B2(new_n981), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n1160), .A2(new_n1161), .B1(new_n1154), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1161), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1154), .A2(new_n1162), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1164), .A2(new_n1165), .A3(new_n1159), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(G378), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1169), .A2(new_n647), .A3(new_n1126), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1120), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1168), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1123), .A2(new_n901), .ZN(new_n1173));
  INV_X1    g0973(.A(G213), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n1151), .A2(new_n1173), .B1(new_n1174), .B2(G343), .ZN(new_n1175));
  OAI21_X1  g0975(.A(KEYINPUT127), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1174), .A2(G343), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1086), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n693), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(G378), .A2(new_n1182), .A3(new_n1118), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n1123), .A2(new_n901), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1177), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT127), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(new_n1168), .C2(new_n1127), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT60), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1130), .A2(new_n1188), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1129), .A2(KEYINPUT60), .A3(new_n1121), .A4(new_n1018), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1189), .A2(new_n647), .A3(new_n1041), .A4(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n1149), .ZN(new_n1192));
  INV_X1    g0992(.A(G384), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1191), .A2(G384), .A3(new_n1149), .ZN(new_n1195));
  OR3_X1    g0995(.A1(new_n1174), .A2(KEYINPUT125), .A3(G343), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1177), .A2(G2897), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1194), .A2(new_n1195), .A3(new_n1198), .A4(new_n1196), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1176), .A2(new_n1187), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1172), .A2(new_n1204), .A3(new_n1175), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT62), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT61), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1203), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1176), .A2(new_n1187), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1204), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1206), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1167), .B1(new_n1209), .B2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1163), .A2(new_n1166), .A3(new_n1208), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT126), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1200), .A2(new_n1215), .A3(new_n1201), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1215), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1185), .B1(new_n1168), .B2(new_n1127), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1214), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(KEYINPUT124), .B1(new_n1205), .B2(KEYINPUT63), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1210), .A2(KEYINPUT63), .A3(new_n1211), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT124), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT63), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(new_n1219), .C2(new_n1204), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .A4(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1213), .A2(new_n1226), .ZN(G405));
  OAI211_X1 g1027(.A(new_n1153), .B(new_n1204), .C1(new_n1168), .C2(new_n1127), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1211), .B1(new_n1172), .B2(new_n1152), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(new_n1167), .Z(G402));
endmodule


