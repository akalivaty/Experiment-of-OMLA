//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  XNOR2_X1  g001(.A(G143), .B(G146), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT68), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  OAI211_X1 g005(.A(new_n190), .B(KEYINPUT1), .C1(new_n191), .C2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G128), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n190), .B1(new_n195), .B2(KEYINPUT1), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n189), .B1(new_n193), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n191), .A2(G146), .ZN(new_n199));
  AND4_X1   g013(.A1(new_n198), .A2(new_n195), .A3(new_n199), .A4(G128), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT11), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G137), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT11), .A3(G134), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n204), .A2(G137), .ZN(new_n208));
  AND3_X1   g022(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT66), .B(G131), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n206), .A2(G134), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n208), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n209), .A2(new_n211), .B1(G131), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n202), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT72), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n209), .A2(new_n211), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n218), .A2(KEYINPUT67), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n205), .A2(new_n207), .A3(new_n220), .A4(new_n208), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G131), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n217), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n195), .A2(new_n199), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT71), .ZN(new_n226));
  OR2_X1    g040(.A1(KEYINPUT0), .A2(G128), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n225), .B(new_n226), .C1(new_n229), .C2(new_n188), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n191), .A2(G146), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n194), .A2(G143), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n228), .B(new_n227), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n226), .B1(new_n234), .B2(new_n225), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n223), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G119), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G116), .ZN(new_n238));
  INV_X1    g052(.A(G116), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G119), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT2), .B(G113), .ZN(new_n242));
  OR2_X1    g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n242), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT72), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n202), .A2(new_n247), .A3(new_n214), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n216), .A2(new_n236), .A3(new_n246), .A4(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT1), .B1(new_n191), .B2(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT68), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(G128), .A3(new_n192), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n200), .B1(new_n253), .B2(new_n189), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n213), .A2(G131), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n255), .B1(new_n218), .B2(new_n210), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n250), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n202), .A2(KEYINPUT69), .A3(new_n214), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n225), .B(new_n259), .C1(new_n229), .C2(new_n188), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n259), .B1(new_n234), .B2(new_n225), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n257), .A2(new_n258), .B1(new_n223), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n249), .B1(new_n264), .B2(new_n246), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT28), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n236), .A2(new_n246), .A3(new_n215), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT28), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G237), .ZN(new_n271));
  INV_X1    g085(.A(G953), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(G210), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n273), .B(KEYINPUT27), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G101), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n274), .B(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT70), .ZN(new_n278));
  XOR2_X1   g092(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n279));
  OAI21_X1  g093(.A(new_n278), .B1(new_n264), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n262), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n223), .A2(new_n281), .A3(new_n260), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n254), .A2(new_n250), .A3(new_n256), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT69), .B1(new_n202), .B2(new_n214), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n279), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(KEYINPUT70), .A3(new_n286), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n216), .A2(new_n236), .A3(KEYINPUT30), .A4(new_n248), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n280), .A2(new_n287), .A3(new_n245), .A4(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n249), .A2(new_n276), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n290), .B1(new_n289), .B2(new_n291), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT31), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT31), .B1(new_n289), .B2(new_n291), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n277), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(G472), .A2(G902), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n187), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n289), .A2(new_n291), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT73), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n295), .B1(new_n304), .B2(KEYINPUT31), .ZN(new_n305));
  OAI211_X1 g119(.A(KEYINPUT32), .B(new_n298), .C1(new_n305), .C2(new_n277), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n270), .A2(KEYINPUT74), .A3(new_n276), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n266), .A2(new_n269), .A3(new_n276), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT29), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n289), .A2(new_n249), .ZN(new_n311));
  INV_X1    g125(.A(new_n276), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n307), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G902), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n216), .A2(new_n236), .A3(new_n248), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n245), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n249), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n318), .A2(KEYINPUT75), .A3(KEYINPUT28), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT75), .B1(new_n318), .B2(KEYINPUT28), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n269), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n276), .A2(KEYINPUT29), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n315), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(G472), .B1(new_n314), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n300), .A2(new_n306), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G128), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(KEYINPUT23), .A3(G119), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n237), .A2(G128), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n237), .A2(G128), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n328), .B(new_n329), .C1(new_n330), .C2(KEYINPUT23), .ZN(new_n331));
  XOR2_X1   g145(.A(KEYINPUT24), .B(G110), .Z(new_n332));
  XNOR2_X1  g146(.A(G119), .B(G128), .ZN(new_n333));
  OAI22_X1  g147(.A1(new_n331), .A2(G110), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G125), .ZN(new_n336));
  INV_X1    g150(.A(G125), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G140), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n338), .A3(KEYINPUT16), .ZN(new_n339));
  OR3_X1    g153(.A1(new_n337), .A2(KEYINPUT16), .A3(G140), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n340), .A3(G146), .ZN(new_n341));
  XNOR2_X1  g155(.A(G125), .B(G140), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n194), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n334), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n331), .A2(G110), .B1(new_n332), .B2(new_n333), .ZN(new_n345));
  INV_X1    g159(.A(new_n341), .ZN(new_n346));
  AOI21_X1  g160(.A(G146), .B1(new_n339), .B2(new_n340), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n345), .B(KEYINPUT76), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n339), .A2(new_n340), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n194), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n341), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT76), .B1(new_n352), .B2(new_n345), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n344), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT22), .B(G137), .ZN(new_n355));
  INV_X1    g169(.A(G221), .ZN(new_n356));
  INV_X1    g170(.A(G234), .ZN(new_n357));
  NOR3_X1   g171(.A1(new_n356), .A2(new_n357), .A3(G953), .ZN(new_n358));
  XOR2_X1   g172(.A(new_n355), .B(new_n358), .Z(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n354), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n344), .B(new_n359), .C1(new_n349), .C2(new_n353), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n315), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT25), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n361), .A2(KEYINPUT25), .A3(new_n315), .A4(new_n362), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(KEYINPUT77), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G217), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n368), .B1(G234), .B2(new_n315), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT77), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n363), .A2(new_n370), .A3(new_n364), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n367), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n367), .A2(KEYINPUT78), .A3(new_n369), .A4(new_n371), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n369), .A2(G902), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n361), .A2(new_n362), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n374), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n326), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(G475), .A2(G902), .ZN(new_n380));
  OR2_X1    g194(.A1(new_n342), .A2(new_n194), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n343), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT87), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT87), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n381), .A2(new_n384), .A3(new_n343), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n271), .A2(new_n272), .A3(G214), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(G143), .ZN(new_n387));
  NAND2_X1  g201(.A1(KEYINPUT18), .A2(G131), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n386), .B(new_n191), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(KEYINPUT18), .A3(G131), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n383), .A2(new_n385), .A3(new_n389), .A4(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(G113), .B(G122), .ZN(new_n393));
  INV_X1    g207(.A(G104), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n393), .B(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n390), .A2(new_n210), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n387), .A2(new_n211), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT17), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n351), .B(new_n341), .C1(new_n396), .C2(new_n398), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n392), .B(new_n395), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n342), .B(KEYINPUT19), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT88), .B1(new_n404), .B2(G146), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n346), .B1(new_n396), .B2(new_n397), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT88), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(new_n407), .A3(new_n194), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n395), .B1(new_n409), .B2(new_n392), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n380), .B1(new_n402), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT20), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT20), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n413), .B(new_n380), .C1(new_n402), .C2(new_n410), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n392), .B1(new_n399), .B2(new_n400), .ZN(new_n416));
  INV_X1    g230(.A(new_n395), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n315), .B1(new_n418), .B2(new_n402), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G475), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n272), .A2(G952), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n357), .B2(new_n271), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  XOR2_X1   g238(.A(KEYINPUT21), .B(G898), .Z(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(KEYINPUT96), .ZN(new_n426));
  AOI211_X1 g240(.A(new_n315), .B(new_n272), .C1(G234), .C2(G237), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n424), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n421), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT9), .B(G234), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n430), .A2(new_n368), .A3(G953), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT89), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n239), .B2(G122), .ZN(new_n433));
  INV_X1    g247(.A(G122), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(KEYINPUT89), .A3(G116), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n239), .A2(G122), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n436), .B1(KEYINPUT14), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT14), .B1(new_n434), .B2(G116), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT92), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT92), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n437), .A2(new_n441), .A3(KEYINPUT14), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G107), .B1(new_n438), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G107), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n433), .A2(new_n435), .B1(new_n239), .B2(G122), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n191), .A2(G128), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n327), .A2(G143), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G134), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n447), .A2(new_n448), .A3(new_n204), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n445), .A2(new_n446), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n444), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT93), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT93), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n444), .A2(new_n452), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n327), .A2(G143), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(KEYINPUT13), .B2(new_n448), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT90), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT13), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT90), .B1(new_n447), .B2(new_n462), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n461), .B(G134), .C1(new_n459), .C2(new_n463), .ZN(new_n464));
  XOR2_X1   g278(.A(new_n451), .B(KEYINPUT91), .Z(new_n465));
  AND2_X1   g279(.A1(new_n446), .A2(new_n445), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n446), .A2(new_n445), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n464), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n431), .B1(new_n457), .B2(new_n468), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n444), .A2(new_n452), .A3(new_n455), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n455), .B1(new_n444), .B2(new_n452), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n468), .B(new_n431), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n315), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT94), .ZN(new_n475));
  INV_X1    g289(.A(G478), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(KEYINPUT15), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n478));
  INV_X1    g292(.A(new_n431), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(G902), .B1(new_n480), .B2(new_n472), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT94), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n475), .A2(new_n477), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n481), .B1(KEYINPUT15), .B2(new_n476), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n484), .A2(KEYINPUT95), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT95), .B1(new_n484), .B2(new_n485), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n429), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  XOR2_X1   g302(.A(KEYINPUT80), .B(G469), .Z(new_n489));
  INV_X1    g303(.A(KEYINPUT82), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT3), .B1(new_n394), .B2(G107), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT3), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n445), .A3(G104), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n394), .A2(G107), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G101), .ZN(new_n496));
  INV_X1    g310(.A(G101), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n491), .A2(new_n493), .A3(new_n497), .A4(new_n494), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n495), .A2(new_n500), .A3(G101), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n499), .B(new_n501), .C1(new_n231), .C2(new_n235), .ZN(new_n502));
  INV_X1    g316(.A(new_n223), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT79), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(new_n445), .A3(G104), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT79), .B1(new_n394), .B2(G107), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n445), .A2(G104), .ZN(new_n507));
  OAI211_X1 g321(.A(G101), .B(new_n505), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n508), .A2(new_n498), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n202), .A2(KEYINPUT10), .A3(new_n509), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n251), .A2(G128), .B1(new_n195), .B2(new_n199), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n498), .B(new_n508), .C1(new_n200), .C2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT10), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n502), .A2(new_n503), .A3(new_n510), .A4(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(G110), .B(G140), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n272), .A2(G227), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n512), .B1(new_n202), .B2(new_n509), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n521), .A2(KEYINPUT12), .A3(new_n223), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT12), .B1(new_n521), .B2(new_n223), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT81), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n520), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT81), .B1(new_n522), .B2(new_n523), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n490), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n521), .A2(new_n223), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT12), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n521), .A2(KEYINPUT12), .A3(new_n223), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n525), .A3(new_n532), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n515), .A2(new_n519), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n527), .A2(new_n533), .A3(new_n534), .A4(new_n490), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n502), .A2(new_n514), .A3(new_n510), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n223), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n515), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n518), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n315), .B(new_n489), .C1(new_n528), .C2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n515), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n518), .B1(new_n524), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n537), .A2(new_n515), .A3(new_n519), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n315), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G469), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n430), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n356), .B1(new_n549), .B2(new_n315), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(G110), .B(G122), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n238), .A2(new_n240), .A3(KEYINPUT5), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n555), .B(G113), .C1(KEYINPUT5), .C2(new_n238), .ZN(new_n556));
  AND4_X1   g370(.A1(new_n243), .A2(new_n556), .A3(new_n498), .A4(new_n508), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n556), .A2(new_n243), .B1(new_n498), .B2(new_n508), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n499), .A2(new_n245), .A3(new_n501), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n509), .A2(new_n243), .A3(new_n556), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(new_n553), .A3(new_n561), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT84), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n225), .B(G125), .C1(new_n229), .C2(new_n188), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(new_n202), .B2(new_n337), .ZN(new_n567));
  INV_X1    g381(.A(G224), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT7), .B1(new_n568), .B2(G953), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n564), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n565), .B1(new_n254), .B2(G125), .ZN(new_n571));
  INV_X1    g385(.A(new_n569), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(KEYINPUT84), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n565), .B(new_n569), .C1(new_n254), .C2(G125), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT83), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n567), .A2(KEYINPUT83), .A3(new_n569), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n563), .A2(new_n574), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n560), .A2(new_n561), .ZN(new_n580));
  INV_X1    g394(.A(new_n553), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(KEYINPUT6), .A3(new_n562), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT6), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n580), .A2(new_n584), .A3(new_n581), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n568), .A2(G953), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n567), .B(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n583), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(G210), .B1(G237), .B2(G902), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n579), .A2(new_n588), .A3(new_n315), .A4(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n589), .B(KEYINPUT86), .Z(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n579), .A2(new_n588), .A3(new_n315), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n593), .B1(new_n594), .B2(KEYINPUT85), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT85), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n579), .A2(new_n588), .A3(new_n596), .A4(new_n315), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n591), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(G214), .B1(G237), .B2(G902), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NOR4_X1   g414(.A1(new_n488), .A2(new_n552), .A3(new_n598), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n379), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  OAI21_X1  g417(.A(G472), .B1(new_n297), .B2(G902), .ZN(new_n604));
  INV_X1    g418(.A(new_n277), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT31), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n302), .B2(new_n303), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n605), .B1(new_n607), .B2(new_n295), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n298), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n610), .A2(new_n378), .A3(new_n552), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n475), .A2(new_n476), .A3(new_n483), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n476), .A2(G902), .ZN(new_n613));
  NOR2_X1   g427(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT97), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI211_X1 g431(.A(new_n614), .B(new_n617), .C1(new_n480), .C2(new_n472), .ZN(new_n618));
  AND4_X1   g432(.A1(new_n615), .A2(new_n480), .A3(new_n616), .A4(new_n472), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n613), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n612), .A2(new_n620), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n621), .A2(new_n421), .ZN(new_n622));
  INV_X1    g436(.A(new_n589), .ZN(new_n623));
  INV_X1    g437(.A(new_n588), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n570), .A2(new_n573), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n577), .A2(new_n578), .A3(new_n562), .A4(new_n559), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n315), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n623), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n600), .B1(new_n628), .B2(new_n590), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n428), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n611), .A2(new_n622), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(new_n394), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  NOR2_X1   g449(.A1(new_n486), .A2(new_n487), .ZN(new_n636));
  INV_X1    g450(.A(new_n421), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n611), .A2(new_n636), .A3(new_n637), .A4(new_n631), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  AND2_X1   g454(.A1(new_n604), .A2(new_n609), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n360), .A2(KEYINPUT36), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT99), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(new_n354), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n376), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n374), .A2(new_n375), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n601), .A2(new_n641), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT37), .B(G110), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G12));
  INV_X1    g463(.A(G900), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n424), .B1(new_n427), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n421), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n636), .A2(new_n629), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n550), .B1(new_n541), .B2(new_n547), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n646), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n325), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G128), .ZN(G30));
  NAND2_X1  g472(.A1(new_n636), .A2(new_n421), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n659), .A2(new_n600), .A3(new_n646), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n594), .A2(KEYINPUT85), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n597), .A3(new_n592), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n590), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT38), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n651), .B(KEYINPUT39), .Z(new_n666));
  NAND2_X1  g480(.A1(new_n654), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n665), .B1(KEYINPUT40), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n304), .B1(new_n312), .B2(new_n318), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n669), .B2(G902), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n300), .A2(new_n670), .A3(new_n306), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n668), .B(new_n671), .C1(KEYINPUT40), .C2(new_n667), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G143), .ZN(G45));
  INV_X1    g487(.A(new_n651), .ZN(new_n674));
  AND4_X1   g488(.A1(new_n421), .A2(new_n621), .A3(new_n629), .A4(new_n674), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n675), .A2(new_n654), .A3(new_n646), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n325), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT100), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n325), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G146), .ZN(G48));
  INV_X1    g496(.A(new_n631), .ZN(new_n683));
  INV_X1    g497(.A(new_n622), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n315), .B1(new_n528), .B2(new_n540), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G469), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n551), .A3(new_n541), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n683), .A2(new_n684), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n379), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  NOR2_X1   g505(.A1(new_n687), .A2(new_n630), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n326), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n487), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n484), .A2(KEYINPUT95), .A3(new_n485), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n695), .A2(new_n696), .A3(new_n637), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n697), .A2(new_n378), .A3(new_n428), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  INV_X1    g514(.A(new_n646), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n488), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n694), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT101), .B(G119), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G21));
  NOR3_X1   g519(.A1(new_n659), .A2(new_n683), .A3(new_n687), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n608), .A2(new_n315), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n321), .A2(new_n312), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n708), .B1(new_n607), .B2(new_n295), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n298), .B(KEYINPUT102), .Z(new_n710));
  AOI22_X1  g524(.A1(new_n707), .A2(G472), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n378), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n706), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G122), .ZN(G24));
  INV_X1    g528(.A(new_n621), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n715), .A2(new_n637), .A3(new_n651), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n709), .A2(new_n710), .ZN(new_n717));
  AND4_X1   g531(.A1(new_n604), .A2(new_n716), .A3(new_n646), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n692), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n306), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n608), .A2(KEYINPUT105), .A3(KEYINPUT32), .A4(new_n298), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n722), .A2(new_n300), .A3(new_n324), .A4(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT104), .B1(new_n663), .B2(new_n600), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n598), .A2(new_n726), .A3(new_n599), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n531), .A2(new_n532), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n519), .B1(new_n728), .B2(new_n515), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n544), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n537), .A2(KEYINPUT103), .A3(new_n515), .A4(new_n519), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n729), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(G469), .B1(new_n733), .B2(G902), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n550), .B1(new_n541), .B2(new_n734), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n725), .A2(new_n727), .A3(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n716), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n724), .A2(new_n712), .A3(new_n736), .A4(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n325), .A2(new_n736), .A3(new_n712), .A4(new_n716), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n738), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g557(.A(KEYINPUT106), .B(G131), .Z(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(G33));
  AND2_X1   g559(.A1(new_n636), .A2(new_n652), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n325), .A2(new_n736), .A3(new_n712), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G134), .ZN(G36));
  NAND2_X1  g562(.A1(new_n610), .A2(new_n646), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n749), .A2(KEYINPUT109), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n715), .A2(new_n421), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n752), .B1(new_n421), .B2(new_n753), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n751), .A2(new_n754), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n757), .B1(new_n749), .B2(KEYINPUT109), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n750), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(KEYINPUT44), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT110), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n733), .A2(KEYINPUT45), .ZN(new_n762));
  INV_X1    g576(.A(G469), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n763), .B1(new_n545), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(G469), .A2(G902), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(KEYINPUT46), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT107), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n766), .A2(KEYINPUT46), .A3(new_n767), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n770), .B1(new_n771), .B2(new_n541), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(new_n770), .A3(new_n541), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n775), .A2(new_n551), .A3(new_n666), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n725), .A2(new_n727), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n779), .B1(KEYINPUT44), .B2(new_n759), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n761), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G137), .ZN(G39));
  XNOR2_X1  g596(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n774), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n785), .A2(new_n769), .A3(new_n772), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n784), .B1(new_n786), .B2(new_n550), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n775), .A2(new_n551), .A3(new_n783), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n777), .A2(new_n737), .A3(new_n712), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n326), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G140), .ZN(G42));
  NAND4_X1  g606(.A1(new_n712), .A2(new_n551), .A3(new_n599), .A4(new_n751), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n686), .A2(new_n541), .ZN(new_n794));
  AOI211_X1 g608(.A(new_n664), .B(new_n793), .C1(KEYINPUT49), .C2(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n300), .A2(new_n306), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n794), .A2(KEYINPUT49), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT112), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n795), .A2(new_n796), .A3(new_n670), .A4(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n794), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n686), .A2(KEYINPUT114), .A3(new_n541), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n550), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n787), .A2(new_n788), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n423), .B1(new_n755), .B2(new_n756), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n604), .A2(new_n717), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n378), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n777), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n804), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT50), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n664), .A2(new_n599), .A3(new_n687), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n811), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n805), .A2(new_n807), .A3(new_n812), .A4(KEYINPUT50), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n777), .A2(new_n687), .A3(new_n378), .A4(new_n423), .ZN(new_n817));
  INV_X1    g631(.A(new_n671), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n817), .A2(new_n818), .A3(new_n637), .A4(new_n715), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n777), .A2(new_n687), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n805), .A2(new_n820), .A3(new_n711), .A4(new_n646), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n810), .A2(new_n816), .A3(KEYINPUT51), .A4(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n817), .A2(new_n622), .A3(new_n818), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n825), .B(new_n422), .C1(new_n693), .C2(new_n808), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n724), .A2(new_n805), .A3(new_n712), .A4(new_n820), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n827), .A2(KEYINPUT48), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(KEYINPUT48), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n826), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n824), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n822), .B1(new_n804), .B2(new_n809), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT51), .B1(new_n832), .B2(new_n816), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT115), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n810), .A2(new_n816), .A3(new_n823), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n838), .A3(new_n824), .A4(new_n830), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n325), .A2(new_n679), .A3(new_n676), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n679), .B1(new_n325), .B2(new_n676), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n657), .B(new_n719), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n695), .A2(new_n696), .A3(new_n421), .A4(new_n629), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n374), .A2(new_n375), .A3(new_n645), .A4(new_n674), .ZN(new_n845));
  INV_X1    g659(.A(new_n735), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n847), .A2(new_n671), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n848), .B1(new_n847), .B2(new_n671), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT52), .B1(new_n843), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n428), .A2(new_n600), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n421), .B1(new_n485), .B2(new_n484), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n663), .B(new_n853), .C1(new_n622), .C2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n641), .A2(new_n712), .A3(new_n654), .A4(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n713), .A3(new_n647), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n325), .B(new_n712), .C1(new_n601), .C2(new_n688), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n325), .B(new_n692), .C1(new_n698), .C2(new_n702), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n711), .A2(new_n736), .A3(new_n646), .A4(new_n716), .ZN(new_n863));
  INV_X1    g677(.A(new_n655), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n652), .A2(new_n485), .A3(new_n484), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n325), .A2(new_n778), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n747), .A2(new_n863), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n742), .B2(new_n740), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n847), .A2(new_n671), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT113), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n847), .A2(new_n671), .A3(new_n848), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT52), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n718), .A2(new_n692), .B1(new_n656), .B2(new_n325), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n872), .A2(new_n681), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n852), .A2(new_n862), .A3(new_n868), .A4(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n857), .A2(new_n713), .A3(new_n647), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n859), .A2(new_n860), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n747), .A2(new_n863), .A3(new_n866), .ZN(new_n881));
  AND4_X1   g695(.A1(new_n743), .A2(new_n879), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(KEYINPUT53), .A3(new_n852), .A4(new_n875), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n878), .A2(new_n883), .A3(KEYINPUT54), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n840), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(G952), .A2(G953), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n799), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT116), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g706(.A(KEYINPUT116), .B(new_n799), .C1(new_n888), .C2(new_n889), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(G75));
  NOR2_X1   g708(.A1(new_n272), .A2(G952), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n315), .B1(new_n878), .B2(new_n883), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT56), .B1(new_n897), .B2(G210), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n583), .A2(new_n585), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(new_n587), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT55), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n896), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT117), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n897), .A2(new_n904), .ZN(new_n905));
  AOI211_X1 g719(.A(KEYINPUT117), .B(new_n315), .C1(new_n878), .C2(new_n883), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n905), .A2(new_n906), .A3(new_n593), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n903), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n884), .A2(G902), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT117), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n897), .A2(new_n904), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n912), .A2(new_n592), .A3(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n914), .A2(KEYINPUT118), .A3(new_n908), .A4(new_n901), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n902), .B1(new_n910), .B2(new_n915), .ZN(G51));
  NOR2_X1   g730(.A1(new_n905), .A2(new_n906), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n917), .A2(new_n762), .A3(new_n765), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n767), .B(KEYINPUT57), .Z(new_n919));
  NAND3_X1  g733(.A1(new_n886), .A2(new_n887), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n920), .B1(new_n528), .B2(new_n540), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n895), .B1(new_n918), .B2(new_n921), .ZN(G54));
  OR2_X1    g736(.A1(new_n402), .A2(new_n410), .ZN(new_n923));
  AND2_X1   g737(.A1(KEYINPUT58), .A2(G475), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n923), .B1(new_n917), .B2(new_n924), .ZN(new_n925));
  AND4_X1   g739(.A1(new_n923), .A2(new_n912), .A3(new_n913), .A4(new_n924), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n925), .A2(new_n926), .A3(new_n895), .ZN(G60));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT119), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT59), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n886), .A2(new_n887), .A3(new_n930), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n618), .A2(new_n619), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n886), .A2(new_n932), .A3(new_n887), .A4(new_n930), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n934), .A2(new_n896), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT120), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT120), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n934), .A2(new_n938), .A3(new_n896), .A4(new_n935), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n939), .ZN(G63));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT121), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT60), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n884), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n361), .A2(new_n362), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n895), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT61), .B1(new_n946), .B2(KEYINPUT122), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n884), .A2(new_n644), .A3(new_n943), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n946), .B(new_n948), .C1(KEYINPUT122), .C2(KEYINPUT61), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(G66));
  OAI21_X1  g766(.A(G953), .B1(new_n426), .B2(new_n568), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n862), .B2(G953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n899), .B1(G898), .B2(new_n272), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(G69));
  NAND3_X1  g770(.A1(new_n280), .A2(new_n287), .A3(new_n288), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(new_n404), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT123), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n843), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n672), .ZN(new_n961));
  AND2_X1   g775(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n667), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n622), .A2(new_n854), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n379), .A2(new_n964), .A3(new_n778), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n791), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n967), .B1(new_n761), .B2(new_n780), .ZN(new_n968));
  NOR2_X1   g782(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n961), .B1(new_n962), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n963), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n958), .B1(new_n971), .B2(new_n272), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n272), .B1(G227), .B2(G900), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n844), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n776), .A2(new_n712), .A3(new_n724), .A4(new_n976), .ZN(new_n977));
  AND4_X1   g791(.A1(new_n743), .A2(new_n791), .A3(new_n747), .A4(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n781), .A2(new_n272), .A3(new_n960), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(G900), .A2(G953), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n979), .A2(new_n958), .A3(new_n980), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n973), .A2(KEYINPUT125), .A3(new_n975), .A4(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(KEYINPUT125), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n974), .B1(new_n983), .B2(new_n972), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(G72));
  NAND4_X1  g799(.A1(new_n781), .A2(new_n862), .A3(new_n960), .A4(new_n978), .ZN(new_n986));
  XNOR2_X1  g800(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n987));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n311), .A2(new_n276), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n895), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n302), .A2(new_n313), .A3(new_n303), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n994), .A2(new_n989), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n993), .B1(new_n884), .B2(new_n995), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n884), .A2(new_n993), .A3(new_n995), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n992), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n311), .A2(new_n276), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n963), .A2(new_n968), .A3(new_n862), .A4(new_n970), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n999), .B1(new_n1000), .B2(new_n989), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n998), .A2(new_n1001), .ZN(G57));
endmodule


