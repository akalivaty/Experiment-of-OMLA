

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798;

  AND2_X1 U373 ( .A1(n411), .A2(KEYINPUT68), .ZN(n656) );
  XNOR2_X1 U374 ( .A(n529), .B(G101), .ZN(n533) );
  NOR2_X1 U375 ( .A1(n785), .A2(n768), .ZN(n352) );
  XOR2_X2 U376 ( .A(KEYINPUT105), .B(n646), .Z(n647) );
  NAND2_X1 U377 ( .A1(n349), .A2(n659), .ZN(n676) );
  NAND2_X1 U378 ( .A1(n423), .A2(KEYINPUT44), .ZN(n349) );
  NAND2_X1 U379 ( .A1(n350), .A2(n447), .ZN(n662) );
  NAND2_X1 U380 ( .A1(n479), .A2(n477), .ZN(n350) );
  XNOR2_X2 U381 ( .A(n548), .B(n782), .ZN(n761) );
  XNOR2_X2 U382 ( .A(n351), .B(n572), .ZN(n782) );
  XOR2_X1 U383 ( .A(G122), .B(G140), .Z(n519) );
  BUF_X1 U384 ( .A(G119), .Z(n409) );
  XNOR2_X2 U385 ( .A(G116), .B(G119), .ZN(n531) );
  XNOR2_X2 U386 ( .A(n561), .B(n488), .ZN(n547) );
  AND2_X1 U387 ( .A1(n355), .A2(n353), .ZN(n371) );
  AND2_X1 U388 ( .A1(n354), .A2(n441), .ZN(n353) );
  AND2_X1 U389 ( .A1(n382), .A2(n644), .ZN(n381) );
  XNOR2_X1 U390 ( .A(n446), .B(KEYINPUT39), .ZN(n632) );
  AND2_X1 U391 ( .A1(n376), .A2(n379), .ZN(n375) );
  XNOR2_X1 U392 ( .A(n727), .B(KEYINPUT107), .ZN(n648) );
  OR2_X1 U393 ( .A1(n761), .A2(n483), .ZN(n482) );
  OR2_X1 U394 ( .A1(n380), .A2(n604), .ZN(n378) );
  INV_X1 U395 ( .A(KEYINPUT47), .ZN(n367) );
  NOR2_X1 U396 ( .A1(n755), .A2(n515), .ZN(n474) );
  NAND2_X1 U397 ( .A1(n369), .A2(n498), .ZN(n504) );
  NAND2_X1 U398 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U399 ( .A1(n371), .A2(n370), .ZN(n785) );
  NAND2_X1 U400 ( .A1(n372), .A2(n356), .ZN(n355) );
  OR2_X1 U401 ( .A1(n357), .A2(n494), .ZN(n354) );
  XNOR2_X1 U402 ( .A(n358), .B(KEYINPUT46), .ZN(n372) );
  NAND2_X1 U403 ( .A1(n405), .A2(n381), .ZN(n659) );
  XNOR2_X1 U404 ( .A(n490), .B(n609), .ZN(n796) );
  NOR2_X1 U405 ( .A1(n418), .A2(n650), .ZN(n694) );
  NAND2_X1 U406 ( .A1(n366), .A2(n365), .ZN(n629) );
  NAND2_X1 U407 ( .A1(n623), .A2(n363), .ZN(n365) );
  NAND2_X1 U408 ( .A1(n368), .A2(n620), .ZN(n700) );
  XNOR2_X1 U409 ( .A(n602), .B(KEYINPUT99), .ZN(n665) );
  NOR2_X1 U410 ( .A1(n662), .A2(n633), .ZN(n424) );
  AND2_X1 U411 ( .A1(KEYINPUT70), .A2(n661), .ZN(n623) );
  XNOR2_X1 U412 ( .A(n359), .B(KEYINPUT28), .ZN(n612) );
  AND2_X1 U413 ( .A1(n610), .A2(n360), .ZN(n359) );
  NOR2_X1 U414 ( .A1(n374), .A2(n373), .ZN(n606) );
  NOR2_X1 U415 ( .A1(n480), .A2(n393), .ZN(n479) );
  OR2_X1 U416 ( .A1(n648), .A2(n378), .ZN(n377) );
  OR2_X1 U417 ( .A1(n652), .A2(KEYINPUT88), .ZN(n396) );
  INV_X1 U418 ( .A(n648), .ZN(n360) );
  AND2_X1 U419 ( .A1(n438), .A2(n397), .ZN(n428) );
  XNOR2_X1 U420 ( .A(n727), .B(n421), .ZN(n652) );
  NOR2_X1 U421 ( .A1(n482), .A2(n481), .ZN(n480) );
  XNOR2_X1 U422 ( .A(n445), .B(n442), .ZN(n766) );
  INV_X1 U423 ( .A(n605), .ZN(n379) );
  NAND2_X1 U424 ( .A1(n380), .A2(n604), .ZN(n376) );
  XNOR2_X1 U425 ( .A(n545), .B(n544), .ZN(n548) );
  OR2_X1 U426 ( .A1(n436), .A2(n391), .ZN(n433) );
  XNOR2_X1 U427 ( .A(n776), .B(KEYINPUT75), .ZN(n539) );
  XNOR2_X1 U428 ( .A(n538), .B(G107), .ZN(n776) );
  XNOR2_X1 U429 ( .A(n416), .B(KEYINPUT35), .ZN(n383) );
  XNOR2_X1 U430 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U431 ( .A(G104), .B(G110), .ZN(n538) );
  XNOR2_X1 U432 ( .A(KEYINPUT18), .B(KEYINPUT80), .ZN(n417) );
  XNOR2_X2 U433 ( .A(G137), .B(G140), .ZN(n572) );
  INV_X1 U434 ( .A(KEYINPUT64), .ZN(n497) );
  XOR2_X1 U435 ( .A(G146), .B(G125), .Z(n535) );
  NAND2_X1 U436 ( .A1(n761), .A2(G469), .ZN(n487) );
  XNOR2_X2 U437 ( .A(n547), .B(n546), .ZN(n351) );
  XNOR2_X1 U438 ( .A(n495), .B(n351), .ZN(n684) );
  NAND2_X1 U439 ( .A1(n352), .A2(n677), .ZN(n681) );
  NAND2_X1 U440 ( .A1(n352), .A2(KEYINPUT2), .ZN(n683) );
  AND2_X1 U441 ( .A1(n357), .A2(n494), .ZN(n356) );
  XNOR2_X1 U442 ( .A(n631), .B(KEYINPUT72), .ZN(n357) );
  NOR2_X1 U443 ( .A1(n796), .A2(n795), .ZN(n358) );
  NAND2_X1 U444 ( .A1(n361), .A2(n367), .ZN(n366) );
  NAND2_X1 U445 ( .A1(n623), .A2(n362), .ZN(n361) );
  INV_X1 U446 ( .A(n700), .ZN(n362) );
  INV_X1 U447 ( .A(n619), .ZN(n368) );
  NOR2_X1 U448 ( .A1(n619), .A2(n364), .ZN(n363) );
  NAND2_X1 U449 ( .A1(n620), .A2(KEYINPUT47), .ZN(n364) );
  XNOR2_X2 U450 ( .A(n682), .B(n492), .ZN(n369) );
  NAND2_X1 U451 ( .A1(n500), .A2(n369), .ZN(n685) );
  NAND2_X1 U452 ( .A1(n499), .A2(n369), .ZN(n760) );
  NAND2_X1 U453 ( .A1(n493), .A2(n369), .ZN(n491) );
  OR2_X1 U454 ( .A1(n372), .A2(n494), .ZN(n370) );
  AND2_X1 U455 ( .A1(n648), .A2(n604), .ZN(n373) );
  NAND2_X1 U456 ( .A1(n377), .A2(n375), .ZN(n374) );
  INV_X1 U457 ( .A(n712), .ZN(n380) );
  XNOR2_X1 U458 ( .A(n643), .B(n383), .ZN(n382) );
  NAND2_X1 U459 ( .A1(n384), .A2(n452), .ZN(n451) );
  OR2_X2 U460 ( .A1(n651), .A2(n396), .ZN(n384) );
  XNOR2_X2 U461 ( .A(n510), .B(n509), .ZN(n651) );
  BUF_X1 U462 ( .A(n768), .Z(n385) );
  BUF_X1 U463 ( .A(n387), .Z(n386) );
  XNOR2_X1 U464 ( .A(n643), .B(KEYINPUT35), .ZN(n387) );
  BUF_X1 U465 ( .A(n413), .Z(n388) );
  NAND2_X1 U466 ( .A1(n639), .A2(n638), .ZN(n389) );
  NAND2_X1 U467 ( .A1(n639), .A2(n638), .ZN(n511) );
  XNOR2_X1 U468 ( .A(n547), .B(n539), .ZN(n540) );
  XNOR2_X1 U469 ( .A(n539), .B(n394), .ZN(n545) );
  NOR2_X1 U470 ( .A1(n451), .A2(n450), .ZN(n390) );
  NOR2_X1 U471 ( .A1(n451), .A2(n450), .ZN(n686) );
  NOR2_X2 U472 ( .A1(n404), .A2(n752), .ZN(n640) );
  AND2_X2 U473 ( .A1(n757), .A2(n392), .ZN(n434) );
  INV_X1 U474 ( .A(KEYINPUT4), .ZN(n488) );
  AND2_X1 U475 ( .A1(n482), .A2(n481), .ZN(n478) );
  AND2_X1 U476 ( .A1(n455), .A2(n710), .ZN(n441) );
  XNOR2_X1 U477 ( .A(n535), .B(KEYINPUT10), .ZN(n783) );
  INV_X1 U478 ( .A(KEYINPUT65), .ZN(n492) );
  BUF_X1 U479 ( .A(n728), .Z(n418) );
  NAND2_X1 U480 ( .A1(n487), .A2(n486), .ZN(n476) );
  NAND2_X1 U481 ( .A1(G469), .A2(G902), .ZN(n486) );
  NAND2_X1 U482 ( .A1(n549), .A2(n484), .ZN(n483) );
  INV_X1 U483 ( .A(G902), .ZN(n484) );
  INV_X1 U484 ( .A(KEYINPUT106), .ZN(n507) );
  XNOR2_X1 U485 ( .A(G113), .B(G104), .ZN(n518) );
  XOR2_X1 U486 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n521) );
  XNOR2_X1 U487 ( .A(G143), .B(G131), .ZN(n523) );
  XNOR2_X1 U488 ( .A(G101), .B(G146), .ZN(n543) );
  NAND2_X1 U489 ( .A1(G234), .A2(G237), .ZN(n589) );
  OR2_X1 U490 ( .A1(n436), .A2(n395), .ZN(n430) );
  XNOR2_X1 U491 ( .A(n603), .B(KEYINPUT30), .ZN(n604) );
  INV_X1 U492 ( .A(KEYINPUT111), .ZN(n603) );
  INV_X1 U493 ( .A(KEYINPUT6), .ZN(n421) );
  XNOR2_X1 U494 ( .A(G131), .B(G134), .ZN(n546) );
  NOR2_X1 U495 ( .A1(G953), .A2(G237), .ZN(n552) );
  XNOR2_X1 U496 ( .A(G146), .B(KEYINPUT5), .ZN(n550) );
  INV_X1 U497 ( .A(KEYINPUT22), .ZN(n509) );
  NOR2_X1 U498 ( .A1(n407), .A2(n672), .ZN(n508) );
  NAND2_X1 U499 ( .A1(n652), .A2(KEYINPUT88), .ZN(n453) );
  XNOR2_X1 U500 ( .A(n444), .B(n443), .ZN(n442) );
  INV_X1 U501 ( .A(G210), .ZN(n502) );
  NOR2_X1 U502 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U503 ( .A1(n754), .A2(G953), .ZN(n516) );
  XNOR2_X1 U504 ( .A(KEYINPUT96), .B(KEYINPUT20), .ZN(n580) );
  INV_X1 U505 ( .A(KEYINPUT68), .ZN(n416) );
  NOR2_X1 U506 ( .A1(G237), .A2(G902), .ZN(n541) );
  XOR2_X1 U507 ( .A(G902), .B(KEYINPUT15), .Z(n677) );
  OR2_X1 U508 ( .A1(n392), .A2(n677), .ZN(n439) );
  XNOR2_X1 U509 ( .A(n475), .B(n535), .ZN(n536) );
  XNOR2_X1 U510 ( .A(n417), .B(KEYINPUT17), .ZN(n475) );
  INV_X1 U511 ( .A(KEYINPUT38), .ZN(n454) );
  INV_X1 U512 ( .A(G953), .ZN(n770) );
  XNOR2_X1 U513 ( .A(G110), .B(KEYINPUT24), .ZN(n577) );
  XNOR2_X1 U514 ( .A(G128), .B(n409), .ZN(n574) );
  XNOR2_X1 U515 ( .A(G134), .B(G116), .ZN(n558) );
  XOR2_X1 U516 ( .A(G122), .B(G107), .Z(n559) );
  XNOR2_X1 U517 ( .A(n525), .B(n426), .ZN(n569) );
  XNOR2_X1 U518 ( .A(n783), .B(n526), .ZN(n426) );
  XNOR2_X1 U519 ( .A(n543), .B(n542), .ZN(n544) );
  INV_X1 U520 ( .A(KEYINPUT85), .ZN(n512) );
  NAND2_X1 U521 ( .A1(n428), .A2(n429), .ZN(n419) );
  INV_X1 U522 ( .A(KEYINPUT78), .ZN(n607) );
  XNOR2_X1 U523 ( .A(n551), .B(n553), .ZN(n496) );
  XNOR2_X1 U524 ( .A(KEYINPUT16), .B(G122), .ZN(n534) );
  INV_X1 U525 ( .A(G217), .ZN(n503) );
  XNOR2_X1 U526 ( .A(n598), .B(n425), .ZN(n599) );
  XNOR2_X1 U527 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n425) );
  XNOR2_X1 U528 ( .A(KEYINPUT32), .B(KEYINPUT81), .ZN(n654) );
  INV_X1 U529 ( .A(KEYINPUT31), .ZN(n449) );
  AND2_X1 U530 ( .A1(n508), .A2(n453), .ZN(n452) );
  INV_X1 U531 ( .A(n766), .ZN(n465) );
  INV_X1 U532 ( .A(KEYINPUT56), .ZN(n460) );
  NAND2_X1 U533 ( .A1(n756), .A2(n516), .ZN(n515) );
  INV_X1 U534 ( .A(G122), .ZN(n415) );
  AND2_X1 U535 ( .A1(n392), .A2(n677), .ZN(n391) );
  AND2_X1 U536 ( .A1(G210), .A2(n596), .ZN(n392) );
  AND2_X1 U537 ( .A1(n476), .A2(KEYINPUT1), .ZN(n393) );
  INV_X1 U538 ( .A(KEYINPUT1), .ZN(n481) );
  AND2_X1 U539 ( .A1(G227), .A2(n786), .ZN(n394) );
  AND2_X1 U540 ( .A1(n712), .A2(n437), .ZN(n395) );
  NOR2_X1 U541 ( .A1(n391), .A2(n437), .ZN(n397) );
  XOR2_X1 U542 ( .A(KEYINPUT67), .B(KEYINPUT0), .Z(n398) );
  XOR2_X1 U543 ( .A(n759), .B(n758), .Z(n399) );
  XOR2_X1 U544 ( .A(n684), .B(KEYINPUT62), .Z(n400) );
  XOR2_X1 U545 ( .A(n763), .B(n762), .Z(n401) );
  XNOR2_X1 U546 ( .A(n528), .B(n527), .ZN(n402) );
  XOR2_X1 U547 ( .A(KEYINPUT66), .B(KEYINPUT60), .Z(n403) );
  AND2_X1 U548 ( .A1(n651), .A2(KEYINPUT88), .ZN(n450) );
  XNOR2_X2 U549 ( .A(n389), .B(n398), .ZN(n404) );
  XNOR2_X1 U550 ( .A(n511), .B(n398), .ZN(n667) );
  NOR2_X1 U551 ( .A1(n412), .A2(n694), .ZN(n405) );
  NOR2_X1 U552 ( .A1(n412), .A2(n694), .ZN(n657) );
  OR2_X1 U553 ( .A1(n757), .A2(n439), .ZN(n406) );
  OR2_X1 U554 ( .A1(n757), .A2(n439), .ZN(n438) );
  NAND2_X1 U555 ( .A1(n479), .A2(n477), .ZN(n407) );
  AND2_X1 U556 ( .A1(n757), .A2(n392), .ZN(n408) );
  BUF_X1 U557 ( .A(n412), .Z(n410) );
  NAND2_X1 U558 ( .A1(n387), .A2(n414), .ZN(n411) );
  XNOR2_X1 U559 ( .A(n424), .B(KEYINPUT33), .ZN(n752) );
  XNOR2_X1 U560 ( .A(n655), .B(n654), .ZN(n412) );
  INV_X1 U561 ( .A(n767), .ZN(n468) );
  XNOR2_X1 U562 ( .A(n410), .B(n798), .ZN(G21) );
  XNOR2_X2 U563 ( .A(n413), .B(KEYINPUT19), .ZN(n639) );
  NOR2_X1 U564 ( .A1(n616), .A2(n388), .ZN(n617) );
  NAND2_X2 U565 ( .A1(n435), .A2(n419), .ZN(n413) );
  INV_X1 U566 ( .A(KEYINPUT89), .ZN(n414) );
  XNOR2_X1 U567 ( .A(n386), .B(n415), .ZN(G24) );
  XNOR2_X2 U568 ( .A(n601), .B(KEYINPUT69), .ZN(n447) );
  XNOR2_X1 U569 ( .A(n579), .B(KEYINPUT95), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n420), .B(n507), .ZN(n471) );
  OR2_X2 U571 ( .A1(n686), .A2(n673), .ZN(n420) );
  INV_X1 U572 ( .A(n504), .ZN(n464) );
  XNOR2_X2 U573 ( .A(n555), .B(n554), .ZN(n727) );
  XNOR2_X2 U574 ( .A(n422), .B(n540), .ZN(n757) );
  XNOR2_X2 U575 ( .A(n777), .B(n506), .ZN(n422) );
  NAND2_X1 U576 ( .A1(n656), .A2(n657), .ZN(n423) );
  NAND2_X1 U577 ( .A1(n464), .A2(G478), .ZN(n764) );
  XNOR2_X1 U578 ( .A(n427), .B(KEYINPUT109), .ZN(n597) );
  AND2_X1 U579 ( .A1(n615), .A2(n712), .ZN(n427) );
  INV_X1 U580 ( .A(n455), .ZN(n711) );
  NOR2_X1 U581 ( .A1(n434), .A2(n433), .ZN(n432) );
  NOR2_X1 U582 ( .A1(n408), .A2(n391), .ZN(n440) );
  INV_X1 U583 ( .A(n408), .ZN(n429) );
  NAND2_X1 U584 ( .A1(n431), .A2(n430), .ZN(n435) );
  NAND2_X1 U585 ( .A1(n432), .A2(n406), .ZN(n431) );
  NAND2_X1 U586 ( .A1(n440), .A2(n406), .ZN(n456) );
  NOR2_X1 U587 ( .A1(n712), .A2(n437), .ZN(n436) );
  INV_X1 U588 ( .A(KEYINPUT90), .ZN(n437) );
  NOR2_X2 U589 ( .A1(n766), .A2(G902), .ZN(n585) );
  XNOR2_X1 U590 ( .A(n517), .B(KEYINPUT23), .ZN(n443) );
  NAND2_X1 U591 ( .A1(n576), .A2(G221), .ZN(n444) );
  XNOR2_X1 U592 ( .A(n505), .B(n575), .ZN(n445) );
  NAND2_X1 U593 ( .A1(n632), .A2(n704), .ZN(n490) );
  NAND2_X1 U594 ( .A1(n627), .A2(n713), .ZN(n446) );
  XNOR2_X1 U595 ( .A(n608), .B(n607), .ZN(n627) );
  NAND2_X1 U596 ( .A1(n447), .A2(n611), .ZN(n602) );
  NOR2_X1 U597 ( .A1(n407), .A2(n447), .ZN(n725) );
  NOR2_X1 U598 ( .A1(n448), .A2(n691), .ZN(n669) );
  NAND2_X1 U599 ( .A1(n448), .A2(n704), .ZN(n705) );
  NAND2_X1 U600 ( .A1(n448), .A2(n706), .ZN(n707) );
  XNOR2_X1 U601 ( .A(n663), .B(n449), .ZN(n448) );
  NOR2_X1 U602 ( .A1(n651), .A2(n652), .ZN(n670) );
  XNOR2_X1 U603 ( .A(n456), .B(n454), .ZN(n713) );
  AND2_X1 U604 ( .A1(n641), .A2(n456), .ZN(n628) );
  OR2_X1 U605 ( .A1(n599), .A2(n456), .ZN(n455) );
  XNOR2_X2 U606 ( .A(n457), .B(n534), .ZN(n777) );
  XNOR2_X1 U607 ( .A(n457), .B(n496), .ZN(n495) );
  XNOR2_X2 U608 ( .A(n532), .B(n533), .ZN(n457) );
  NAND2_X1 U609 ( .A1(n768), .A2(n744), .ZN(n513) );
  XNOR2_X1 U610 ( .A(n513), .B(n512), .ZN(n746) );
  XNOR2_X1 U611 ( .A(n458), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U612 ( .A1(n459), .A2(n468), .ZN(n458) );
  XNOR2_X1 U613 ( .A(n685), .B(n400), .ZN(n459) );
  XNOR2_X1 U614 ( .A(n461), .B(n460), .ZN(G51) );
  NAND2_X1 U615 ( .A1(n463), .A2(n468), .ZN(n461) );
  NOR2_X1 U616 ( .A1(n749), .A2(n501), .ZN(n493) );
  XNOR2_X1 U617 ( .A(n462), .B(n403), .ZN(G60) );
  NAND2_X1 U618 ( .A1(n469), .A2(n468), .ZN(n462) );
  XNOR2_X1 U619 ( .A(n760), .B(n399), .ZN(n463) );
  XNOR2_X1 U620 ( .A(n466), .B(n465), .ZN(n472) );
  NOR2_X1 U621 ( .A1(n504), .A2(n503), .ZN(n466) );
  XNOR2_X1 U622 ( .A(n467), .B(n401), .ZN(n470) );
  NOR2_X1 U623 ( .A1(n504), .A2(n549), .ZN(n467) );
  XNOR2_X1 U624 ( .A(n491), .B(n402), .ZN(n469) );
  NOR2_X1 U625 ( .A1(n470), .A2(n767), .ZN(G54) );
  XNOR2_X1 U626 ( .A(n764), .B(n765), .ZN(n473) );
  NAND2_X1 U627 ( .A1(n471), .A2(n674), .ZN(n675) );
  NOR2_X1 U628 ( .A1(n472), .A2(n767), .ZN(G66) );
  NOR2_X1 U629 ( .A1(n473), .A2(n767), .ZN(G63) );
  XNOR2_X1 U630 ( .A(n474), .B(KEYINPUT53), .ZN(G75) );
  INV_X1 U631 ( .A(n476), .ZN(n485) );
  NAND2_X1 U632 ( .A1(n485), .A2(n482), .ZN(n611) );
  NAND2_X1 U633 ( .A1(n478), .A2(n485), .ZN(n477) );
  XNOR2_X2 U634 ( .A(n489), .B(G128), .ZN(n561) );
  XNOR2_X2 U635 ( .A(G143), .B(KEYINPUT82), .ZN(n489) );
  XNOR2_X2 U636 ( .A(n683), .B(KEYINPUT77), .ZN(n749) );
  INV_X1 U637 ( .A(KEYINPUT48), .ZN(n494) );
  NOR2_X2 U638 ( .A1(n667), .A2(n647), .ZN(n510) );
  XNOR2_X1 U639 ( .A(n536), .B(n537), .ZN(n506) );
  XNOR2_X2 U640 ( .A(n497), .B(G953), .ZN(n786) );
  NAND2_X1 U641 ( .A1(n786), .A2(G234), .ZN(n557) );
  INV_X1 U642 ( .A(n749), .ZN(n498) );
  NOR2_X1 U643 ( .A1(n749), .A2(n502), .ZN(n499) );
  NOR2_X1 U644 ( .A1(n749), .A2(n554), .ZN(n500) );
  INV_X1 U645 ( .A(G475), .ZN(n501) );
  XNOR2_X2 U646 ( .A(n514), .B(KEYINPUT45), .ZN(n768) );
  NOR2_X2 U647 ( .A1(n675), .A2(n676), .ZN(n514) );
  XNOR2_X1 U648 ( .A(n748), .B(n747), .ZN(n750) );
  XNOR2_X2 U649 ( .A(G113), .B(KEYINPUT3), .ZN(n529) );
  INV_X1 U650 ( .A(n727), .ZN(n664) );
  NOR2_X1 U651 ( .A1(n786), .A2(G952), .ZN(n767) );
  XOR2_X1 U652 ( .A(n578), .B(n577), .Z(n517) );
  INV_X1 U653 ( .A(KEYINPUT79), .ZN(n542) );
  INV_X1 U654 ( .A(KEYINPUT74), .ZN(n530) );
  INV_X1 U655 ( .A(G469), .ZN(n549) );
  INV_X1 U656 ( .A(G472), .ZN(n554) );
  XNOR2_X1 U657 ( .A(KEYINPUT122), .B(KEYINPUT92), .ZN(n528) );
  XNOR2_X1 U658 ( .A(n519), .B(n518), .ZN(n526) );
  NAND2_X1 U659 ( .A1(G214), .A2(n552), .ZN(n520) );
  XNOR2_X1 U660 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U661 ( .A(n522), .B(KEYINPUT101), .Z(n524) );
  XNOR2_X1 U662 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U663 ( .A(n569), .B(KEYINPUT59), .ZN(n527) );
  NAND2_X1 U664 ( .A1(G224), .A2(n786), .ZN(n537) );
  XOR2_X1 U665 ( .A(KEYINPUT76), .B(n541), .Z(n596) );
  XNOR2_X1 U666 ( .A(n550), .B(G137), .ZN(n551) );
  NAND2_X1 U667 ( .A1(n552), .A2(G210), .ZN(n553) );
  NOR2_X1 U668 ( .A1(n684), .A2(G902), .ZN(n555) );
  INV_X1 U669 ( .A(n652), .ZN(n633) );
  XNOR2_X1 U670 ( .A(KEYINPUT71), .B(KEYINPUT8), .ZN(n556) );
  XNOR2_X1 U671 ( .A(n557), .B(n556), .ZN(n576) );
  NAND2_X1 U672 ( .A1(n576), .A2(G217), .ZN(n565) );
  XNOR2_X1 U673 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U674 ( .A(n560), .B(KEYINPUT7), .Z(n563) );
  XNOR2_X1 U675 ( .A(n561), .B(KEYINPUT9), .ZN(n562) );
  XNOR2_X1 U676 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U677 ( .A(n565), .B(n564), .ZN(n765) );
  NOR2_X1 U678 ( .A1(G902), .A2(n765), .ZN(n566) );
  XOR2_X1 U679 ( .A(G478), .B(n566), .Z(n624) );
  INV_X1 U680 ( .A(n624), .ZN(n621) );
  XOR2_X1 U681 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n568) );
  XNOR2_X1 U682 ( .A(KEYINPUT13), .B(G475), .ZN(n567) );
  XNOR2_X1 U683 ( .A(n568), .B(n567), .ZN(n571) );
  NOR2_X1 U684 ( .A1(G902), .A2(n569), .ZN(n570) );
  XNOR2_X1 U685 ( .A(n571), .B(n570), .ZN(n625) );
  NAND2_X1 U686 ( .A1(n621), .A2(n625), .ZN(n701) );
  INV_X1 U687 ( .A(n701), .ZN(n704) );
  INV_X1 U688 ( .A(n572), .ZN(n573) );
  XNOR2_X1 U689 ( .A(n574), .B(n573), .ZN(n579) );
  INV_X1 U690 ( .A(n783), .ZN(n575) );
  XOR2_X1 U691 ( .A(KEYINPUT94), .B(KEYINPUT84), .Z(n578) );
  XOR2_X1 U692 ( .A(KEYINPUT25), .B(KEYINPUT97), .Z(n583) );
  INV_X1 U693 ( .A(n677), .ZN(n678) );
  NAND2_X1 U694 ( .A1(n678), .A2(G234), .ZN(n581) );
  XNOR2_X1 U695 ( .A(n581), .B(n580), .ZN(n586) );
  NAND2_X1 U696 ( .A1(G217), .A2(n586), .ZN(n582) );
  XNOR2_X1 U697 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X2 U698 ( .A(n585), .B(n584), .ZN(n728) );
  NAND2_X1 U699 ( .A1(n586), .A2(G221), .ZN(n587) );
  XNOR2_X1 U700 ( .A(n587), .B(KEYINPUT21), .ZN(n588) );
  XNOR2_X1 U701 ( .A(KEYINPUT98), .B(n588), .ZN(n600) );
  XNOR2_X1 U702 ( .A(n589), .B(KEYINPUT14), .ZN(n636) );
  NAND2_X1 U703 ( .A1(G952), .A2(n770), .ZN(n634) );
  NOR2_X1 U704 ( .A1(G900), .A2(n786), .ZN(n590) );
  NAND2_X1 U705 ( .A1(G902), .A2(n590), .ZN(n591) );
  NAND2_X1 U706 ( .A1(n634), .A2(n591), .ZN(n592) );
  NAND2_X1 U707 ( .A1(n636), .A2(n592), .ZN(n605) );
  NOR2_X1 U708 ( .A1(n600), .A2(n605), .ZN(n593) );
  XNOR2_X1 U709 ( .A(n593), .B(KEYINPUT73), .ZN(n594) );
  NOR2_X1 U710 ( .A1(n728), .A2(n594), .ZN(n610) );
  NAND2_X1 U711 ( .A1(n704), .A2(n610), .ZN(n595) );
  NOR2_X1 U712 ( .A1(n633), .A2(n595), .ZN(n615) );
  NAND2_X1 U713 ( .A1(n596), .A2(G214), .ZN(n712) );
  NOR2_X1 U714 ( .A1(n407), .A2(n597), .ZN(n598) );
  XOR2_X1 U715 ( .A(KEYINPUT112), .B(KEYINPUT40), .Z(n609) );
  INV_X1 U716 ( .A(n600), .ZN(n729) );
  NAND2_X1 U717 ( .A1(n728), .A2(n729), .ZN(n601) );
  NAND2_X1 U718 ( .A1(n665), .A2(n606), .ZN(n608) );
  NAND2_X1 U719 ( .A1(n612), .A2(n611), .ZN(n619) );
  NOR2_X1 U720 ( .A1(n625), .A2(n624), .ZN(n645) );
  INV_X1 U721 ( .A(n645), .ZN(n716) );
  NAND2_X1 U722 ( .A1(n713), .A2(n712), .ZN(n717) );
  NOR2_X1 U723 ( .A1(n716), .A2(n717), .ZN(n613) );
  XNOR2_X1 U724 ( .A(KEYINPUT41), .B(n613), .ZN(n753) );
  NOR2_X1 U725 ( .A1(n619), .A2(n753), .ZN(n614) );
  XNOR2_X1 U726 ( .A(KEYINPUT42), .B(n614), .ZN(n795) );
  INV_X1 U727 ( .A(n407), .ZN(n671) );
  INV_X1 U728 ( .A(n615), .ZN(n616) );
  XOR2_X1 U729 ( .A(KEYINPUT36), .B(n617), .Z(n618) );
  NOR2_X1 U730 ( .A1(n671), .A2(n618), .ZN(n708) );
  BUF_X1 U731 ( .A(n639), .Z(n620) );
  OR2_X1 U732 ( .A1(n625), .A2(n621), .ZN(n622) );
  XNOR2_X1 U733 ( .A(n622), .B(KEYINPUT104), .ZN(n695) );
  NAND2_X1 U734 ( .A1(n695), .A2(n701), .ZN(n661) );
  NAND2_X1 U735 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U736 ( .A(n626), .B(KEYINPUT108), .Z(n641) );
  NAND2_X1 U737 ( .A1(n628), .A2(n627), .ZN(n699) );
  NAND2_X1 U738 ( .A1(n629), .A2(n699), .ZN(n630) );
  NOR2_X1 U739 ( .A1(n708), .A2(n630), .ZN(n631) );
  INV_X1 U740 ( .A(n695), .ZN(n706) );
  NAND2_X1 U741 ( .A1(n632), .A2(n706), .ZN(n710) );
  XOR2_X1 U742 ( .A(G898), .B(KEYINPUT93), .Z(n772) );
  NOR2_X1 U743 ( .A1(n772), .A2(n770), .ZN(n779) );
  NAND2_X1 U744 ( .A1(G902), .A2(n779), .ZN(n635) );
  AND2_X1 U745 ( .A1(n635), .A2(n634), .ZN(n637) );
  INV_X1 U746 ( .A(n636), .ZN(n741) );
  NOR2_X1 U747 ( .A1(n637), .A2(n741), .ZN(n638) );
  XNOR2_X1 U748 ( .A(n640), .B(KEYINPUT34), .ZN(n642) );
  NAND2_X1 U749 ( .A1(n642), .A2(n641), .ZN(n643) );
  INV_X1 U750 ( .A(KEYINPUT44), .ZN(n644) );
  NAND2_X1 U751 ( .A1(n729), .A2(n645), .ZN(n646) );
  NOR2_X1 U752 ( .A1(n651), .A2(n407), .ZN(n649) );
  NAND2_X1 U753 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U754 ( .A1(n418), .A2(n671), .ZN(n653) );
  NAND2_X1 U755 ( .A1(n670), .A2(n653), .ZN(n655) );
  NAND2_X1 U756 ( .A1(n386), .A2(KEYINPUT44), .ZN(n660) );
  NAND2_X1 U757 ( .A1(n660), .A2(KEYINPUT89), .ZN(n674) );
  INV_X1 U758 ( .A(n661), .ZN(n718) );
  OR2_X1 U759 ( .A1(n664), .A2(n662), .ZN(n734) );
  NOR2_X1 U760 ( .A1(n404), .A2(n734), .ZN(n663) );
  NAND2_X1 U761 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U762 ( .A1(n404), .A2(n666), .ZN(n668) );
  XNOR2_X1 U763 ( .A(KEYINPUT100), .B(n668), .ZN(n691) );
  NOR2_X1 U764 ( .A1(n718), .A2(n669), .ZN(n673) );
  INV_X1 U765 ( .A(n418), .ZN(n672) );
  XNOR2_X1 U766 ( .A(n678), .B(KEYINPUT87), .ZN(n679) );
  NAND2_X1 U767 ( .A1(n679), .A2(KEYINPUT2), .ZN(n680) );
  XOR2_X1 U768 ( .A(n390), .B(G101), .Z(G3) );
  NAND2_X1 U769 ( .A1(n691), .A2(n704), .ZN(n687) );
  XNOR2_X1 U770 ( .A(n687), .B(G104), .ZN(G6) );
  XOR2_X1 U771 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n689) );
  XNOR2_X1 U772 ( .A(G107), .B(KEYINPUT113), .ZN(n688) );
  XNOR2_X1 U773 ( .A(n689), .B(n688), .ZN(n690) );
  XOR2_X1 U774 ( .A(KEYINPUT26), .B(n690), .Z(n693) );
  NAND2_X1 U775 ( .A1(n691), .A2(n706), .ZN(n692) );
  XNOR2_X1 U776 ( .A(n693), .B(n692), .ZN(G9) );
  XOR2_X1 U777 ( .A(G110), .B(n694), .Z(G12) );
  NOR2_X1 U778 ( .A1(n695), .A2(n700), .ZN(n697) );
  XNOR2_X1 U779 ( .A(KEYINPUT115), .B(KEYINPUT29), .ZN(n696) );
  XNOR2_X1 U780 ( .A(n697), .B(n696), .ZN(n698) );
  XOR2_X1 U781 ( .A(G128), .B(n698), .Z(G30) );
  XNOR2_X1 U782 ( .A(G143), .B(n699), .ZN(G45) );
  NOR2_X1 U783 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U784 ( .A(KEYINPUT116), .B(n702), .Z(n703) );
  XNOR2_X1 U785 ( .A(G146), .B(n703), .ZN(G48) );
  XNOR2_X1 U786 ( .A(n705), .B(G113), .ZN(G15) );
  XNOR2_X1 U787 ( .A(n707), .B(G116), .ZN(G18) );
  XNOR2_X1 U788 ( .A(G125), .B(n708), .ZN(n709) );
  XNOR2_X1 U789 ( .A(n709), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U790 ( .A(G134), .B(n710), .ZN(G36) );
  XOR2_X1 U791 ( .A(G140), .B(n711), .Z(G42) );
  NOR2_X1 U792 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U793 ( .A(KEYINPUT117), .B(n714), .Z(n715) );
  NOR2_X1 U794 ( .A1(n716), .A2(n715), .ZN(n720) );
  NOR2_X1 U795 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U796 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U797 ( .A(n721), .B(KEYINPUT118), .ZN(n722) );
  NOR2_X1 U798 ( .A1(n752), .A2(n722), .ZN(n723) );
  XOR2_X1 U799 ( .A(KEYINPUT119), .B(n723), .Z(n738) );
  XNOR2_X1 U800 ( .A(n725), .B(KEYINPUT50), .ZN(n726) );
  NOR2_X1 U801 ( .A1(n727), .A2(n726), .ZN(n732) );
  NOR2_X1 U802 ( .A1(n729), .A2(n418), .ZN(n730) );
  XNOR2_X1 U803 ( .A(n730), .B(KEYINPUT49), .ZN(n731) );
  NAND2_X1 U804 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U805 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U806 ( .A(KEYINPUT51), .B(n735), .ZN(n736) );
  NOR2_X1 U807 ( .A1(n753), .A2(n736), .ZN(n737) );
  NOR2_X1 U808 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U809 ( .A(n739), .B(KEYINPUT52), .ZN(n740) );
  NOR2_X1 U810 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U811 ( .A1(n742), .A2(G952), .ZN(n743) );
  XNOR2_X1 U812 ( .A(n743), .B(KEYINPUT120), .ZN(n756) );
  INV_X1 U813 ( .A(KEYINPUT2), .ZN(n744) );
  NAND2_X1 U814 ( .A1(n744), .A2(n785), .ZN(n745) );
  NAND2_X1 U815 ( .A1(n746), .A2(n745), .ZN(n748) );
  INV_X1 U816 ( .A(KEYINPUT83), .ZN(n747) );
  XNOR2_X1 U817 ( .A(n751), .B(KEYINPUT86), .ZN(n755) );
  NOR2_X1 U818 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U819 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n759) );
  XNOR2_X1 U820 ( .A(n757), .B(KEYINPUT91), .ZN(n758) );
  XNOR2_X1 U821 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n763) );
  XNOR2_X1 U822 ( .A(n761), .B(KEYINPUT57), .ZN(n762) );
  INV_X1 U823 ( .A(n385), .ZN(n769) );
  NAND2_X1 U824 ( .A1(n770), .A2(n769), .ZN(n775) );
  NAND2_X1 U825 ( .A1(G953), .A2(G224), .ZN(n771) );
  XNOR2_X1 U826 ( .A(KEYINPUT61), .B(n771), .ZN(n773) );
  NAND2_X1 U827 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U828 ( .A1(n775), .A2(n774), .ZN(n781) );
  XOR2_X1 U829 ( .A(n777), .B(n776), .Z(n778) );
  NOR2_X1 U830 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U831 ( .A(n781), .B(n780), .ZN(G69) );
  XNOR2_X1 U832 ( .A(n782), .B(KEYINPUT123), .ZN(n784) );
  XNOR2_X1 U833 ( .A(n783), .B(n784), .ZN(n789) );
  XNOR2_X1 U834 ( .A(n785), .B(n789), .ZN(n787) );
  NAND2_X1 U835 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U836 ( .A(n788), .B(KEYINPUT124), .ZN(n793) );
  XNOR2_X1 U837 ( .A(G227), .B(n789), .ZN(n790) );
  NAND2_X1 U838 ( .A1(n790), .A2(G900), .ZN(n791) );
  NAND2_X1 U839 ( .A1(G953), .A2(n791), .ZN(n792) );
  NAND2_X1 U840 ( .A1(n793), .A2(n792), .ZN(G72) );
  XOR2_X1 U841 ( .A(G137), .B(KEYINPUT126), .Z(n794) );
  XNOR2_X1 U842 ( .A(n795), .B(n794), .ZN(G39) );
  XNOR2_X1 U843 ( .A(n796), .B(G131), .ZN(n797) );
  XNOR2_X1 U844 ( .A(n797), .B(KEYINPUT127), .ZN(G33) );
  XNOR2_X1 U845 ( .A(n409), .B(KEYINPUT125), .ZN(n798) );
endmodule

