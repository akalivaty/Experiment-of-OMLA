//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n562,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n601, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1204, new_n1205, new_n1206, new_n1207;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n454), .A2(G567), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT66), .ZN(new_n458));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n451), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT67), .Z(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n462), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(G137), .ZN(new_n471));
  NAND2_X1  g046(.A1(G101), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n467), .A2(new_n462), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  INV_X1    g054(.A(G100), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n480), .A2(new_n462), .A3(KEYINPUT68), .ZN(new_n481));
  AOI21_X1  g056(.A(KEYINPUT68), .B1(new_n480), .B2(new_n462), .ZN(new_n482));
  OAI221_X1 g057(.A(G2104), .B1(G112), .B2(new_n462), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  AND3_X1   g058(.A1(new_n477), .A2(new_n479), .A3(new_n483), .ZN(G162));
  OAI21_X1  g059(.A(G2104), .B1(new_n462), .B2(G114), .ZN(new_n485));
  NOR2_X1   g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(G126), .A2(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n465), .B2(new_n466), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AND2_X1   g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  NOR2_X1   g066(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n492));
  OAI211_X1 g067(.A(G138), .B(new_n462), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n467), .A2(KEYINPUT4), .A3(G138), .A4(new_n462), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n490), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n500), .A2(G543), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G50), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n506), .A2(new_n510), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n509), .A2(new_n515), .ZN(G166));
  OR2_X1    g091(.A1(KEYINPUT70), .A2(KEYINPUT7), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT70), .A2(KEYINPUT7), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n519), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n517), .A2(new_n521), .A3(new_n518), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n520), .A2(new_n522), .B1(new_n511), .B2(G51), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n504), .A2(G89), .A3(new_n505), .A4(new_n510), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n504), .A2(G63), .A3(G651), .A4(new_n505), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n523), .A2(KEYINPUT71), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n520), .A2(new_n522), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n510), .A2(G51), .A3(G543), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n527), .A2(new_n524), .A3(new_n525), .A4(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n526), .A2(new_n531), .ZN(G168));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n504), .A2(new_n505), .ZN(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n511), .A2(G52), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n506), .A2(G90), .A3(new_n510), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND2_X1  g116(.A1(new_n511), .A2(G43), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n504), .A2(G81), .A3(new_n505), .A4(new_n510), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n534), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n544), .B1(G651), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g125(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n551));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NAND3_X1  g129(.A1(new_n510), .A2(G53), .A3(G543), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT9), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n506), .A2(G91), .A3(new_n510), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n556), .B(new_n557), .C1(new_n558), .C2(new_n508), .ZN(G299));
  INV_X1    g134(.A(G168), .ZN(G286));
  INV_X1    g135(.A(G166), .ZN(G303));
  AND2_X1   g136(.A1(new_n506), .A2(new_n510), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G87), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n511), .A2(G49), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(G288));
  AOI22_X1  g141(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n567), .A2(new_n508), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n511), .A2(G48), .ZN(new_n569));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n513), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G305));
  XOR2_X1   g148(.A(KEYINPUT74), .B(G85), .Z(new_n574));
  AOI22_X1  g149(.A1(new_n562), .A2(new_n574), .B1(G47), .B2(new_n511), .ZN(new_n575));
  NAND2_X1  g150(.A1(G72), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G60), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n534), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n578), .A2(KEYINPUT73), .A3(G651), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(G651), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT73), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n575), .A2(new_n579), .A3(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n585));
  INV_X1    g160(.A(G92), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n513), .B2(new_n586), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n506), .A2(KEYINPUT10), .A3(G92), .A4(new_n510), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G66), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n534), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(G54), .B2(new_n511), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n584), .B1(new_n595), .B2(G868), .ZN(G284));
  OAI21_X1  g171(.A(new_n584), .B1(new_n595), .B2(G868), .ZN(G321));
  NOR2_X1   g172(.A1(G299), .A2(G868), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g174(.A(new_n598), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n595), .B1(new_n601), .B2(G860), .ZN(G148));
  NAND2_X1  g177(.A1(new_n595), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n476), .A2(G2104), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT75), .B(KEYINPUT12), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n607), .B(new_n608), .Z(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT13), .Z(new_n610));
  INV_X1    g185(.A(G2100), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n476), .A2(G135), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT76), .Z(new_n615));
  NAND2_X1  g190(.A1(new_n478), .A2(G123), .ZN(new_n616));
  NOR2_X1   g191(.A1(G99), .A2(G2105), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n615), .B(new_n616), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(G2096), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n612), .A2(new_n613), .A3(new_n621), .ZN(G156));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT78), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2438), .ZN(new_n625));
  XOR2_X1   g200(.A(G2427), .B(G2430), .Z(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n627), .A2(KEYINPUT14), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(G1341), .B(G1348), .Z(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n629), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G14), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n633), .A2(new_n636), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT79), .Z(G401));
  XNOR2_X1  g216(.A(G2072), .B(G2078), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT81), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT17), .Z(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT80), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n648), .B(new_n650), .C1(new_n647), .C2(new_n642), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n649), .A2(new_n646), .A3(new_n642), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT18), .ZN(new_n653));
  INV_X1    g228(.A(new_n645), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n647), .A2(new_n650), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(new_n620), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2100), .ZN(G227));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT82), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1956), .B(G2474), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT83), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1961), .B(G1966), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT85), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n669), .B(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n665), .A2(new_n667), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n663), .A2(new_n668), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n663), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G1986), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  INV_X1    g257(.A(G1981), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n684), .B1(new_n679), .B2(new_n680), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(G229));
  INV_X1    g263(.A(G288), .ZN(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n690), .B2(G23), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT33), .B(G1976), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n690), .A2(G22), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G166), .B2(new_n690), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n694), .B1(new_n696), .B2(G1971), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n690), .A2(G6), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(new_n572), .B2(new_n690), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT32), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n700), .A2(G1981), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(G1981), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n696), .A2(G1971), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n692), .B2(new_n693), .ZN(new_n704));
  NAND4_X1  g279(.A1(new_n697), .A2(new_n701), .A3(new_n702), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT87), .B(KEYINPUT34), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  INV_X1    g283(.A(G290), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G16), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G16), .B2(G24), .ZN(new_n711));
  INV_X1    g286(.A(G1986), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n478), .A2(G119), .ZN(new_n715));
  NOR2_X1   g290(.A1(G95), .A2(G2105), .ZN(new_n716));
  OAI21_X1  g291(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n717));
  INV_X1    g292(.A(G131), .ZN(new_n718));
  OAI221_X1 g293(.A(new_n715), .B1(new_n716), .B2(new_n717), .C1(new_n718), .C2(new_n475), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT86), .B(G29), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  MUX2_X1   g296(.A(G25), .B(new_n719), .S(new_n721), .Z(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT35), .B(G1991), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NOR3_X1   g299(.A1(new_n713), .A2(new_n714), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n707), .A2(new_n708), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT36), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n595), .A2(new_n690), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G4), .B2(new_n690), .ZN(new_n730));
  INV_X1    g305(.A(G1348), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n690), .A2(G20), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT23), .ZN(new_n734));
  INV_X1    g309(.A(G299), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n690), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(G1956), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n730), .A2(new_n731), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n690), .A2(G5), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G171), .B2(new_n690), .ZN(new_n740));
  INV_X1    g315(.A(G1961), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n732), .A2(new_n737), .A3(new_n738), .A4(new_n742), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT25), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n476), .A2(G139), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n467), .A2(G127), .ZN(new_n750));
  NAND2_X1  g325(.A1(G115), .A2(G2104), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n462), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G29), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n754), .B2(G33), .ZN(new_n756));
  INV_X1    g331(.A(G2072), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT91), .B(KEYINPUT31), .Z(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G11), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT92), .B(G28), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(KEYINPUT30), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(KEYINPUT30), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(new_n754), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n760), .B1(new_n762), .B2(new_n764), .C1(new_n619), .C2(new_n720), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n758), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n757), .B2(new_n756), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT88), .B(KEYINPUT24), .Z(new_n768));
  OR2_X1    g343(.A1(new_n768), .A2(G34), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(G34), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n769), .A2(new_n720), .A3(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(G160), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(new_n754), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(G2084), .Z(new_n774));
  NAND3_X1  g349(.A1(new_n467), .A2(G140), .A3(new_n462), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n467), .A2(G128), .A3(G2105), .ZN(new_n776));
  OR2_X1    g351(.A1(G104), .A2(G2105), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n777), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G29), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n720), .A2(G26), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT28), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G2067), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n690), .A2(G19), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n548), .B2(new_n690), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1341), .ZN(new_n787));
  NOR4_X1   g362(.A1(new_n767), .A2(new_n774), .A3(new_n784), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n721), .A2(G35), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G162), .B2(new_n721), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n792), .A2(G2090), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT27), .B(G1996), .ZN(new_n794));
  OR2_X1    g369(.A1(KEYINPUT89), .A2(KEYINPUT26), .ZN(new_n795));
  NAND2_X1  g370(.A1(KEYINPUT89), .A2(KEYINPUT26), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n795), .A2(new_n798), .A3(new_n796), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n478), .A2(G129), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n467), .A2(G141), .A3(new_n462), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n802), .A2(new_n803), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(new_n754), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT90), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G29), .B2(G32), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n793), .B1(new_n794), .B2(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n809), .A2(new_n794), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n721), .A2(G27), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G164), .B2(new_n721), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(G2078), .Z(new_n814));
  NAND4_X1  g389(.A1(new_n788), .A2(new_n810), .A3(new_n811), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n792), .A2(G2090), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT94), .ZN(new_n817));
  NOR2_X1   g392(.A1(G16), .A2(G21), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G168), .B2(G16), .ZN(new_n819));
  INV_X1    g394(.A(G1966), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n817), .A2(new_n821), .ZN(new_n822));
  NOR4_X1   g397(.A1(new_n728), .A2(new_n743), .A3(new_n815), .A4(new_n822), .ZN(G311));
  OR4_X1    g398(.A1(new_n728), .A2(new_n743), .A3(new_n815), .A4(new_n822), .ZN(G150));
  NAND2_X1  g399(.A1(G80), .A2(G543), .ZN(new_n825));
  INV_X1    g400(.A(G67), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n534), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G651), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n504), .A2(G93), .A3(new_n505), .A4(new_n510), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n510), .A2(G55), .A3(G543), .ZN(new_n830));
  AND3_X1   g405(.A1(new_n829), .A2(KEYINPUT95), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(KEYINPUT95), .B1(new_n829), .B2(new_n830), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n828), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n548), .B(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT38), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n595), .A2(G559), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n838), .A2(new_n839), .A3(G860), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n833), .A2(G860), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n840), .A2(new_n842), .ZN(G145));
  XNOR2_X1  g418(.A(new_n619), .B(G160), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G162), .ZN(new_n845));
  OAI21_X1  g420(.A(KEYINPUT96), .B1(new_n487), .B2(new_n489), .ZN(new_n846));
  OAI211_X1 g421(.A(G126), .B(G2105), .C1(new_n491), .C2(new_n492), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT96), .ZN(new_n848));
  OR2_X1    g423(.A1(G102), .A2(G2105), .ZN(new_n849));
  INV_X1    g424(.A(G114), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G2105), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n849), .A2(new_n851), .A3(G2104), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n847), .A2(new_n848), .A3(new_n852), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n846), .A2(new_n495), .A3(new_n496), .A4(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n779), .A2(KEYINPUT97), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT97), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n775), .A2(new_n776), .A3(new_n857), .A4(new_n778), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n806), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n856), .A2(new_n806), .A3(new_n858), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n855), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n861), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n863), .A2(new_n859), .A3(new_n854), .ZN(new_n864));
  INV_X1    g439(.A(new_n753), .ZN(new_n865));
  NOR3_X1   g440(.A1(new_n862), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT98), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(new_n862), .B2(new_n864), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n860), .A2(new_n855), .A3(new_n861), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n854), .B1(new_n863), .B2(new_n859), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT98), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n753), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n867), .B1(new_n873), .B2(KEYINPUT99), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT98), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT98), .B1(new_n870), .B2(new_n871), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n865), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT99), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n609), .B1(new_n874), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n866), .B1(new_n877), .B2(new_n878), .ZN(new_n881));
  INV_X1    g456(.A(new_n609), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n873), .A2(KEYINPUT99), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n719), .B(KEYINPUT100), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n478), .A2(G130), .ZN(new_n886));
  NOR2_X1   g461(.A1(G106), .A2(G2105), .ZN(new_n887));
  OAI21_X1  g462(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n888));
  INV_X1    g463(.A(G142), .ZN(new_n889));
  OAI221_X1 g464(.A(new_n886), .B1(new_n887), .B2(new_n888), .C1(new_n889), .C2(new_n475), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n885), .B(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n880), .A2(new_n884), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n891), .B1(new_n880), .B2(new_n884), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n845), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  INV_X1    g471(.A(new_n891), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n874), .A2(new_n879), .A3(new_n609), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n882), .B1(new_n881), .B2(new_n883), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n845), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n901), .A3(new_n892), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n895), .A2(new_n896), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g479(.A1(new_n594), .A2(new_n735), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n589), .A2(G299), .A3(new_n593), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT101), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n907), .B(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n548), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n833), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n548), .B(new_n828), .C1(new_n832), .C2(new_n831), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n603), .B(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  INV_X1    g491(.A(new_n906), .ZN(new_n917));
  AOI21_X1  g492(.A(G299), .B1(new_n589), .B2(new_n593), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n905), .A2(KEYINPUT41), .A3(new_n906), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n915), .B1(new_n914), .B2(new_n921), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n922), .A2(KEYINPUT42), .ZN(new_n923));
  XNOR2_X1  g498(.A(G290), .B(new_n572), .ZN(new_n924));
  XNOR2_X1  g499(.A(G166), .B(G288), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n924), .B(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n922), .A2(KEYINPUT42), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n923), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n927), .B1(new_n923), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g505(.A(G868), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(G868), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n833), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(G295));
  INV_X1    g509(.A(KEYINPUT102), .ZN(new_n935));
  XNOR2_X1  g510(.A(G295), .B(new_n935), .ZN(G331));
  NAND2_X1  g511(.A1(G301), .A2(KEYINPUT103), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n537), .A2(new_n938), .A3(new_n538), .A4(new_n539), .ZN(new_n939));
  NAND3_X1  g514(.A1(G168), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(G301), .A2(new_n526), .A3(new_n531), .A4(KEYINPUT103), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT104), .B1(new_n942), .B2(new_n913), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n913), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n834), .A2(new_n945), .A3(new_n941), .A4(new_n940), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n943), .A2(new_n907), .A3(new_n944), .A4(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n942), .A2(new_n913), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n834), .B1(new_n941), .B2(new_n940), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n921), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n926), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT105), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n926), .A2(new_n947), .A3(new_n950), .A4(new_n953), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n952), .A2(new_n896), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n919), .A2(KEYINPUT106), .A3(new_n920), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n907), .A2(new_n959), .A3(new_n916), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n944), .A2(new_n946), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n961), .B1(new_n962), .B2(new_n943), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n909), .A2(new_n948), .A3(new_n949), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n927), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n955), .A2(new_n956), .A3(new_n957), .A4(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(G37), .B1(new_n951), .B2(KEYINPUT105), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n965), .A2(new_n967), .A3(new_n957), .A4(new_n954), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT107), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n947), .A2(new_n950), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n927), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n967), .A2(new_n954), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n966), .A2(new_n969), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n955), .A2(new_n957), .A3(new_n971), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n955), .A2(new_n965), .ZN(new_n978));
  OAI211_X1 g553(.A(KEYINPUT44), .B(new_n977), .C1(new_n978), .C2(new_n957), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n979), .A2(new_n980), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n976), .B1(new_n981), .B2(new_n982), .ZN(G397));
  AND2_X1   g558(.A1(G160), .A2(G40), .ZN(new_n984));
  XNOR2_X1  g559(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n986), .B1(new_n854), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n984), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(G290), .A2(G1986), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  XOR2_X1   g567(.A(new_n779), .B(G2067), .Z(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n806), .B(G1996), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g571(.A(new_n719), .B(new_n723), .Z(new_n997));
  NAND3_X1  g572(.A1(new_n992), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n709), .A2(new_n712), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n990), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n497), .A2(new_n987), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n985), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n854), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n984), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  XOR2_X1   g579(.A(KEYINPUT110), .B(G1971), .Z(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g581(.A(new_n1006), .B(KEYINPUT111), .Z(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT114), .B(G2090), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n854), .A2(new_n987), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n854), .A2(KEYINPUT112), .A3(new_n987), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT113), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1012), .A2(new_n1017), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1001), .A2(KEYINPUT50), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1016), .A2(new_n984), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1007), .B1(new_n1009), .B2(new_n1020), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1021), .A2(G8), .ZN(new_n1022));
  INV_X1    g597(.A(G8), .ZN(new_n1023));
  NOR2_X1   g598(.A1(G166), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1024), .B(KEYINPUT55), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT49), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n572), .A2(new_n683), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n572), .A2(new_n683), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1026), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1029), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1031), .A2(KEYINPUT49), .A3(new_n1027), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1012), .A2(new_n984), .A3(new_n1014), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1033), .A2(G8), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1030), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n689), .A2(G1976), .ZN(new_n1036));
  INV_X1    g611(.A(G1976), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT52), .B1(G288), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1034), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1040), .B1(KEYINPUT52), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1022), .A2(new_n1025), .A3(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1035), .A2(new_n1037), .A3(new_n689), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1034), .B1(new_n1044), .B2(new_n1028), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1021), .A2(G8), .A3(new_n1025), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1047), .A2(new_n1042), .ZN(new_n1048));
  NAND2_X1  g623(.A1(G160), .A2(G40), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(G2084), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1016), .A2(new_n1018), .A3(new_n1019), .A4(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT45), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n854), .A2(KEYINPUT112), .A3(new_n987), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT112), .B1(new_n854), .B2(new_n987), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(new_n1001), .B2(new_n985), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n497), .A2(KEYINPUT115), .A3(new_n987), .A4(new_n986), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1055), .A2(new_n1059), .A3(new_n984), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n820), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n1023), .B(G286), .C1(new_n1051), .C2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT63), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1048), .B(new_n1065), .C1(new_n1025), .C2(new_n1022), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT50), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1001), .A2(KEYINPUT50), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1068), .A2(new_n1049), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n1008), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1023), .B1(new_n1071), .B2(new_n1006), .ZN(new_n1072));
  OR2_X1    g647(.A1(new_n1072), .A2(new_n1025), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1047), .A2(new_n1042), .A3(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1064), .B1(new_n1074), .B2(new_n1063), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1046), .B1(new_n1066), .B2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(G299), .B(KEYINPUT57), .ZN(new_n1077));
  AOI21_X1  g652(.A(G1956), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT56), .B(G2072), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1004), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1077), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1033), .A2(KEYINPUT116), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1012), .A2(new_n984), .A3(new_n1084), .A4(new_n1014), .ZN(new_n1085));
  AOI21_X1  g660(.A(G2067), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1020), .A2(new_n1087), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1015), .A2(KEYINPUT113), .B1(KEYINPUT50), .B2(new_n1001), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1089), .A2(KEYINPUT117), .A3(new_n984), .A4(new_n1018), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1086), .B1(new_n1091), .B2(new_n731), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1082), .B1(new_n1092), .B2(new_n594), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1078), .A2(new_n1077), .A3(new_n1081), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT118), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1093), .A2(new_n1098), .A3(new_n1095), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1091), .A2(new_n731), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1086), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1100), .A2(KEYINPUT60), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT60), .ZN(new_n1103));
  AOI21_X1  g678(.A(G1348), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1103), .B1(new_n1104), .B2(new_n1086), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1102), .A2(new_n595), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1095), .A2(KEYINPUT61), .A3(new_n1082), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT58), .B(G1341), .Z(new_n1109));
  NAND3_X1  g684(.A1(new_n1083), .A2(new_n1085), .A3(new_n1109), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1004), .A2(G1996), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1108), .B1(new_n1112), .B2(new_n548), .ZN(new_n1113));
  AOI211_X1 g688(.A(KEYINPUT59), .B(new_n910), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1107), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT119), .B(KEYINPUT61), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1082), .B1(new_n1094), .B2(KEYINPUT120), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1118), .B(new_n1077), .C1(new_n1078), .C2(new_n1081), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1116), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1115), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1092), .A2(KEYINPUT60), .A3(new_n594), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1106), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1097), .A2(new_n1099), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1051), .A2(new_n1061), .A3(G168), .ZN(new_n1125));
  AND2_X1   g700(.A1(KEYINPUT121), .A2(G8), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT51), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT51), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1125), .A2(new_n1129), .A3(new_n1126), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1051), .A2(new_n1061), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1131), .A2(G8), .A3(G286), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1128), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(KEYINPUT122), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1128), .A2(new_n1135), .A3(new_n1130), .A4(new_n1132), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT54), .ZN(new_n1138));
  AOI21_X1  g713(.A(G1961), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n984), .A2(new_n1003), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT53), .ZN(new_n1141));
  NOR4_X1   g716(.A1(new_n1140), .A2(new_n988), .A3(new_n1141), .A4(G2078), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1142), .B(KEYINPUT123), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1141), .B1(new_n1004), .B2(G2078), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  NOR4_X1   g720(.A1(new_n1139), .A2(new_n1143), .A3(new_n1145), .A4(G171), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1091), .A2(new_n741), .ZN(new_n1147));
  OR3_X1    g722(.A1(new_n1060), .A2(new_n1141), .A3(G2078), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1148), .A2(new_n1144), .ZN(new_n1149));
  AOI21_X1  g724(.A(G301), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1138), .B1(new_n1146), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1074), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1147), .A2(G301), .A3(new_n1144), .A4(new_n1148), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1139), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1153), .B(KEYINPUT54), .C1(new_n1154), .C2(G301), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1137), .A2(new_n1151), .A3(new_n1152), .A4(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1076), .B1(new_n1124), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT124), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1158), .B1(new_n1137), .B2(KEYINPUT62), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n1160));
  AOI211_X1 g735(.A(KEYINPUT124), .B(new_n1160), .C1(new_n1134), .C2(new_n1136), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1134), .A2(new_n1160), .A3(new_n1136), .ZN(new_n1162));
  AND4_X1   g737(.A1(new_n1073), .A2(new_n1150), .A3(new_n1047), .A4(new_n1042), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1159), .A2(new_n1161), .A3(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1000), .B1(new_n1157), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT46), .ZN(new_n1167));
  OR3_X1    g742(.A1(new_n989), .A2(new_n1167), .A3(G1996), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n990), .B1(new_n806), .B2(new_n994), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1167), .B1(new_n989), .B2(G1996), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  XOR2_X1   g746(.A(new_n1171), .B(KEYINPUT47), .Z(new_n1172));
  NOR2_X1   g747(.A1(new_n992), .A2(new_n989), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(KEYINPUT48), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1173), .A2(KEYINPUT48), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n989), .B1(new_n996), .B2(new_n997), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1172), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n996), .A2(new_n989), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1179), .A2(new_n723), .A3(new_n719), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n779), .A2(G2067), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT125), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n990), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1184), .B1(new_n1183), .B2(new_n1182), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1178), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(new_n1186), .B2(new_n1185), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1166), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g764(.A(G319), .ZN(new_n1191));
  NOR3_X1   g765(.A1(G227), .A2(new_n640), .A3(new_n1191), .ZN(new_n1192));
  OAI21_X1  g766(.A(new_n1192), .B1(new_n686), .B2(new_n687), .ZN(new_n1193));
  NAND2_X1  g767(.A1(new_n900), .A2(new_n892), .ZN(new_n1194));
  AOI21_X1  g768(.A(G37), .B1(new_n1194), .B2(new_n845), .ZN(new_n1195));
  AOI21_X1  g769(.A(new_n1193), .B1(new_n1195), .B2(new_n902), .ZN(new_n1196));
  AOI21_X1  g770(.A(KEYINPUT127), .B1(new_n1196), .B2(new_n974), .ZN(new_n1197));
  OR3_X1    g771(.A1(G227), .A2(new_n640), .A3(new_n1191), .ZN(new_n1198));
  INV_X1    g772(.A(new_n686), .ZN(new_n1199));
  INV_X1    g773(.A(new_n687), .ZN(new_n1200));
  AOI21_X1  g774(.A(new_n1198), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  AND4_X1   g775(.A1(KEYINPUT127), .A2(new_n974), .A3(new_n1201), .A4(new_n903), .ZN(new_n1202));
  NOR2_X1   g776(.A1(new_n1197), .A2(new_n1202), .ZN(G308));
  NAND3_X1  g777(.A1(new_n974), .A2(new_n1201), .A3(new_n903), .ZN(new_n1204));
  INV_X1    g778(.A(KEYINPUT127), .ZN(new_n1205));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g780(.A1(new_n1196), .A2(KEYINPUT127), .A3(new_n974), .ZN(new_n1207));
  NAND2_X1  g781(.A1(new_n1206), .A2(new_n1207), .ZN(G225));
endmodule


