//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT84), .Z(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT92), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n193), .B1(G143), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n194), .A2(G143), .ZN(new_n199));
  OAI22_X1  g013(.A1(new_n195), .A2(new_n196), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT64), .B1(new_n197), .B2(G146), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(new_n194), .A3(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n197), .A2(G146), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n196), .A2(KEYINPUT1), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n201), .A2(new_n203), .A3(new_n204), .A4(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n200), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G125), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT87), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT0), .A2(G128), .ZN(new_n210));
  OR2_X1    g024(.A1(KEYINPUT0), .A2(G128), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n210), .B(new_n211), .C1(new_n198), .C2(new_n199), .ZN(new_n212));
  INV_X1    g026(.A(new_n210), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n201), .A2(new_n203), .A3(new_n204), .A4(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G125), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n208), .B1(new_n209), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n216), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT87), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G224), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(G953), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n220), .B(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G110), .B(G122), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n226));
  INV_X1    g040(.A(G104), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT3), .B1(new_n227), .B2(G107), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT81), .ZN(new_n229));
  INV_X1    g043(.A(G107), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G104), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT81), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n232), .A3(KEYINPUT3), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n227), .A2(G107), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n235), .B1(new_n231), .B2(KEYINPUT3), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n226), .B1(new_n238), .B2(G101), .ZN(new_n239));
  INV_X1    g053(.A(G101), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n234), .A2(new_n240), .A3(new_n237), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT82), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n236), .B1(new_n233), .B2(new_n229), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT82), .B1(new_n244), .B2(new_n240), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n239), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G119), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G116), .ZN(new_n248));
  INV_X1    g062(.A(G116), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G119), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT2), .B(G113), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n251), .A2(new_n253), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n251), .A2(new_n253), .A3(KEYINPUT67), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n244), .A2(KEYINPUT4), .A3(new_n240), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n246), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n240), .B1(new_n231), .B2(new_n235), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n241), .A2(new_n242), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n244), .A2(KEYINPUT82), .A3(new_n240), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(KEYINPUT85), .A2(KEYINPUT5), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT85), .A2(KEYINPUT5), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(G113), .B1(new_n272), .B2(new_n248), .ZN(new_n273));
  INV_X1    g087(.A(new_n271), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n248), .B(new_n250), .C1(new_n274), .C2(new_n269), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n255), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n268), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n225), .B1(new_n264), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n266), .A2(new_n267), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n262), .B1(new_n282), .B2(new_n239), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n283), .A2(new_n261), .B1(new_n268), .B2(new_n278), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT86), .B1(new_n284), .B2(new_n225), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n264), .A2(KEYINPUT86), .A3(new_n279), .A4(new_n225), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n281), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT6), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT6), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n281), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n224), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n217), .A2(KEYINPUT7), .A3(new_n219), .A4(new_n223), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT90), .B(KEYINPUT7), .Z(new_n294));
  OAI22_X1  g108(.A1(new_n218), .A2(new_n208), .B1(new_n222), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n252), .A2(KEYINPUT88), .A3(KEYINPUT5), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT88), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT5), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n297), .B1(new_n251), .B2(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n296), .B(new_n299), .C1(new_n273), .C2(KEYINPUT89), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n273), .A2(KEYINPUT89), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n255), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n302), .A2(new_n268), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n225), .B(KEYINPUT8), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n304), .B1(new_n268), .B2(new_n277), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n293), .B(new_n295), .C1(new_n303), .C2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n307), .B1(new_n285), .B2(new_n287), .ZN(new_n308));
  INV_X1    g122(.A(G902), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(KEYINPUT91), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT91), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n264), .A2(new_n279), .A3(new_n225), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT86), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n306), .B1(new_n314), .B2(new_n286), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n311), .B1(new_n315), .B2(G902), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n192), .B1(new_n292), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n280), .B1(new_n314), .B2(new_n286), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n291), .B1(new_n319), .B2(new_n290), .ZN(new_n320));
  INV_X1    g134(.A(new_n224), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n322), .A2(new_n316), .A3(new_n310), .A4(new_n191), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n188), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n197), .A2(G128), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n196), .A2(G143), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G134), .ZN(new_n328));
  INV_X1    g142(.A(G134), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n325), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT98), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n249), .A2(G122), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n249), .A2(G122), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n334), .B1(new_n335), .B2(KEYINPUT14), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(KEYINPUT14), .B2(new_n334), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G107), .ZN(new_n338));
  XNOR2_X1  g152(.A(G116), .B(G122), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n230), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n328), .A2(KEYINPUT98), .A3(new_n330), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n333), .A2(new_n338), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n339), .B(new_n230), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n196), .A2(G143), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n344), .B1(KEYINPUT13), .B2(new_n326), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n344), .A2(KEYINPUT13), .ZN(new_n346));
  OAI21_X1  g160(.A(G134), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n343), .A2(new_n347), .A3(new_n330), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n342), .A2(new_n348), .ZN(new_n349));
  XOR2_X1   g163(.A(KEYINPUT9), .B(G234), .Z(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(KEYINPUT80), .ZN(new_n351));
  INV_X1    g165(.A(G953), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(G217), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT99), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n349), .A2(KEYINPUT99), .A3(new_n353), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n349), .A2(new_n353), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G478), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(KEYINPUT15), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n359), .A2(KEYINPUT100), .A3(new_n309), .A4(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n359), .A2(new_n309), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT100), .ZN(new_n364));
  OAI22_X1  g178(.A1(new_n363), .A2(new_n364), .B1(KEYINPUT15), .B2(new_n360), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT100), .B1(new_n359), .B2(new_n309), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n362), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n352), .A2(G952), .ZN(new_n368));
  NAND2_X1  g182(.A1(G234), .A2(G237), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n369), .A2(G902), .A3(G953), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT21), .B(G898), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n367), .A2(new_n374), .ZN(new_n375));
  NOR3_X1   g189(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G113), .B(G122), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(new_n227), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT18), .ZN(new_n380));
  INV_X1    g194(.A(G131), .ZN(new_n381));
  NOR3_X1   g195(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT93), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT69), .B(G237), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(G214), .A3(new_n352), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(new_n197), .ZN(new_n385));
  OR2_X1    g199(.A1(KEYINPUT69), .A2(G237), .ZN(new_n386));
  NAND2_X1  g200(.A1(KEYINPUT69), .A2(G237), .ZN(new_n387));
  AOI21_X1  g201(.A(G953), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(G143), .B1(new_n388), .B2(G214), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n382), .B1(new_n385), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n384), .A2(new_n197), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(G143), .A3(G214), .ZN(new_n392));
  INV_X1    g206(.A(new_n382), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G140), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G125), .ZN(new_n396));
  INV_X1    g210(.A(G125), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G140), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT77), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G125), .B(G140), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT77), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n401), .A2(new_n403), .A3(new_n194), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n404), .B1(new_n194), .B2(new_n402), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n390), .A2(new_n394), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT94), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n390), .A2(new_n405), .A3(KEYINPUT94), .A4(new_n394), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT65), .B(G131), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n412), .B1(new_n385), .B2(new_n389), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n391), .A2(new_n411), .A3(new_n392), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n396), .A2(KEYINPUT16), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n416), .B1(new_n402), .B2(KEYINPUT16), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G146), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT19), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n401), .A2(new_n403), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT95), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n402), .B2(new_n419), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n399), .A2(KEYINPUT95), .A3(KEYINPUT19), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n420), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n415), .B(new_n418), .C1(G146), .C2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n379), .B1(new_n410), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT17), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n413), .A2(new_n428), .A3(new_n414), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT96), .ZN(new_n430));
  OAI21_X1  g244(.A(KEYINPUT76), .B1(new_n417), .B2(G146), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT76), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n402), .A2(KEYINPUT16), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n432), .B(new_n194), .C1(new_n433), .C2(new_n416), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n431), .A2(new_n434), .A3(new_n418), .ZN(new_n435));
  AOI211_X1 g249(.A(new_n428), .B(new_n411), .C1(new_n391), .C2(new_n392), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT96), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n413), .A2(new_n438), .A3(new_n428), .A4(new_n414), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n430), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(new_n379), .A3(new_n410), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n377), .B1(new_n427), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT97), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n440), .A2(new_n379), .A3(new_n410), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n443), .B1(new_n444), .B2(new_n426), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n427), .A2(KEYINPUT97), .A3(new_n441), .ZN(new_n446));
  NOR2_X1   g260(.A1(G475), .A2(G902), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n442), .B1(new_n448), .B2(KEYINPUT20), .ZN(new_n449));
  INV_X1    g263(.A(G475), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n379), .B1(new_n440), .B2(new_n410), .ZN(new_n451));
  OR2_X1    g265(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n450), .B1(new_n452), .B2(new_n309), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n375), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G221), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(new_n351), .B2(new_n309), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT11), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n329), .B2(G137), .ZN(new_n458));
  INV_X1    g272(.A(G137), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(KEYINPUT11), .A3(G134), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n329), .A2(G137), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n412), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT66), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n458), .A2(new_n460), .A3(KEYINPUT66), .A4(new_n461), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n464), .B1(new_n468), .B2(new_n381), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n201), .A2(new_n203), .A3(new_n204), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n470), .B1(new_n196), .B2(new_n195), .ZN(new_n471));
  AOI221_X4 g285(.A(new_n265), .B1(new_n206), .B2(new_n471), .C1(new_n266), .C2(new_n267), .ZN(new_n472));
  INV_X1    g286(.A(new_n265), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n207), .B1(new_n282), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n469), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT12), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g291(.A(KEYINPUT12), .B(new_n469), .C1(new_n472), .C2(new_n474), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n471), .A2(new_n206), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n282), .A2(new_n473), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT10), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n215), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n246), .A2(new_n484), .A3(new_n263), .ZN(new_n485));
  INV_X1    g299(.A(new_n469), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n200), .A2(new_n206), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(new_n482), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n268), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n483), .A2(new_n485), .A3(new_n486), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n479), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(G110), .B(G140), .ZN(new_n492));
  INV_X1    g306(.A(G227), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(G953), .ZN(new_n494));
  XOR2_X1   g308(.A(new_n492), .B(new_n494), .Z(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n283), .A2(new_n484), .B1(new_n268), .B2(new_n488), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n486), .B1(new_n497), .B2(new_n483), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n490), .A2(new_n495), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n491), .A2(new_n496), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(G469), .B1(new_n502), .B2(G902), .ZN(new_n503));
  INV_X1    g317(.A(new_n490), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n496), .B1(new_n498), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n490), .A2(KEYINPUT83), .A3(new_n495), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n479), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT83), .B1(new_n490), .B2(new_n495), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G469), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n510), .A3(new_n309), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n456), .B1(new_n503), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n324), .A2(new_n454), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT79), .ZN(new_n514));
  INV_X1    g328(.A(G472), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n381), .B1(new_n466), .B2(new_n467), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n484), .B1(new_n516), .B2(new_n463), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n459), .A2(G134), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n518), .A2(new_n461), .ZN(new_n519));
  OAI22_X1  g333(.A1(new_n412), .A2(new_n462), .B1(new_n519), .B2(new_n381), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT68), .ZN(new_n521));
  NOR3_X1   g335(.A1(new_n487), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n381), .B1(new_n518), .B2(new_n461), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n523), .B1(new_n524), .B2(new_n411), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT68), .B1(new_n525), .B2(new_n207), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n517), .B(new_n260), .C1(new_n522), .C2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n525), .A2(new_n207), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n517), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n521), .B1(new_n487), .B2(new_n520), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n525), .A2(KEYINPUT68), .A3(new_n207), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n469), .A2(new_n484), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n531), .B1(new_n534), .B2(new_n529), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n528), .B1(new_n535), .B2(new_n261), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n388), .A2(G210), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(KEYINPUT27), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT26), .B(G101), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT72), .B1(new_n536), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT71), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n517), .A2(new_n530), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n527), .A2(new_n542), .B1(new_n261), .B2(new_n543), .ZN(new_n544));
  AOI211_X1 g358(.A(KEYINPUT71), .B(new_n260), .C1(new_n517), .C2(new_n530), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT28), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT70), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n540), .B(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT28), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n543), .B2(new_n261), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n546), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n532), .A2(new_n533), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n529), .B1(new_n552), .B2(new_n517), .ZN(new_n553));
  INV_X1    g367(.A(new_n531), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n261), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n527), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT72), .ZN(new_n557));
  INV_X1    g371(.A(new_n540), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT29), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n541), .A2(new_n551), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n550), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n534), .B(new_n260), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n562), .B1(new_n563), .B2(KEYINPUT28), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n558), .A2(new_n560), .ZN(new_n565));
  AOI21_X1  g379(.A(G902), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n515), .B1(new_n561), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT31), .B1(new_n536), .B2(new_n540), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n555), .A2(KEYINPUT31), .A3(new_n527), .A4(new_n540), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n548), .B1(new_n546), .B2(new_n550), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n515), .B(new_n309), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT32), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n555), .A2(new_n527), .A3(new_n540), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT31), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n569), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n527), .A2(new_n542), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n543), .A2(new_n261), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n545), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n550), .B1(new_n581), .B2(new_n549), .ZN(new_n582));
  INV_X1    g396(.A(new_n548), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(G902), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT32), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n586), .A3(new_n515), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n567), .B1(new_n574), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT25), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(KEYINPUT78), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT74), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n591), .A2(new_n592), .B1(new_n247), .B2(G128), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n196), .A2(G119), .ZN(new_n594));
  AND2_X1   g408(.A1(KEYINPUT75), .A2(KEYINPUT23), .ZN(new_n595));
  NOR2_X1   g409(.A1(KEYINPUT75), .A2(KEYINPUT23), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n593), .B(new_n597), .C1(new_n592), .C2(new_n591), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(G110), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n247), .A2(G128), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT24), .B(G110), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT73), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n435), .A2(new_n599), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n601), .A2(new_n602), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n606), .B1(new_n598), .B2(G110), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(new_n418), .A3(new_n404), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT22), .B(G137), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n352), .A2(G221), .A3(G234), .ZN(new_n611));
  XOR2_X1   g425(.A(new_n610), .B(new_n611), .Z(new_n612));
  NOR2_X1   g426(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n612), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n605), .B2(new_n608), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n590), .B1(new_n616), .B2(G902), .ZN(new_n617));
  OAI221_X1 g431(.A(new_n309), .B1(KEYINPUT78), .B2(new_n589), .C1(new_n613), .C2(new_n615), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n617), .A2(new_n618), .B1(KEYINPUT78), .B2(new_n589), .ZN(new_n619));
  INV_X1    g433(.A(G217), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(G234), .B2(new_n309), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n616), .A2(G902), .A3(new_n621), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n514), .B1(new_n588), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n567), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n586), .B1(new_n585), .B2(new_n515), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n577), .A2(new_n569), .B1(new_n582), .B2(new_n583), .ZN(new_n629));
  NOR4_X1   g443(.A1(new_n629), .A2(KEYINPUT32), .A3(G472), .A4(G902), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n627), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n623), .A2(new_n624), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n631), .A2(KEYINPUT79), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n513), .B1(new_n626), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(new_n240), .ZN(G3));
  NAND4_X1  g449(.A1(new_n322), .A2(new_n316), .A3(new_n310), .A4(new_n189), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT101), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n322), .A2(new_n316), .A3(new_n310), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n190), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n638), .A2(KEYINPUT101), .A3(new_n190), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n188), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(G472), .B1(new_n629), .B2(G902), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n573), .A2(new_n643), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n512), .A2(new_n644), .A3(new_n632), .ZN(new_n645));
  INV_X1    g459(.A(new_n453), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n448), .A2(KEYINPUT20), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n646), .B1(new_n647), .B2(new_n442), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n363), .A2(new_n360), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT33), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n359), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n358), .A2(KEYINPUT33), .A3(new_n354), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n309), .A2(G478), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n648), .A2(new_n374), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n642), .A2(new_n645), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT34), .B(G104), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  NAND2_X1  g474(.A1(new_n448), .A2(KEYINPUT20), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n445), .A2(new_n446), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n661), .B1(new_n663), .B2(new_n377), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n646), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n665), .A2(new_n367), .A3(new_n373), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n642), .A2(new_n645), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT35), .B(G107), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  NOR2_X1   g483(.A1(new_n614), .A2(KEYINPUT36), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n609), .B(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n621), .A2(G902), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n673), .B1(new_n619), .B2(new_n622), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n644), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n675), .A2(new_n324), .A3(new_n454), .A4(new_n512), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT37), .B(G110), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G12));
  NAND2_X1  g492(.A1(new_n631), .A2(new_n674), .ZN(new_n679));
  INV_X1    g493(.A(new_n367), .ZN(new_n680));
  INV_X1    g494(.A(G900), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n370), .B1(new_n371), .B2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n664), .A2(new_n646), .A3(new_n680), .A4(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n512), .A3(new_n642), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  INV_X1    g501(.A(new_n188), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n574), .A2(new_n587), .ZN(new_n689));
  INV_X1    g503(.A(new_n575), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n690), .B1(new_n583), .B2(new_n563), .ZN(new_n691));
  OAI21_X1  g505(.A(G472), .B1(new_n691), .B2(G902), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n674), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n449), .A2(new_n453), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n367), .ZN(new_n696));
  AND4_X1   g510(.A1(new_n688), .A2(new_n693), .A3(new_n694), .A4(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n682), .B(KEYINPUT39), .Z(new_n698));
  NAND2_X1  g512(.A1(new_n512), .A2(new_n698), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n699), .A2(KEYINPUT40), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(KEYINPUT40), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n318), .A2(new_n323), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT38), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n697), .A2(new_n700), .A3(new_n701), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G143), .ZN(G45));
  NOR2_X1   g519(.A1(new_n588), .A2(new_n694), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n648), .A2(new_n655), .A3(new_n683), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n642), .A2(new_n512), .A3(new_n706), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  INV_X1    g524(.A(KEYINPUT103), .ZN(new_n711));
  NAND2_X1  g525(.A1(KEYINPUT102), .A2(G469), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT83), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n500), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n506), .A3(new_n479), .ZN(new_n716));
  AOI211_X1 g530(.A(G902), .B(new_n713), .C1(new_n716), .C2(new_n505), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n712), .B1(new_n509), .B2(new_n309), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n456), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n711), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR4_X1   g535(.A1(new_n717), .A2(new_n718), .A3(KEYINPUT103), .A4(new_n456), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n631), .A2(new_n632), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n723), .A2(new_n725), .A3(new_n642), .A4(new_n657), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT41), .B(G113), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT104), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n726), .B(new_n728), .ZN(G15));
  NAND4_X1  g543(.A1(new_n723), .A2(new_n725), .A3(new_n642), .A4(new_n666), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G116), .ZN(G18));
  NAND4_X1  g545(.A1(new_n723), .A2(new_n642), .A3(new_n454), .A4(new_n706), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G119), .ZN(G21));
  OAI21_X1  g547(.A(new_n578), .B1(new_n548), .B2(new_n564), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n515), .A3(new_n309), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n643), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n625), .A2(new_n736), .A3(new_n373), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n723), .A2(new_n642), .A3(new_n696), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  NAND3_X1  g553(.A1(new_n735), .A2(new_n643), .A3(new_n674), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n707), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n723), .A2(new_n642), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G125), .ZN(G27));
  AND3_X1   g557(.A1(new_n318), .A2(new_n688), .A3(new_n323), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n491), .A2(new_n496), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n501), .A2(new_n499), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(G469), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(G469), .A2(G902), .ZN(new_n748));
  XOR2_X1   g562(.A(new_n748), .B(KEYINPUT105), .Z(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  AOI211_X1 g564(.A(G469), .B(G902), .C1(new_n716), .C2(new_n505), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n720), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT106), .B1(new_n744), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n318), .A2(new_n688), .A3(new_n323), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n755), .A2(new_n752), .A3(new_n756), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n725), .B(new_n708), .C1(new_n754), .C2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT42), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n744), .A2(new_n753), .A3(KEYINPUT106), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n756), .B1(new_n755), .B2(new_n752), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n724), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(KEYINPUT42), .A3(new_n708), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G131), .ZN(G33));
  INV_X1    g580(.A(new_n684), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT107), .B1(new_n763), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n763), .A2(KEYINPUT107), .A3(new_n767), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  INV_X1    g586(.A(new_n749), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n502), .B(KEYINPUT45), .Z(new_n774));
  AOI21_X1  g588(.A(new_n773), .B1(new_n774), .B2(G469), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n751), .B1(new_n775), .B2(KEYINPUT46), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n776), .B1(KEYINPUT46), .B2(new_n775), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n720), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n779), .A2(new_n698), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n695), .A2(new_n655), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT43), .ZN(new_n783));
  OR3_X1    g597(.A1(new_n783), .A2(new_n644), .A3(new_n694), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n780), .B1(new_n781), .B2(new_n784), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n784), .A2(new_n781), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n785), .A2(new_n755), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(new_n459), .ZN(G39));
  INV_X1    g602(.A(KEYINPUT47), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n789), .A2(KEYINPUT108), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(KEYINPUT108), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n779), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n778), .A2(KEYINPUT108), .A3(new_n789), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n707), .A2(new_n631), .A3(new_n755), .A4(new_n632), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G140), .ZN(G42));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n645), .A2(new_n324), .A3(new_n657), .ZN(new_n799));
  OAI21_X1  g613(.A(KEYINPUT110), .B1(new_n634), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT111), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n449), .A2(new_n367), .A3(new_n453), .A4(new_n373), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n324), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n645), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n801), .B1(new_n324), .B2(new_n802), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n676), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n324), .A2(new_n454), .A3(new_n512), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n588), .A2(new_n514), .A3(new_n625), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT79), .B1(new_n631), .B2(new_n632), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT110), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n645), .A2(new_n657), .A3(new_n324), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n800), .A2(new_n807), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT112), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n800), .A2(new_n807), .A3(new_n814), .A4(KEYINPUT112), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n741), .B1(new_n754), .B2(new_n757), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n665), .A2(new_n680), .A3(new_n682), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n706), .A2(new_n512), .A3(new_n821), .A4(new_n744), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n769), .B2(new_n770), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n726), .A2(new_n730), .A3(new_n732), .A4(new_n738), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(new_n760), .B2(new_n764), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n819), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n694), .A2(new_n683), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(new_n689), .B2(new_n692), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n642), .A2(new_n696), .A3(new_n829), .A4(new_n753), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n686), .A2(new_n709), .A3(new_n830), .A4(new_n742), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n679), .A2(new_n707), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n512), .B(new_n642), .C1(new_n834), .C2(new_n685), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n835), .A2(KEYINPUT52), .A3(new_n742), .A4(new_n830), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT113), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n833), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n798), .B1(new_n827), .B2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n811), .A2(new_n813), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n806), .B1(new_n844), .B2(KEYINPUT110), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT112), .B1(new_n845), .B2(new_n814), .ZN(new_n846));
  AND4_X1   g660(.A1(KEYINPUT112), .A2(new_n800), .A3(new_n814), .A4(new_n807), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n824), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n732), .A2(new_n738), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT114), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n849), .A2(new_n850), .A3(new_n726), .A4(new_n730), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n825), .A2(KEYINPUT114), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n798), .B1(new_n760), .B2(new_n764), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n837), .A2(new_n851), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n848), .A2(new_n854), .A3(KEYINPUT115), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n833), .A2(new_n836), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n823), .ZN(new_n860));
  INV_X1    g674(.A(new_n770), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n860), .B1(new_n861), .B2(new_n768), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n817), .B2(new_n818), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n856), .B1(new_n859), .B2(new_n863), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n842), .B(new_n843), .C1(new_n855), .C2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n863), .A2(new_n826), .A3(new_n838), .A4(new_n840), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT53), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n863), .A2(new_n798), .A3(new_n826), .A4(new_n837), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n867), .A2(KEYINPUT54), .A3(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n865), .A2(new_n869), .A3(KEYINPUT116), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n723), .A2(new_n744), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT118), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n648), .A2(new_n655), .ZN(new_n873));
  INV_X1    g687(.A(new_n370), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n693), .A2(new_n625), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n723), .A2(new_n642), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n783), .A2(new_n874), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n625), .A2(new_n736), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n876), .B(new_n368), .C1(new_n877), .C2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n872), .A2(new_n725), .A3(new_n878), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n882), .A2(KEYINPUT48), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(KEYINPUT48), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n880), .A2(new_n755), .ZN(new_n886));
  INV_X1    g700(.A(new_n719), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(new_n720), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n886), .B1(new_n794), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n648), .A2(new_n655), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n872), .A2(new_n875), .A3(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n703), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(new_n188), .A3(new_n723), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n880), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT50), .ZN(new_n895));
  INV_X1    g709(.A(new_n740), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n872), .A2(new_n896), .A3(new_n878), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n889), .A2(new_n891), .A3(new_n895), .A4(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT117), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT51), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT51), .B1(new_n898), .B2(new_n899), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n885), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT116), .B1(new_n865), .B2(new_n869), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n870), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(G952), .A2(G953), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n632), .A2(new_n688), .A3(new_n720), .ZN(new_n906));
  AOI211_X1 g720(.A(new_n782), .B(new_n906), .C1(KEYINPUT49), .C2(new_n887), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(KEYINPUT109), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(KEYINPUT109), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT49), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n693), .B1(new_n910), .B2(new_n719), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n909), .A2(new_n892), .A3(new_n911), .ZN(new_n912));
  OAI22_X1  g726(.A1(new_n904), .A2(new_n905), .B1(new_n908), .B2(new_n912), .ZN(G75));
  OAI21_X1  g727(.A(KEYINPUT115), .B1(new_n848), .B2(new_n854), .ZN(new_n914));
  INV_X1    g728(.A(new_n857), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n863), .A2(new_n915), .A3(new_n856), .A4(new_n837), .ZN(new_n916));
  AOI22_X1  g730(.A1(new_n914), .A2(new_n916), .B1(new_n866), .B2(new_n798), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n917), .A2(new_n309), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(G210), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT56), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n320), .B(new_n224), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT55), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n922), .B1(new_n919), .B2(new_n920), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n352), .A2(G952), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT119), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n923), .A2(new_n924), .A3(new_n927), .ZN(G51));
  XNOR2_X1  g742(.A(new_n509), .B(KEYINPUT121), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n914), .A2(new_n916), .ZN(new_n930));
  AOI211_X1 g744(.A(KEYINPUT120), .B(new_n843), .C1(new_n930), .C2(new_n842), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n842), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT54), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT120), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n865), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n931), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n749), .B(KEYINPUT57), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n929), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n774), .A2(G469), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT122), .Z(new_n940));
  NAND2_X1  g754(.A1(new_n918), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n925), .B1(new_n938), .B2(new_n941), .ZN(G54));
  NAND3_X1  g756(.A1(new_n918), .A2(KEYINPUT58), .A3(G475), .ZN(new_n943));
  OAI22_X1  g757(.A1(new_n943), .A2(new_n663), .B1(G952), .B2(new_n352), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n663), .B2(new_n943), .ZN(G60));
  NAND2_X1  g759(.A1(G478), .A2(G902), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT59), .Z(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n948), .B1(new_n870), .B2(new_n903), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n653), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n932), .A2(new_n934), .A3(KEYINPUT54), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT120), .B1(new_n917), .B2(new_n843), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n917), .A2(new_n843), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n653), .A2(new_n947), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n927), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n950), .A2(new_n956), .ZN(G63));
  OAI21_X1  g771(.A(new_n926), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n958));
  NAND2_X1  g772(.A1(G217), .A2(G902), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT123), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT60), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n932), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n958), .B1(new_n962), .B2(new_n616), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n932), .A2(new_n671), .A3(new_n961), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(G66));
  INV_X1    g781(.A(new_n825), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n819), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n352), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n971), .A2(KEYINPUT125), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(KEYINPUT125), .ZN(new_n973));
  OAI21_X1  g787(.A(G953), .B1(new_n372), .B2(new_n221), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n289), .B(new_n291), .C1(G898), .C2(new_n352), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G69));
  XNOR2_X1  g791(.A(new_n535), .B(new_n424), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(new_n493), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n979), .A2(new_n681), .A3(new_n352), .ZN(new_n980));
  INV_X1    g794(.A(new_n796), .ZN(new_n981));
  AND4_X1   g795(.A1(new_n725), .A2(new_n780), .A3(new_n642), .A4(new_n696), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n787), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n835), .A2(new_n742), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n983), .A2(new_n765), .A3(new_n771), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n704), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT62), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n809), .A2(new_n810), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n873), .B1(new_n695), .B2(new_n680), .ZN(new_n989));
  NOR4_X1   g803(.A1(new_n988), .A2(new_n989), .A3(new_n699), .A4(new_n755), .ZN(new_n990));
  NOR4_X1   g804(.A1(new_n787), .A2(new_n981), .A3(new_n987), .A4(new_n990), .ZN(new_n991));
  MUX2_X1   g805(.A(new_n985), .B(new_n991), .S(new_n978), .Z(new_n992));
  AOI21_X1  g806(.A(new_n980), .B1(new_n992), .B2(new_n352), .ZN(G72));
  NAND2_X1  g807(.A1(G472), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT63), .Z(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n985), .B2(new_n969), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n556), .A2(new_n540), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n925), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n991), .A2(new_n819), .A3(new_n968), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n995), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n1000), .A2(new_n540), .A3(new_n556), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n541), .A2(new_n559), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT126), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n995), .B1(new_n1003), .B2(new_n690), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT127), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n867), .A2(new_n868), .A3(new_n1005), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n998), .A2(new_n1001), .A3(new_n1006), .ZN(G57));
endmodule


