

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U554 ( .A(KEYINPUT27), .ZN(n713) );
  XNOR2_X1 U555 ( .A(n714), .B(n713), .ZN(n715) );
  NAND2_X1 U556 ( .A1(n711), .A2(n710), .ZN(n751) );
  OR2_X1 U557 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U558 ( .A1(n533), .A2(G2105), .ZN(n900) );
  XNOR2_X1 U559 ( .A(G543), .B(KEYINPUT0), .ZN(n519) );
  XNOR2_X1 U560 ( .A(n519), .B(KEYINPUT67), .ZN(n635) );
  INV_X1 U561 ( .A(G651), .ZN(n520) );
  NOR2_X1 U562 ( .A1(n635), .A2(n520), .ZN(n642) );
  NAND2_X1 U563 ( .A1(G78), .A2(n642), .ZN(n523) );
  NOR2_X1 U564 ( .A1(G543), .A2(n520), .ZN(n521) );
  XOR2_X1 U565 ( .A(KEYINPUT1), .B(n521), .Z(n651) );
  NAND2_X1 U566 ( .A1(G65), .A2(n651), .ZN(n522) );
  NAND2_X1 U567 ( .A1(n523), .A2(n522), .ZN(n527) );
  NOR2_X1 U568 ( .A1(G651), .A2(G543), .ZN(n645) );
  NAND2_X1 U569 ( .A1(G91), .A2(n645), .ZN(n525) );
  NOR2_X1 U570 ( .A1(G651), .A2(n635), .ZN(n646) );
  NAND2_X1 U571 ( .A1(G53), .A2(n646), .ZN(n524) );
  NAND2_X1 U572 ( .A1(n525), .A2(n524), .ZN(n526) );
  OR2_X1 U573 ( .A1(n527), .A2(n526), .ZN(G299) );
  AND2_X1 U574 ( .A1(G2105), .A2(G2104), .ZN(n901) );
  NAND2_X1 U575 ( .A1(n901), .A2(G113), .ZN(n531) );
  NOR2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  XOR2_X1 U577 ( .A(KEYINPUT66), .B(n528), .Z(n529) );
  XNOR2_X1 U578 ( .A(KEYINPUT17), .B(n529), .ZN(n879) );
  NAND2_X1 U579 ( .A1(G137), .A2(n879), .ZN(n530) );
  AND2_X1 U580 ( .A1(n531), .A2(n530), .ZN(n706) );
  INV_X1 U581 ( .A(G2104), .ZN(n533) );
  NOR2_X1 U582 ( .A1(G2105), .A2(n533), .ZN(n557) );
  NAND2_X1 U583 ( .A1(n557), .A2(G101), .ZN(n532) );
  XOR2_X1 U584 ( .A(n532), .B(KEYINPUT23), .Z(n535) );
  NAND2_X1 U585 ( .A1(n900), .A2(G125), .ZN(n534) );
  NAND2_X1 U586 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U587 ( .A(n536), .B(KEYINPUT65), .ZN(n704) );
  AND2_X1 U588 ( .A1(n706), .A2(n704), .ZN(G160) );
  NAND2_X1 U589 ( .A1(G72), .A2(n642), .ZN(n538) );
  NAND2_X1 U590 ( .A1(G60), .A2(n651), .ZN(n537) );
  NAND2_X1 U591 ( .A1(n538), .A2(n537), .ZN(n542) );
  NAND2_X1 U592 ( .A1(G85), .A2(n645), .ZN(n540) );
  NAND2_X1 U593 ( .A1(G47), .A2(n646), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n540), .A2(n539), .ZN(n541) );
  OR2_X1 U595 ( .A1(n542), .A2(n541), .ZN(G290) );
  XOR2_X1 U596 ( .A(G2446), .B(G2430), .Z(n544) );
  XNOR2_X1 U597 ( .A(G2451), .B(G2454), .ZN(n543) );
  XNOR2_X1 U598 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U599 ( .A(n545), .B(G2427), .Z(n547) );
  XNOR2_X1 U600 ( .A(G1348), .B(G1341), .ZN(n546) );
  XNOR2_X1 U601 ( .A(n547), .B(n546), .ZN(n551) );
  XOR2_X1 U602 ( .A(G2443), .B(KEYINPUT106), .Z(n549) );
  XNOR2_X1 U603 ( .A(G2438), .B(G2435), .ZN(n548) );
  XNOR2_X1 U604 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U605 ( .A(n551), .B(n550), .Z(n552) );
  AND2_X1 U606 ( .A1(G14), .A2(n552), .ZN(G401) );
  AND2_X1 U607 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U608 ( .A1(n900), .A2(G123), .ZN(n554) );
  XNOR2_X1 U609 ( .A(KEYINPUT18), .B(KEYINPUT74), .ZN(n553) );
  XNOR2_X1 U610 ( .A(n554), .B(n553), .ZN(n562) );
  NAND2_X1 U611 ( .A1(n901), .A2(G111), .ZN(n556) );
  BUF_X1 U612 ( .A(n879), .Z(n905) );
  NAND2_X1 U613 ( .A1(G135), .A2(n905), .ZN(n555) );
  NAND2_X1 U614 ( .A1(n556), .A2(n555), .ZN(n560) );
  BUF_X1 U615 ( .A(n557), .Z(n904) );
  NAND2_X1 U616 ( .A1(G99), .A2(n904), .ZN(n558) );
  XNOR2_X1 U617 ( .A(KEYINPUT75), .B(n558), .ZN(n559) );
  NOR2_X1 U618 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U619 ( .A1(n562), .A2(n561), .ZN(n1001) );
  XNOR2_X1 U620 ( .A(G2096), .B(n1001), .ZN(n563) );
  OR2_X1 U621 ( .A1(G2100), .A2(n563), .ZN(G156) );
  INV_X1 U622 ( .A(G57), .ZN(G237) );
  INV_X1 U623 ( .A(G132), .ZN(G219) );
  INV_X1 U624 ( .A(G82), .ZN(G220) );
  NAND2_X1 U625 ( .A1(n651), .A2(G62), .ZN(n564) );
  XOR2_X1 U626 ( .A(KEYINPUT81), .B(n564), .Z(n566) );
  NAND2_X1 U627 ( .A1(n646), .A2(G50), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U629 ( .A(KEYINPUT82), .B(n567), .Z(n571) );
  NAND2_X1 U630 ( .A1(G75), .A2(n642), .ZN(n569) );
  NAND2_X1 U631 ( .A1(G88), .A2(n645), .ZN(n568) );
  AND2_X1 U632 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U633 ( .A1(n571), .A2(n570), .ZN(G303) );
  NAND2_X1 U634 ( .A1(G64), .A2(n651), .ZN(n573) );
  NAND2_X1 U635 ( .A1(G52), .A2(n646), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n573), .A2(n572), .ZN(n578) );
  NAND2_X1 U637 ( .A1(G77), .A2(n642), .ZN(n575) );
  NAND2_X1 U638 ( .A1(G90), .A2(n645), .ZN(n574) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U640 ( .A(KEYINPUT9), .B(n576), .Z(n577) );
  NOR2_X1 U641 ( .A1(n578), .A2(n577), .ZN(G171) );
  INV_X1 U642 ( .A(G171), .ZN(G301) );
  NAND2_X1 U643 ( .A1(G89), .A2(n645), .ZN(n579) );
  XOR2_X1 U644 ( .A(KEYINPUT71), .B(n579), .Z(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(KEYINPUT4), .ZN(n582) );
  NAND2_X1 U646 ( .A1(G76), .A2(n642), .ZN(n581) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(KEYINPUT5), .ZN(n589) );
  NAND2_X1 U649 ( .A1(n651), .A2(G63), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n584), .B(KEYINPUT72), .ZN(n586) );
  NAND2_X1 U651 ( .A1(G51), .A2(n646), .ZN(n585) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U653 ( .A(KEYINPUT6), .B(n587), .Z(n588) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n590), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U656 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U657 ( .A(KEYINPUT68), .B(KEYINPUT11), .Z(n593) );
  NAND2_X1 U658 ( .A1(G7), .A2(G661), .ZN(n591) );
  XOR2_X1 U659 ( .A(n591), .B(KEYINPUT10), .Z(n928) );
  NAND2_X1 U660 ( .A1(G567), .A2(n928), .ZN(n592) );
  XNOR2_X1 U661 ( .A(n593), .B(n592), .ZN(G234) );
  NAND2_X1 U662 ( .A1(G56), .A2(n651), .ZN(n594) );
  XOR2_X1 U663 ( .A(KEYINPUT14), .B(n594), .Z(n602) );
  NAND2_X1 U664 ( .A1(n642), .A2(G68), .ZN(n595) );
  XNOR2_X1 U665 ( .A(KEYINPUT70), .B(n595), .ZN(n599) );
  XOR2_X1 U666 ( .A(KEYINPUT69), .B(KEYINPUT12), .Z(n597) );
  NAND2_X1 U667 ( .A1(G81), .A2(n645), .ZN(n596) );
  XNOR2_X1 U668 ( .A(n597), .B(n596), .ZN(n598) );
  NAND2_X1 U669 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U670 ( .A(KEYINPUT13), .B(n600), .Z(n601) );
  NOR2_X1 U671 ( .A1(n602), .A2(n601), .ZN(n604) );
  NAND2_X1 U672 ( .A1(n646), .A2(G43), .ZN(n603) );
  NAND2_X1 U673 ( .A1(n604), .A2(n603), .ZN(n929) );
  INV_X1 U674 ( .A(G860), .ZN(n624) );
  OR2_X1 U675 ( .A1(n929), .A2(n624), .ZN(G153) );
  NAND2_X1 U676 ( .A1(G868), .A2(G301), .ZN(n613) );
  NAND2_X1 U677 ( .A1(G92), .A2(n645), .ZN(n606) );
  NAND2_X1 U678 ( .A1(G54), .A2(n646), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U680 ( .A1(G79), .A2(n642), .ZN(n608) );
  NAND2_X1 U681 ( .A1(G66), .A2(n651), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U683 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U684 ( .A(n611), .B(KEYINPUT15), .Z(n932) );
  INV_X1 U685 ( .A(n932), .ZN(n728) );
  INV_X1 U686 ( .A(G868), .ZN(n618) );
  NAND2_X1 U687 ( .A1(n728), .A2(n618), .ZN(n612) );
  NAND2_X1 U688 ( .A1(n613), .A2(n612), .ZN(G284) );
  NOR2_X1 U689 ( .A1(G868), .A2(G299), .ZN(n615) );
  NOR2_X1 U690 ( .A1(G286), .A2(n618), .ZN(n614) );
  NOR2_X1 U691 ( .A1(n615), .A2(n614), .ZN(G297) );
  NAND2_X1 U692 ( .A1(n624), .A2(G559), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n616), .A2(n932), .ZN(n617) );
  XNOR2_X1 U694 ( .A(n617), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U695 ( .A1(n728), .A2(n618), .ZN(n619) );
  XNOR2_X1 U696 ( .A(n619), .B(KEYINPUT73), .ZN(n620) );
  NOR2_X1 U697 ( .A1(G559), .A2(n620), .ZN(n622) );
  NOR2_X1 U698 ( .A1(G868), .A2(n929), .ZN(n621) );
  NOR2_X1 U699 ( .A1(n622), .A2(n621), .ZN(G282) );
  NAND2_X1 U700 ( .A1(G559), .A2(n932), .ZN(n623) );
  XOR2_X1 U701 ( .A(n929), .B(n623), .Z(n660) );
  NAND2_X1 U702 ( .A1(n624), .A2(n660), .ZN(n633) );
  NAND2_X1 U703 ( .A1(G80), .A2(n642), .ZN(n626) );
  NAND2_X1 U704 ( .A1(G93), .A2(n645), .ZN(n625) );
  NAND2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U706 ( .A(KEYINPUT76), .B(n627), .Z(n629) );
  NAND2_X1 U707 ( .A1(n646), .A2(G55), .ZN(n628) );
  NAND2_X1 U708 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U709 ( .A1(G67), .A2(n651), .ZN(n630) );
  XNOR2_X1 U710 ( .A(KEYINPUT77), .B(n630), .ZN(n631) );
  NOR2_X1 U711 ( .A1(n632), .A2(n631), .ZN(n662) );
  XOR2_X1 U712 ( .A(n633), .B(n662), .Z(G145) );
  NAND2_X1 U713 ( .A1(G49), .A2(n646), .ZN(n634) );
  XNOR2_X1 U714 ( .A(n634), .B(KEYINPUT78), .ZN(n640) );
  NAND2_X1 U715 ( .A1(G87), .A2(n635), .ZN(n637) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U718 ( .A1(n651), .A2(n638), .ZN(n639) );
  NAND2_X1 U719 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U720 ( .A(KEYINPUT79), .B(n641), .Z(G288) );
  XOR2_X1 U721 ( .A(KEYINPUT80), .B(KEYINPUT2), .Z(n644) );
  NAND2_X1 U722 ( .A1(G73), .A2(n642), .ZN(n643) );
  XNOR2_X1 U723 ( .A(n644), .B(n643), .ZN(n650) );
  NAND2_X1 U724 ( .A1(G86), .A2(n645), .ZN(n648) );
  NAND2_X1 U725 ( .A1(G48), .A2(n646), .ZN(n647) );
  NAND2_X1 U726 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U727 ( .A1(n650), .A2(n649), .ZN(n653) );
  NAND2_X1 U728 ( .A1(n651), .A2(G61), .ZN(n652) );
  NAND2_X1 U729 ( .A1(n653), .A2(n652), .ZN(G305) );
  XOR2_X1 U730 ( .A(G303), .B(G288), .Z(n659) );
  XNOR2_X1 U731 ( .A(KEYINPUT19), .B(n662), .ZN(n655) );
  XNOR2_X1 U732 ( .A(G290), .B(KEYINPUT83), .ZN(n654) );
  XNOR2_X1 U733 ( .A(n655), .B(n654), .ZN(n656) );
  XOR2_X1 U734 ( .A(n656), .B(G305), .Z(n657) );
  XNOR2_X1 U735 ( .A(G299), .B(n657), .ZN(n658) );
  XNOR2_X1 U736 ( .A(n659), .B(n658), .ZN(n848) );
  XNOR2_X1 U737 ( .A(n660), .B(n848), .ZN(n661) );
  NAND2_X1 U738 ( .A1(n661), .A2(G868), .ZN(n664) );
  OR2_X1 U739 ( .A1(G868), .A2(n662), .ZN(n663) );
  NAND2_X1 U740 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2078), .A2(G2084), .ZN(n665) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n666), .ZN(n667) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n667), .ZN(n668) );
  NAND2_X1 U745 ( .A1(n668), .A2(G2072), .ZN(n669) );
  XNOR2_X1 U746 ( .A(KEYINPUT84), .B(n669), .ZN(G158) );
  XNOR2_X1 U747 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U748 ( .A1(G220), .A2(G219), .ZN(n670) );
  XNOR2_X1 U749 ( .A(KEYINPUT22), .B(n670), .ZN(n671) );
  NAND2_X1 U750 ( .A1(n671), .A2(G96), .ZN(n672) );
  NOR2_X1 U751 ( .A1(n672), .A2(G218), .ZN(n673) );
  XNOR2_X1 U752 ( .A(n673), .B(KEYINPUT85), .ZN(n925) );
  NAND2_X1 U753 ( .A1(G2106), .A2(n925), .ZN(n674) );
  XNOR2_X1 U754 ( .A(KEYINPUT86), .B(n674), .ZN(n678) );
  NAND2_X1 U755 ( .A1(G120), .A2(G69), .ZN(n675) );
  NOR2_X1 U756 ( .A1(G237), .A2(n675), .ZN(n676) );
  NAND2_X1 U757 ( .A1(G108), .A2(n676), .ZN(n926) );
  NAND2_X1 U758 ( .A1(G567), .A2(n926), .ZN(n677) );
  NAND2_X1 U759 ( .A1(n678), .A2(n677), .ZN(n927) );
  NAND2_X1 U760 ( .A1(G661), .A2(G483), .ZN(n679) );
  NOR2_X1 U761 ( .A1(n927), .A2(n679), .ZN(n845) );
  NAND2_X1 U762 ( .A1(n845), .A2(G36), .ZN(G176) );
  NAND2_X1 U763 ( .A1(n904), .A2(G102), .ZN(n681) );
  NAND2_X1 U764 ( .A1(G138), .A2(n879), .ZN(n680) );
  NAND2_X1 U765 ( .A1(n681), .A2(n680), .ZN(n685) );
  NAND2_X1 U766 ( .A1(G126), .A2(n900), .ZN(n683) );
  NAND2_X1 U767 ( .A1(G114), .A2(n901), .ZN(n682) );
  NAND2_X1 U768 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U769 ( .A1(n685), .A2(n684), .ZN(G164) );
  NAND2_X1 U770 ( .A1(n904), .A2(G95), .ZN(n687) );
  NAND2_X1 U771 ( .A1(G131), .A2(n905), .ZN(n686) );
  NAND2_X1 U772 ( .A1(n687), .A2(n686), .ZN(n691) );
  NAND2_X1 U773 ( .A1(G119), .A2(n900), .ZN(n689) );
  NAND2_X1 U774 ( .A1(G107), .A2(n901), .ZN(n688) );
  NAND2_X1 U775 ( .A1(n689), .A2(n688), .ZN(n690) );
  OR2_X1 U776 ( .A1(n691), .A2(n690), .ZN(n892) );
  AND2_X1 U777 ( .A1(n892), .A2(G1991), .ZN(n703) );
  NAND2_X1 U778 ( .A1(n905), .A2(G141), .ZN(n692) );
  XNOR2_X1 U779 ( .A(n692), .B(KEYINPUT92), .ZN(n701) );
  NAND2_X1 U780 ( .A1(G105), .A2(n904), .ZN(n693) );
  XOR2_X1 U781 ( .A(KEYINPUT38), .B(n693), .Z(n694) );
  XNOR2_X1 U782 ( .A(n694), .B(KEYINPUT91), .ZN(n696) );
  NAND2_X1 U783 ( .A1(G129), .A2(n900), .ZN(n695) );
  NAND2_X1 U784 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U785 ( .A1(n901), .A2(G117), .ZN(n697) );
  XOR2_X1 U786 ( .A(KEYINPUT90), .B(n697), .Z(n698) );
  NOR2_X1 U787 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U788 ( .A1(n701), .A2(n700), .ZN(n915) );
  AND2_X1 U789 ( .A1(n915), .A2(G1996), .ZN(n702) );
  NOR2_X1 U790 ( .A1(n703), .A2(n702), .ZN(n1006) );
  NOR2_X1 U791 ( .A1(G164), .A2(G1384), .ZN(n710) );
  AND2_X1 U792 ( .A1(G40), .A2(n704), .ZN(n705) );
  NAND2_X1 U793 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U794 ( .A(n707), .B(KEYINPUT88), .ZN(n709) );
  NOR2_X1 U795 ( .A1(n710), .A2(n709), .ZN(n837) );
  INV_X1 U796 ( .A(n837), .ZN(n708) );
  NOR2_X1 U797 ( .A1(n1006), .A2(n708), .ZN(n828) );
  XNOR2_X1 U798 ( .A(KEYINPUT93), .B(n709), .ZN(n711) );
  XNOR2_X1 U799 ( .A(KEYINPUT95), .B(n751), .ZN(n712) );
  BUF_X1 U800 ( .A(n712), .Z(n718) );
  INV_X1 U801 ( .A(n718), .ZN(n741) );
  XNOR2_X1 U802 ( .A(G1956), .B(KEYINPUT96), .ZN(n967) );
  NAND2_X1 U803 ( .A1(n741), .A2(n967), .ZN(n716) );
  NAND2_X1 U804 ( .A1(n712), .A2(G2072), .ZN(n714) );
  NAND2_X1 U805 ( .A1(n716), .A2(n715), .ZN(n734) );
  NOR2_X1 U806 ( .A1(G299), .A2(n734), .ZN(n717) );
  XOR2_X1 U807 ( .A(KEYINPUT97), .B(n717), .Z(n722) );
  NAND2_X1 U808 ( .A1(G2067), .A2(n718), .ZN(n720) );
  NAND2_X1 U809 ( .A1(G1348), .A2(n751), .ZN(n719) );
  NAND2_X1 U810 ( .A1(n720), .A2(n719), .ZN(n729) );
  NOR2_X1 U811 ( .A1(n728), .A2(n729), .ZN(n721) );
  NOR2_X1 U812 ( .A1(n722), .A2(n721), .ZN(n733) );
  INV_X1 U813 ( .A(G1996), .ZN(n868) );
  NOR2_X1 U814 ( .A1(n751), .A2(n868), .ZN(n723) );
  XOR2_X1 U815 ( .A(n723), .B(KEYINPUT26), .Z(n725) );
  NAND2_X1 U816 ( .A1(n751), .A2(G1341), .ZN(n724) );
  NAND2_X1 U817 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U818 ( .A1(n929), .A2(n726), .ZN(n727) );
  XNOR2_X1 U819 ( .A(n727), .B(KEYINPUT64), .ZN(n731) );
  NAND2_X1 U820 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U821 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U822 ( .A1(n733), .A2(n732), .ZN(n737) );
  NAND2_X1 U823 ( .A1(G299), .A2(n734), .ZN(n735) );
  XNOR2_X1 U824 ( .A(n735), .B(KEYINPUT28), .ZN(n736) );
  NAND2_X1 U825 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U826 ( .A(n738), .B(KEYINPUT29), .ZN(n767) );
  INV_X1 U827 ( .A(n751), .ZN(n739) );
  NOR2_X1 U828 ( .A1(n739), .A2(G1961), .ZN(n740) );
  XNOR2_X1 U829 ( .A(n740), .B(KEYINPUT94), .ZN(n743) );
  XOR2_X1 U830 ( .A(KEYINPUT25), .B(G2078), .Z(n979) );
  NOR2_X1 U831 ( .A1(n741), .A2(n979), .ZN(n742) );
  NOR2_X1 U832 ( .A1(n743), .A2(n742), .ZN(n755) );
  NOR2_X1 U833 ( .A1(G301), .A2(n755), .ZN(n766) );
  INV_X1 U834 ( .A(G8), .ZN(n748) );
  NAND2_X1 U835 ( .A1(G8), .A2(n751), .ZN(n800) );
  NOR2_X1 U836 ( .A1(G1971), .A2(n800), .ZN(n745) );
  NOR2_X1 U837 ( .A1(G2090), .A2(n751), .ZN(n744) );
  NOR2_X1 U838 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U839 ( .A1(n746), .A2(G303), .ZN(n747) );
  NOR2_X1 U840 ( .A1(n748), .A2(n747), .ZN(n759) );
  OR2_X1 U841 ( .A1(n759), .A2(G286), .ZN(n761) );
  INV_X1 U842 ( .A(n761), .ZN(n749) );
  OR2_X1 U843 ( .A1(n766), .A2(n749), .ZN(n750) );
  NOR2_X1 U844 ( .A1(n767), .A2(n750), .ZN(n763) );
  NOR2_X1 U845 ( .A1(G1966), .A2(n800), .ZN(n771) );
  NOR2_X1 U846 ( .A1(G2084), .A2(n751), .ZN(n770) );
  NOR2_X1 U847 ( .A1(n771), .A2(n770), .ZN(n752) );
  NAND2_X1 U848 ( .A1(G8), .A2(n752), .ZN(n753) );
  XNOR2_X1 U849 ( .A(KEYINPUT30), .B(n753), .ZN(n754) );
  NOR2_X1 U850 ( .A1(G168), .A2(n754), .ZN(n757) );
  AND2_X1 U851 ( .A1(G301), .A2(n755), .ZN(n756) );
  NOR2_X1 U852 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U853 ( .A(n758), .B(KEYINPUT31), .ZN(n768) );
  OR2_X1 U854 ( .A1(n768), .A2(n759), .ZN(n760) );
  AND2_X1 U855 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U856 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U857 ( .A(n764), .B(KEYINPUT32), .ZN(n765) );
  XNOR2_X1 U858 ( .A(n765), .B(KEYINPUT98), .ZN(n794) );
  NOR2_X1 U859 ( .A1(n767), .A2(n766), .ZN(n769) );
  OR2_X1 U860 ( .A1(n769), .A2(n768), .ZN(n774) );
  AND2_X1 U861 ( .A1(n770), .A2(G8), .ZN(n772) );
  NOR2_X1 U862 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U863 ( .A1(n774), .A2(n773), .ZN(n787) );
  AND2_X1 U864 ( .A1(n787), .A2(n800), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n794), .A2(n775), .ZN(n779) );
  INV_X1 U866 ( .A(n800), .ZN(n788) );
  NOR2_X1 U867 ( .A1(G2090), .A2(G303), .ZN(n776) );
  NAND2_X1 U868 ( .A1(G8), .A2(n776), .ZN(n777) );
  OR2_X1 U869 ( .A1(n788), .A2(n777), .ZN(n778) );
  NAND2_X1 U870 ( .A1(n779), .A2(n778), .ZN(n781) );
  INV_X1 U871 ( .A(KEYINPUT102), .ZN(n780) );
  XNOR2_X1 U872 ( .A(n781), .B(n780), .ZN(n785) );
  NOR2_X1 U873 ( .A1(G1981), .A2(G305), .ZN(n782) );
  XOR2_X1 U874 ( .A(n782), .B(KEYINPUT24), .Z(n783) );
  OR2_X1 U875 ( .A1(n800), .A2(n783), .ZN(n784) );
  AND2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n809) );
  NAND2_X1 U877 ( .A1(G288), .A2(G1976), .ZN(n786) );
  XOR2_X1 U878 ( .A(KEYINPUT101), .B(n786), .Z(n947) );
  AND2_X1 U879 ( .A1(n787), .A2(n947), .ZN(n789) );
  AND2_X1 U880 ( .A1(n789), .A2(n788), .ZN(n792) );
  NOR2_X1 U881 ( .A1(G1976), .A2(G288), .ZN(n790) );
  XOR2_X1 U882 ( .A(KEYINPUT99), .B(n790), .Z(n796) );
  NAND2_X1 U883 ( .A1(n796), .A2(KEYINPUT33), .ZN(n791) );
  OR2_X1 U884 ( .A1(n800), .A2(n791), .ZN(n804) );
  AND2_X1 U885 ( .A1(n792), .A2(n804), .ZN(n793) );
  AND2_X1 U886 ( .A1(n794), .A2(n793), .ZN(n806) );
  INV_X1 U887 ( .A(n947), .ZN(n798) );
  NOR2_X1 U888 ( .A1(G1971), .A2(G303), .ZN(n795) );
  NOR2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n940) );
  XNOR2_X1 U890 ( .A(KEYINPUT100), .B(n940), .ZN(n797) );
  OR2_X1 U891 ( .A1(n798), .A2(n797), .ZN(n799) );
  OR2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n802) );
  INV_X1 U893 ( .A(KEYINPUT33), .ZN(n801) );
  NAND2_X1 U894 ( .A1(n802), .A2(n801), .ZN(n803) );
  AND2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U896 ( .A(G1981), .B(G305), .Z(n943) );
  NAND2_X1 U897 ( .A1(n807), .A2(n943), .ZN(n808) );
  AND2_X1 U898 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U899 ( .A1(n828), .A2(n810), .ZN(n825) );
  XNOR2_X1 U900 ( .A(KEYINPUT87), .B(G1986), .ZN(n811) );
  XNOR2_X1 U901 ( .A(n811), .B(G290), .ZN(n936) );
  XNOR2_X1 U902 ( .A(G2067), .B(KEYINPUT37), .ZN(n835) );
  NAND2_X1 U903 ( .A1(n900), .A2(G128), .ZN(n812) );
  XOR2_X1 U904 ( .A(KEYINPUT89), .B(n812), .Z(n814) );
  NAND2_X1 U905 ( .A1(n901), .A2(G116), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U907 ( .A(n815), .B(KEYINPUT35), .ZN(n820) );
  NAND2_X1 U908 ( .A1(n904), .A2(G104), .ZN(n817) );
  NAND2_X1 U909 ( .A1(G140), .A2(n879), .ZN(n816) );
  NAND2_X1 U910 ( .A1(n817), .A2(n816), .ZN(n818) );
  XOR2_X1 U911 ( .A(KEYINPUT34), .B(n818), .Z(n819) );
  NAND2_X1 U912 ( .A1(n820), .A2(n819), .ZN(n821) );
  XOR2_X1 U913 ( .A(n821), .B(KEYINPUT36), .Z(n914) );
  NOR2_X1 U914 ( .A1(n835), .A2(n914), .ZN(n1015) );
  INV_X1 U915 ( .A(n1015), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n936), .A2(n822), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n823), .A2(n837), .ZN(n824) );
  NAND2_X1 U918 ( .A1(n825), .A2(n824), .ZN(n840) );
  NOR2_X1 U919 ( .A1(G1996), .A2(n915), .ZN(n1012) );
  NOR2_X1 U920 ( .A1(G1986), .A2(G290), .ZN(n826) );
  NOR2_X1 U921 ( .A1(G1991), .A2(n892), .ZN(n1004) );
  NOR2_X1 U922 ( .A1(n826), .A2(n1004), .ZN(n827) );
  NOR2_X1 U923 ( .A1(n828), .A2(n827), .ZN(n829) );
  XOR2_X1 U924 ( .A(KEYINPUT103), .B(n829), .Z(n830) );
  NOR2_X1 U925 ( .A1(n1012), .A2(n830), .ZN(n831) );
  XOR2_X1 U926 ( .A(KEYINPUT104), .B(n831), .Z(n832) );
  XNOR2_X1 U927 ( .A(n832), .B(KEYINPUT39), .ZN(n833) );
  NOR2_X1 U928 ( .A1(n1015), .A2(n833), .ZN(n834) );
  XNOR2_X1 U929 ( .A(n834), .B(KEYINPUT105), .ZN(n836) );
  NAND2_X1 U930 ( .A1(n835), .A2(n914), .ZN(n1021) );
  NAND2_X1 U931 ( .A1(n836), .A2(n1021), .ZN(n838) );
  NAND2_X1 U932 ( .A1(n838), .A2(n837), .ZN(n839) );
  NAND2_X1 U933 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U934 ( .A(KEYINPUT40), .B(n841), .ZN(G329) );
  NAND2_X1 U935 ( .A1(G2106), .A2(n928), .ZN(G217) );
  AND2_X1 U936 ( .A1(G15), .A2(G2), .ZN(n842) );
  NAND2_X1 U937 ( .A1(G661), .A2(n842), .ZN(G259) );
  NAND2_X1 U938 ( .A1(G3), .A2(G1), .ZN(n843) );
  XOR2_X1 U939 ( .A(KEYINPUT107), .B(n843), .Z(n844) );
  NAND2_X1 U940 ( .A1(n845), .A2(n844), .ZN(G188) );
  XOR2_X1 U941 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  XOR2_X1 U942 ( .A(n932), .B(KEYINPUT118), .Z(n847) );
  XOR2_X1 U943 ( .A(G286), .B(G301), .Z(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n850) );
  XOR2_X1 U945 ( .A(n929), .B(n848), .Z(n849) );
  XNOR2_X1 U946 ( .A(n850), .B(n849), .ZN(n851) );
  NOR2_X1 U947 ( .A1(G37), .A2(n851), .ZN(G397) );
  XOR2_X1 U948 ( .A(KEYINPUT42), .B(G2084), .Z(n853) );
  XNOR2_X1 U949 ( .A(G2090), .B(G2072), .ZN(n852) );
  XNOR2_X1 U950 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U951 ( .A(n854), .B(G2100), .Z(n856) );
  XNOR2_X1 U952 ( .A(G2078), .B(G2067), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U954 ( .A(G2096), .B(KEYINPUT43), .Z(n858) );
  XNOR2_X1 U955 ( .A(KEYINPUT109), .B(G2678), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U957 ( .A(n860), .B(n859), .Z(G227) );
  XOR2_X1 U958 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n862) );
  XNOR2_X1 U959 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U961 ( .A(n863), .B(G2474), .Z(n865) );
  XNOR2_X1 U962 ( .A(G1981), .B(G1986), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n865), .B(n864), .ZN(n874) );
  XOR2_X1 U964 ( .A(G1966), .B(G1961), .Z(n867) );
  XNOR2_X1 U965 ( .A(G1976), .B(G1971), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(n872) );
  XOR2_X1 U967 ( .A(KEYINPUT112), .B(G1991), .Z(n870) );
  XOR2_X1 U968 ( .A(n868), .B(G1956), .Z(n869) );
  XNOR2_X1 U969 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U970 ( .A(n872), .B(n871), .Z(n873) );
  XNOR2_X1 U971 ( .A(n874), .B(n873), .ZN(G229) );
  NAND2_X1 U972 ( .A1(G124), .A2(n900), .ZN(n875) );
  XNOR2_X1 U973 ( .A(n875), .B(KEYINPUT44), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n876), .B(KEYINPUT114), .ZN(n878) );
  NAND2_X1 U975 ( .A1(G112), .A2(n901), .ZN(n877) );
  NAND2_X1 U976 ( .A1(n878), .A2(n877), .ZN(n883) );
  NAND2_X1 U977 ( .A1(n904), .A2(G100), .ZN(n881) );
  NAND2_X1 U978 ( .A1(G136), .A2(n879), .ZN(n880) );
  NAND2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n882) );
  NOR2_X1 U980 ( .A1(n883), .A2(n882), .ZN(G162) );
  NAND2_X1 U981 ( .A1(G127), .A2(n900), .ZN(n885) );
  NAND2_X1 U982 ( .A1(G115), .A2(n901), .ZN(n884) );
  NAND2_X1 U983 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U984 ( .A(n886), .B(KEYINPUT47), .ZN(n888) );
  NAND2_X1 U985 ( .A1(G103), .A2(n904), .ZN(n887) );
  NAND2_X1 U986 ( .A1(n888), .A2(n887), .ZN(n891) );
  NAND2_X1 U987 ( .A1(G139), .A2(n905), .ZN(n889) );
  XNOR2_X1 U988 ( .A(KEYINPUT115), .B(n889), .ZN(n890) );
  NOR2_X1 U989 ( .A1(n891), .A2(n890), .ZN(n1007) );
  XOR2_X1 U990 ( .A(n892), .B(n1007), .Z(n896) );
  XOR2_X1 U991 ( .A(KEYINPUT46), .B(KEYINPUT116), .Z(n894) );
  XNOR2_X1 U992 ( .A(KEYINPUT117), .B(KEYINPUT48), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U995 ( .A(G162), .B(n897), .Z(n899) );
  XNOR2_X1 U996 ( .A(G164), .B(G160), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n913) );
  NAND2_X1 U998 ( .A1(G130), .A2(n900), .ZN(n903) );
  NAND2_X1 U999 ( .A1(G118), .A2(n901), .ZN(n902) );
  NAND2_X1 U1000 ( .A1(n903), .A2(n902), .ZN(n910) );
  NAND2_X1 U1001 ( .A1(n904), .A2(G106), .ZN(n907) );
  NAND2_X1 U1002 ( .A1(G142), .A2(n905), .ZN(n906) );
  NAND2_X1 U1003 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1004 ( .A(n908), .B(KEYINPUT45), .Z(n909) );
  NOR2_X1 U1005 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(n911), .B(n1001), .ZN(n912) );
  XOR2_X1 U1007 ( .A(n913), .B(n912), .Z(n917) );
  XNOR2_X1 U1008 ( .A(n915), .B(n914), .ZN(n916) );
  XNOR2_X1 U1009 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n918), .ZN(G395) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n919) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n919), .ZN(n920) );
  NOR2_X1 U1013 ( .A1(G397), .A2(n920), .ZN(n924) );
  NOR2_X1 U1014 ( .A1(G401), .A2(n927), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(KEYINPUT119), .B(n921), .ZN(n922) );
  NOR2_X1 U1016 ( .A1(G395), .A2(n922), .ZN(n923) );
  NAND2_X1 U1017 ( .A1(n924), .A2(n923), .ZN(G225) );
  XOR2_X1 U1018 ( .A(KEYINPUT120), .B(G225), .Z(G308) );
  INV_X1 U1020 ( .A(G120), .ZN(G236) );
  INV_X1 U1021 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(G325) );
  INV_X1 U1023 ( .A(G325), .ZN(G261) );
  INV_X1 U1024 ( .A(n927), .ZN(G319) );
  INV_X1 U1025 ( .A(G108), .ZN(G238) );
  INV_X1 U1026 ( .A(n928), .ZN(G223) );
  XOR2_X1 U1027 ( .A(G16), .B(KEYINPUT56), .Z(n952) );
  XNOR2_X1 U1028 ( .A(G1341), .B(n929), .ZN(n950) );
  XOR2_X1 U1029 ( .A(G1956), .B(G299), .Z(n931) );
  NAND2_X1 U1030 ( .A1(G1971), .A2(G303), .ZN(n930) );
  NAND2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n938) );
  XOR2_X1 U1032 ( .A(G171), .B(G1961), .Z(n934) );
  XOR2_X1 U1033 ( .A(n932), .B(G1348), .Z(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n946) );
  XNOR2_X1 U1038 ( .A(G168), .B(G1966), .ZN(n941) );
  XNOR2_X1 U1039 ( .A(n941), .B(KEYINPUT124), .ZN(n942) );
  NAND2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1041 ( .A(KEYINPUT57), .B(n944), .Z(n945) );
  NOR2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n948) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n1030) );
  XNOR2_X1 U1046 ( .A(G1976), .B(G23), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(G22), .B(G1971), .ZN(n953) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1049 ( .A(KEYINPUT126), .B(n955), .Z(n957) );
  XNOR2_X1 U1050 ( .A(G1986), .B(G24), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(KEYINPUT58), .B(n958), .ZN(n962) );
  XNOR2_X1 U1053 ( .A(G1961), .B(G5), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(G1966), .B(G21), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n974) );
  XNOR2_X1 U1057 ( .A(G1981), .B(G6), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(KEYINPUT59), .B(G4), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(n963), .B(KEYINPUT125), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(n964), .B(G1348), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(n967), .B(G20), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(G19), .B(G1341), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(KEYINPUT60), .B(n972), .ZN(n973) );
  NOR2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1068 ( .A(KEYINPUT61), .B(n975), .Z(n976) );
  NOR2_X1 U1069 ( .A1(G16), .A2(n976), .ZN(n1000) );
  XOR2_X1 U1070 ( .A(KEYINPUT123), .B(KEYINPUT53), .Z(n989) );
  XOR2_X1 U1071 ( .A(G2067), .B(G26), .Z(n978) );
  XOR2_X1 U1072 ( .A(G1996), .B(G32), .Z(n977) );
  NAND2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(G27), .B(n979), .ZN(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n987) );
  XOR2_X1 U1076 ( .A(G25), .B(G1991), .Z(n982) );
  NAND2_X1 U1077 ( .A1(n982), .A2(G28), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(KEYINPUT122), .B(G2072), .ZN(n983) );
  XNOR2_X1 U1079 ( .A(G33), .B(n983), .ZN(n984) );
  NOR2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(n989), .B(n988), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(G2084), .B(G34), .ZN(n990) );
  XNOR2_X1 U1084 ( .A(n990), .B(KEYINPUT54), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(G35), .B(G2090), .ZN(n991) );
  NOR2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1088 ( .A(KEYINPUT55), .B(n995), .Z(n997) );
  INV_X1 U1089 ( .A(G29), .ZN(n996) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1091 ( .A1(G11), .A2(n998), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1028) );
  XNOR2_X1 U1093 ( .A(G160), .B(G2084), .ZN(n1002) );
  NAND2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1019) );
  XOR2_X1 U1097 ( .A(G2072), .B(n1007), .Z(n1009) );
  XOR2_X1 U1098 ( .A(G164), .B(G2078), .Z(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(KEYINPUT50), .B(n1010), .ZN(n1017) );
  XOR2_X1 U1101 ( .A(G2090), .B(G162), .Z(n1011) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(n1013), .B(KEYINPUT51), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(n1022), .B(KEYINPUT52), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(KEYINPUT121), .B(n1023), .ZN(n1025) );
  INV_X1 U1110 ( .A(KEYINPUT55), .ZN(n1024) );
  NAND2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(G29), .ZN(n1027) );
  NAND2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1115 ( .A(KEYINPUT127), .B(n1031), .Z(n1032) );
  XOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1032), .Z(G150) );
  INV_X1 U1117 ( .A(G150), .ZN(G311) );
  INV_X1 U1118 ( .A(G303), .ZN(G166) );
endmodule

