//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n202), .A2(G77), .A3(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n208));
  INV_X1    g0008(.A(G50), .ZN(new_n209));
  INV_X1    g0009(.A(G226), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n207), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT1), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n207), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT0), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n204), .A2(G50), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(new_n220), .A2(new_n221), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n227), .B1(new_n221), .B2(new_n220), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n218), .A2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT65), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n233), .B(new_n237), .Z(G358));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(G107), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G97), .ZN(new_n243));
  INV_X1    g0043(.A(G97), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G107), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n241), .B(new_n248), .Z(G351));
  INV_X1    g0049(.A(KEYINPUT11), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G50), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT77), .ZN(new_n253));
  INV_X1    g0053(.A(G68), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n252), .A2(new_n253), .B1(G20), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n251), .A2(KEYINPUT77), .A3(G50), .ZN(new_n256));
  INV_X1    g0056(.A(G77), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT68), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n258), .B1(new_n259), .B2(G20), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n225), .A2(KEYINPUT68), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n255), .B(new_n256), .C1(new_n257), .C2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT78), .ZN(new_n264));
  NAND3_X1  g0064(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n224), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n263), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n264), .B1(new_n263), .B2(new_n266), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n250), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n269), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(KEYINPUT11), .A3(new_n267), .ZN(new_n272));
  INV_X1    g0072(.A(G1), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G13), .A3(G20), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G68), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT12), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n265), .A2(new_n224), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(new_n274), .A3(KEYINPUT72), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT72), .ZN(new_n279));
  INV_X1    g0079(.A(new_n274), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n279), .B1(new_n280), .B2(new_n266), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n273), .A2(G20), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n276), .B1(new_n284), .B2(G68), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n270), .A2(new_n272), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G200), .ZN(new_n287));
  OR2_X1    g0087(.A1(KEYINPUT66), .A2(G45), .ZN(new_n288));
  NAND2_X1  g0088(.A1(KEYINPUT66), .A2(G45), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G41), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT74), .ZN(new_n293));
  INV_X1    g0093(.A(G274), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G1), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n292), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(G41), .B1(new_n288), .B2(new_n289), .ZN(new_n297));
  INV_X1    g0097(.A(new_n295), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT74), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G41), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n300), .A2(G1), .A3(G13), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n273), .B1(G41), .B2(G45), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n296), .A2(new_n299), .B1(G238), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT3), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G33), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n306), .A2(new_n308), .A3(G232), .A4(G1698), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G97), .ZN(new_n310));
  AND2_X1   g0110(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n311));
  NOR2_X1   g0111(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n306), .B(new_n308), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n309), .B(new_n310), .C1(new_n313), .C2(new_n210), .ZN(new_n314));
  INV_X1    g0114(.A(new_n301), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n305), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT13), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT13), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n305), .A2(new_n319), .A3(new_n316), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n287), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n286), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G190), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT75), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n318), .A2(new_n324), .A3(new_n320), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n317), .A2(KEYINPUT75), .A3(KEYINPUT13), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n323), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT76), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n322), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n327), .A2(new_n328), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n305), .A2(new_n319), .A3(new_n316), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n319), .B1(new_n305), .B2(new_n316), .ZN(new_n333));
  OAI21_X1  g0133(.A(G169), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT14), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT14), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n336), .B(G169), .C1(new_n332), .C2(new_n333), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G179), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n339), .B1(new_n325), .B2(new_n326), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n286), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n331), .A2(new_n341), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n297), .A2(new_n298), .B1(new_n303), .B2(new_n210), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n306), .A2(new_n308), .A3(G1698), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n306), .A2(new_n308), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n344), .A2(G223), .B1(G77), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G222), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n346), .B1(new_n347), .B2(new_n313), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n343), .B1(new_n348), .B2(new_n315), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n349), .A2(G169), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n350), .B1(new_n339), .B2(new_n349), .ZN(new_n351));
  OR2_X1    g0151(.A1(KEYINPUT8), .A2(G58), .ZN(new_n352));
  NAND2_X1  g0152(.A1(KEYINPUT8), .A2(G58), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n260), .A2(new_n261), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n251), .A2(G150), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT69), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n225), .B1(new_n201), .B2(new_n203), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n354), .A2(KEYINPUT69), .A3(new_n355), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n277), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n277), .A2(new_n274), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT70), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n277), .A2(new_n274), .A3(KEYINPUT70), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n363), .A2(G50), .A3(new_n283), .A4(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n280), .A2(new_n209), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n351), .B1(new_n360), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n349), .A2(G190), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n287), .B2(new_n349), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n365), .A2(new_n366), .ZN(new_n371));
  INV_X1    g0171(.A(new_n359), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n372), .A2(new_n357), .A3(new_n356), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n371), .B(KEYINPUT73), .C1(new_n277), .C2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT73), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n360), .B2(new_n367), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n370), .B1(new_n377), .B2(KEYINPUT9), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT10), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT9), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n374), .A2(new_n380), .A3(new_n376), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n378), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n379), .B1(new_n378), .B2(new_n381), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n368), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n344), .A2(G238), .B1(G107), .B2(new_n345), .ZN(new_n385));
  INV_X1    g0185(.A(G232), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n385), .B1(new_n386), .B2(new_n313), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n315), .ZN(new_n388));
  AOI22_X1  g0188(.A1(G244), .A2(new_n304), .B1(new_n292), .B2(new_n295), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n339), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n352), .A2(new_n353), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n393), .A2(new_n251), .B1(G20), .B2(G77), .ZN(new_n394));
  XNOR2_X1  g0194(.A(KEYINPUT15), .B(G87), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n395), .B(KEYINPUT71), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n394), .B1(new_n396), .B2(new_n262), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(new_n266), .B1(new_n257), .B2(new_n280), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n284), .A2(G77), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G169), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n390), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n392), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n390), .A2(G200), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n400), .B1(new_n391), .B2(G190), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT79), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n301), .A2(G232), .A3(new_n302), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n297), .B2(new_n298), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n306), .A2(new_n308), .A3(G226), .A4(G1698), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G87), .ZN(new_n412));
  INV_X1    g0212(.A(G223), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n411), .B(new_n412), .C1(new_n313), .C2(new_n413), .ZN(new_n414));
  AOI211_X1 g0214(.A(G190), .B(new_n410), .C1(new_n315), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n315), .ZN(new_n416));
  INV_X1    g0216(.A(new_n410), .ZN(new_n417));
  AOI21_X1  g0217(.A(G200), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n408), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n410), .B1(new_n414), .B2(new_n315), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n323), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n421), .B(KEYINPUT79), .C1(G200), .C2(new_n420), .ZN(new_n422));
  XNOR2_X1  g0222(.A(KEYINPUT3), .B(G33), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT7), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n423), .A2(new_n424), .A3(G20), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT7), .B1(new_n345), .B2(new_n225), .ZN(new_n426));
  OAI21_X1  g0226(.A(G68), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(G58), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(new_n254), .ZN(new_n429));
  OAI21_X1  g0229(.A(G20), .B1(new_n429), .B2(new_n203), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n251), .A2(G159), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n427), .A2(KEYINPUT16), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT16), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n424), .B1(new_n423), .B2(G20), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n345), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n254), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n435), .B1(new_n438), .B2(new_n432), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n434), .A2(new_n439), .A3(new_n266), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n393), .A2(new_n274), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n363), .A2(new_n283), .A3(new_n364), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n441), .B1(new_n442), .B2(new_n393), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n419), .A2(new_n422), .A3(new_n440), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT17), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n440), .A2(new_n443), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT17), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(new_n422), .A4(new_n419), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n420), .A2(new_n339), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n420), .A2(G169), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n446), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT18), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT18), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n446), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n407), .A2(new_n450), .A3(new_n459), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n342), .A2(new_n384), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n462), .B(new_n225), .C1(G33), .C2(new_n244), .ZN(new_n463));
  INV_X1    g0263(.A(G116), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G20), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(new_n266), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT20), .ZN(new_n467));
  OR2_X1    g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n467), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n468), .A2(new_n469), .B1(new_n464), .B2(new_n280), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n273), .A2(G33), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G116), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT87), .B1(new_n282), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT87), .ZN(new_n475));
  AOI211_X1 g0275(.A(new_n475), .B(new_n472), .C1(new_n278), .C2(new_n281), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n470), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT81), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT5), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n478), .B1(new_n479), .B2(G41), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n291), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n481));
  INV_X1    g0281(.A(G45), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(G1), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n479), .A2(G41), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n480), .A2(new_n481), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(G270), .A3(new_n301), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n273), .A2(G45), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n487), .B1(new_n479), .B2(G41), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n488), .A2(G274), .A3(new_n481), .A4(new_n480), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n345), .A2(G303), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n306), .A2(new_n308), .A3(G264), .A4(G1698), .ZN(new_n492));
  INV_X1    g0292(.A(G257), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n491), .B(new_n492), .C1(new_n493), .C2(new_n313), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n315), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n401), .B1(new_n490), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT21), .B1(new_n477), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n490), .A2(new_n495), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(new_n323), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n287), .B1(new_n490), .B2(new_n495), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n499), .A2(new_n477), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT88), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n486), .A2(new_n489), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n315), .B2(new_n494), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n496), .A2(KEYINPUT21), .B1(new_n504), .B2(G179), .ZN(new_n505));
  INV_X1    g0305(.A(new_n477), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n498), .A2(KEYINPUT21), .A3(G169), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n490), .A2(new_n495), .A3(G179), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(KEYINPUT88), .A3(new_n477), .ZN(new_n511));
  AOI211_X1 g0311(.A(new_n497), .B(new_n501), .C1(new_n507), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n485), .A2(new_n301), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n489), .B1(new_n513), .B2(new_n493), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n306), .A2(new_n308), .A3(G250), .A4(G1698), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n515), .A2(new_n462), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT4), .ZN(new_n517));
  INV_X1    g0317(.A(G244), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n517), .B1(new_n313), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g0319(.A(KEYINPUT67), .B(G1698), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n423), .A2(new_n520), .A3(KEYINPUT4), .A4(G244), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n516), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n514), .B1(new_n315), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(G107), .B1(new_n425), .B2(new_n426), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n242), .A2(KEYINPUT6), .A3(G97), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n246), .B2(KEYINPUT6), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n526), .A2(G20), .B1(G77), .B2(new_n251), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n277), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n280), .A2(new_n244), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n277), .A2(new_n274), .A3(new_n471), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n529), .B1(new_n530), .B2(new_n244), .ZN(new_n531));
  OAI22_X1  g0331(.A1(new_n523), .A2(G169), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n522), .A2(new_n315), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT80), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n522), .A2(KEYINPUT80), .A3(new_n315), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n514), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n532), .B1(new_n537), .B2(new_n339), .ZN(new_n538));
  INV_X1    g0338(.A(new_n514), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n522), .A2(KEYINPUT80), .A3(new_n315), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT80), .B1(new_n522), .B2(new_n315), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT82), .B1(new_n542), .B2(G200), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n533), .A2(new_n539), .A3(G190), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT83), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n528), .A2(new_n531), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n523), .A2(KEYINPUT83), .A3(G190), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n542), .A2(KEYINPUT82), .A3(G200), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n538), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n396), .A2(new_n530), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT85), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n260), .A2(G97), .A3(new_n261), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n225), .B1(new_n310), .B2(new_n557), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n211), .A2(new_n244), .A3(new_n242), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n306), .A2(new_n308), .A3(new_n225), .A4(G68), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n555), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n556), .A2(new_n557), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n565), .A2(KEYINPUT85), .A3(new_n561), .A4(new_n562), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n266), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT86), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n396), .A2(new_n280), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n568), .B1(new_n567), .B2(new_n569), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n554), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n306), .A2(new_n308), .A3(G244), .A4(G1698), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G33), .A2(G116), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n423), .A2(new_n520), .A3(G238), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n301), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n487), .A2(KEYINPUT84), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT84), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n579), .A2(new_n273), .A3(G45), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n301), .A2(G250), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n581), .A2(new_n582), .B1(new_n294), .B2(new_n487), .ZN(new_n583));
  OAI21_X1  g0383(.A(G169), .B1(new_n577), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n576), .A2(new_n574), .A3(new_n573), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n315), .ZN(new_n586));
  INV_X1    g0386(.A(new_n583), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(G179), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n572), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n306), .A2(new_n308), .A3(G257), .A4(G1698), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G294), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n591), .B(new_n592), .C1(new_n313), .C2(new_n212), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n315), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n485), .A2(G264), .A3(new_n301), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n489), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G169), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(KEYINPUT92), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT92), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n485), .A2(new_n599), .A3(G264), .A4(new_n301), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n485), .A2(new_n294), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n602), .B1(new_n593), .B2(new_n315), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(G179), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n597), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n306), .A2(new_n308), .A3(new_n225), .A4(G87), .ZN(new_n606));
  AND2_X1   g0406(.A1(KEYINPUT89), .A2(KEYINPUT22), .ZN(new_n607));
  NOR2_X1   g0407(.A1(KEYINPUT89), .A2(KEYINPUT22), .ZN(new_n608));
  OR2_X1    g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n607), .A2(new_n608), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n611), .A2(new_n423), .A3(new_n225), .A4(G87), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT90), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n242), .A2(G20), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n613), .B1(new_n614), .B2(KEYINPUT23), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n225), .A2(G107), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT23), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(KEYINPUT90), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n574), .A2(G20), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n620), .B1(KEYINPUT23), .B2(new_n614), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n610), .A2(new_n612), .A3(new_n619), .A4(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT24), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI22_X1  g0424(.A1(new_n616), .A2(new_n617), .B1(G20), .B2(new_n574), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(new_n615), .B2(new_n618), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n626), .A2(KEYINPUT24), .A3(new_n610), .A4(new_n612), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n624), .A2(new_n266), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n280), .A2(KEYINPUT25), .A3(new_n242), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(KEYINPUT91), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT25), .B1(new_n280), .B2(new_n242), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n629), .A2(KEYINPUT91), .ZN(new_n633));
  INV_X1    g0433(.A(new_n530), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n632), .A2(new_n633), .B1(new_n634), .B2(G107), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n628), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n605), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(G200), .B1(new_n601), .B2(new_n603), .ZN(new_n638));
  AND4_X1   g0438(.A1(new_n323), .A2(new_n594), .A3(new_n489), .A4(new_n595), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n628), .B(new_n635), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n287), .B1(new_n586), .B2(new_n587), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n577), .A2(new_n583), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n642), .B1(G190), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n634), .A2(G87), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n644), .B(new_n645), .C1(new_n570), .C2(new_n571), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n590), .A2(new_n641), .A3(new_n646), .ZN(new_n647));
  AND4_X1   g0447(.A1(new_n461), .A2(new_n512), .A3(new_n552), .A4(new_n647), .ZN(G372));
  INV_X1    g0448(.A(new_n368), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n455), .A2(KEYINPUT95), .A3(new_n457), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT95), .B1(new_n455), .B2(new_n457), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n338), .A2(new_n340), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n331), .A2(new_n404), .B1(new_n286), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n450), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n382), .A2(new_n383), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n649), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n567), .A2(new_n569), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(KEYINPUT86), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n553), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT93), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n584), .A2(new_n663), .A3(new_n588), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n663), .B1(new_n584), .B2(new_n588), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n538), .B(new_n646), .C1(new_n662), .C2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n589), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n538), .B(new_n646), .C1(new_n662), .C2(new_n670), .ZN(new_n671));
  XOR2_X1   g0471(.A(KEYINPUT94), .B(KEYINPUT26), .Z(new_n672));
  OAI22_X1  g0472(.A1(new_n669), .A2(KEYINPUT26), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n660), .A2(new_n661), .B1(G87), .B2(new_n634), .ZN(new_n674));
  INV_X1    g0474(.A(new_n666), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n664), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n674), .A2(new_n644), .B1(new_n676), .B2(new_n572), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n497), .B1(new_n477), .B2(new_n510), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n637), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n552), .A2(new_n640), .A3(new_n677), .A4(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n676), .A2(new_n572), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n673), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n461), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n658), .A2(new_n683), .ZN(G369));
  INV_X1    g0484(.A(G13), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G20), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n273), .ZN(new_n687));
  XOR2_X1   g0487(.A(new_n687), .B(KEYINPUT96), .Z(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G213), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g0492(.A(KEYINPUT97), .B(G343), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n477), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n512), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n678), .B2(new_n696), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n695), .A2(new_n636), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n641), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n637), .B2(new_n694), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n507), .A2(new_n511), .ZN(new_n705));
  INV_X1    g0505(.A(new_n497), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n695), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n641), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n637), .B2(new_n695), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n704), .A2(new_n710), .ZN(G399));
  INV_X1    g0511(.A(new_n219), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G41), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n560), .A2(G116), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(G1), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(new_n222), .B2(new_n714), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT28), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT29), .ZN(new_n719));
  INV_X1    g0519(.A(new_n681), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT82), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n537), .B2(new_n287), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n721), .A2(new_n723), .A3(new_n551), .ZN(new_n724));
  INV_X1    g0524(.A(new_n538), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n681), .A2(new_n640), .A3(new_n646), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n705), .A2(new_n706), .A3(new_n637), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n720), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n671), .A2(new_n672), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT100), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n669), .A2(KEYINPUT26), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n671), .A2(KEYINPUT100), .A3(new_n672), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n730), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n719), .B1(new_n737), .B2(new_n694), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n682), .A2(new_n719), .A3(new_n694), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n504), .A2(new_n643), .A3(G179), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n601), .A2(new_n603), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n741), .A2(new_n542), .A3(new_n742), .ZN(new_n743));
  AND3_X1   g0543(.A1(new_n643), .A2(new_n594), .A3(new_n601), .ZN(new_n744));
  INV_X1    g0544(.A(new_n509), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n744), .A2(new_n745), .A3(KEYINPUT30), .A4(new_n523), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT30), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n523), .A2(new_n504), .A3(G179), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n643), .A2(new_n594), .A3(new_n601), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n743), .A2(new_n746), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(KEYINPUT99), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT99), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n743), .A2(new_n746), .A3(new_n750), .A4(new_n753), .ZN(new_n754));
  AND3_X1   g0554(.A1(new_n752), .A2(new_n695), .A3(new_n754), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n647), .A2(new_n552), .A3(new_n512), .A4(new_n694), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n755), .B1(new_n756), .B2(KEYINPUT31), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n751), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT98), .ZN(new_n759));
  OAI21_X1  g0559(.A(G330), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n739), .A2(new_n740), .A3(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n718), .B1(new_n762), .B2(G1), .ZN(G364));
  XNOR2_X1  g0563(.A(new_n699), .B(KEYINPUT101), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n273), .B1(new_n686), .B2(G45), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n713), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n764), .B(new_n768), .C1(G330), .C2(new_n698), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n769), .A2(KEYINPUT102), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n712), .A2(new_n345), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G355), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(G116), .B2(new_n219), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n712), .A2(new_n423), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(new_n223), .B2(new_n290), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n241), .A2(G45), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n773), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n224), .B1(G20), .B2(new_n401), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n767), .B1(new_n778), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n339), .A2(new_n287), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n225), .A2(new_n323), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G326), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n287), .A2(G179), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G303), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n788), .A2(new_n789), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n339), .A2(G200), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n787), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n423), .B(new_n793), .C1(G322), .C2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n225), .A2(G190), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n794), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G179), .A2(G200), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G311), .A2(new_n800), .B1(new_n803), .B2(G329), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n786), .A2(new_n798), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(KEYINPUT33), .B(G317), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n798), .A2(new_n790), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n806), .A2(new_n807), .B1(new_n809), .B2(G283), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n225), .B1(new_n801), .B2(G190), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G294), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n797), .A2(new_n804), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n423), .B1(new_n788), .B2(new_n209), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n803), .A2(G159), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n815), .B1(KEYINPUT32), .B2(new_n816), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n816), .A2(KEYINPUT32), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n808), .A2(new_n242), .ZN(new_n819));
  INV_X1    g0619(.A(new_n791), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(G87), .B2(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G58), .A2(new_n796), .B1(new_n800), .B2(G77), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n817), .A2(new_n818), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n811), .A2(new_n244), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G68), .B2(new_n806), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT103), .Z(new_n826));
  OAI21_X1  g0626(.A(new_n814), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n785), .B1(new_n827), .B2(new_n782), .ZN(new_n828));
  INV_X1    g0628(.A(new_n781), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n698), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n769), .A2(KEYINPUT102), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n770), .A2(new_n830), .A3(new_n831), .ZN(G396));
  AOI22_X1  g0632(.A1(G87), .A2(new_n809), .B1(new_n803), .B2(G311), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n833), .B1(new_n242), .B2(new_n791), .C1(new_n792), .C2(new_n788), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n345), .B1(new_n799), .B2(new_n464), .ZN(new_n835));
  INV_X1    g0635(.A(G283), .ZN(new_n836));
  INV_X1    g0636(.A(G294), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n836), .A2(new_n805), .B1(new_n795), .B2(new_n837), .ZN(new_n838));
  NOR4_X1   g0638(.A1(new_n834), .A2(new_n824), .A3(new_n835), .A4(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT104), .ZN(new_n840));
  INV_X1    g0640(.A(G132), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n423), .B1(new_n802), .B2(new_n841), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n791), .A2(new_n209), .B1(new_n808), .B2(new_n254), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n842), .B(new_n843), .C1(G58), .C2(new_n812), .ZN(new_n844));
  INV_X1    g0644(.A(G137), .ZN(new_n845));
  INV_X1    g0645(.A(G150), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n788), .A2(new_n845), .B1(new_n805), .B2(new_n846), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT105), .Z(new_n848));
  AOI22_X1  g0648(.A1(G143), .A2(new_n796), .B1(new_n800), .B2(G159), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT34), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n844), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(new_n851), .B2(new_n850), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n782), .B1(new_n840), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n782), .A2(new_n779), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n768), .B1(new_n257), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n404), .A2(new_n694), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n405), .A2(new_n406), .B1(new_n695), .B2(new_n400), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n857), .B1(new_n858), .B2(new_n404), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n854), .B(new_n856), .C1(new_n860), .C2(new_n780), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n682), .A2(new_n694), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n859), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n682), .A2(new_n694), .A3(new_n860), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n767), .B1(new_n865), .B2(new_n760), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n865), .A2(new_n760), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n861), .B1(new_n867), .B2(new_n868), .ZN(G384));
  NOR2_X1   g0669(.A1(new_n202), .A2(new_n254), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n222), .A2(new_n257), .A3(new_n429), .ZN(new_n871));
  OAI211_X1 g0671(.A(G1), .B(new_n685), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n872), .B(KEYINPUT106), .Z(new_n873));
  OR2_X1    g0673(.A1(new_n526), .A2(KEYINPUT35), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n874), .A2(G116), .A3(new_n226), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(KEYINPUT35), .B2(new_n526), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n873), .B1(KEYINPUT36), .B2(new_n876), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n755), .A2(KEYINPUT31), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n461), .B1(new_n757), .B2(new_n878), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT109), .Z(new_n880));
  NAND2_X1  g0680(.A1(new_n446), .A2(new_n692), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(new_n459), .B2(new_n450), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n444), .A2(new_n454), .A3(new_n881), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT37), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n883), .B(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n882), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n450), .B1(new_n650), .B2(new_n651), .ZN(new_n888));
  INV_X1    g0688(.A(new_n881), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n444), .A2(new_n881), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(new_n884), .A3(new_n454), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n446), .A2(new_n453), .A3(KEYINPUT95), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT95), .B1(new_n446), .B2(new_n453), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n884), .B1(new_n895), .B2(new_n891), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n892), .B1(new_n896), .B2(KEYINPUT108), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT95), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n454), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n446), .A2(new_n453), .A3(KEYINPUT95), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n899), .A2(new_n444), .A3(new_n881), .A4(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(KEYINPUT108), .A3(KEYINPUT37), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n890), .B1(new_n897), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n887), .B1(new_n904), .B2(new_n886), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n695), .A2(new_n286), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n341), .B(new_n906), .C1(new_n330), .C2(new_n329), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n653), .A2(new_n286), .A3(new_n695), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n859), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n757), .B2(new_n878), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT40), .B1(new_n905), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n907), .A2(new_n908), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n860), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n756), .A2(KEYINPUT31), .ZN(new_n914));
  INV_X1    g0714(.A(new_n755), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n755), .A2(KEYINPUT31), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n886), .B1(new_n885), .B2(new_n882), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n889), .B1(new_n655), .B2(new_n458), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n883), .A2(KEYINPUT37), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n892), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(KEYINPUT38), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT40), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n918), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n911), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(G330), .B1(new_n880), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n926), .B2(new_n880), .ZN(new_n928));
  INV_X1    g0728(.A(new_n912), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT38), .B1(new_n920), .B2(new_n922), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n887), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n857), .B(KEYINPUT107), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n929), .B(new_n931), .C1(new_n864), .C2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n653), .A2(new_n286), .A3(new_n694), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT39), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n883), .A2(KEYINPUT37), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT108), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n939), .A2(new_n902), .B1(new_n889), .B2(new_n888), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n935), .B(new_n923), .C1(new_n940), .C2(KEYINPUT38), .ZN(new_n941));
  OAI21_X1  g0741(.A(KEYINPUT39), .B1(new_n887), .B2(new_n930), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n934), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n652), .A2(new_n692), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n933), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n740), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n461), .B1(new_n738), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n658), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n945), .B(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n928), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT110), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n928), .A2(new_n949), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n951), .B(new_n952), .C1(new_n273), .C2(new_n686), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n950), .A2(KEYINPUT110), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n877), .B1(KEYINPUT36), .B2(new_n876), .C1(new_n953), .C2(new_n954), .ZN(G367));
  NOR2_X1   g0755(.A1(new_n694), .A2(new_n547), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n726), .A2(new_n956), .B1(new_n725), .B2(new_n694), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n957), .A2(KEYINPUT111), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(KEYINPUT111), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n710), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT45), .Z(new_n962));
  NOR2_X1   g0762(.A1(new_n958), .A2(new_n959), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n709), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT44), .Z(new_n965));
  NAND2_X1  g0765(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n704), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n708), .B1(new_n703), .B2(new_n707), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n967), .B1(new_n764), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n761), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n713), .B(KEYINPUT41), .Z(new_n971));
  OAI21_X1  g0771(.A(new_n765), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n963), .A2(new_n708), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT42), .Z(new_n974));
  INV_X1    g0774(.A(KEYINPUT43), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n674), .A2(new_n694), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n720), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n677), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n977), .B1(new_n978), .B2(new_n976), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n963), .A2(new_n637), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n695), .B1(new_n981), .B2(new_n725), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n974), .A2(new_n975), .A3(new_n980), .A4(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n704), .A2(new_n963), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n980), .A2(new_n975), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n979), .A2(KEYINPUT43), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n973), .B(KEYINPUT42), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n986), .B(new_n987), .C1(new_n988), .C2(new_n982), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n984), .A2(new_n985), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n984), .A2(new_n989), .ZN(new_n991));
  INV_X1    g0791(.A(new_n985), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n972), .A2(new_n990), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n980), .A2(new_n781), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n237), .A2(new_n775), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n783), .B1(new_n396), .B2(new_n219), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n767), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n808), .A2(new_n257), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n795), .A2(new_n846), .B1(new_n802), .B2(new_n845), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n788), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n999), .B(new_n1000), .C1(G143), .C2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n811), .A2(new_n254), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n345), .B1(new_n806), .B2(G159), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n800), .A2(new_n202), .B1(new_n820), .B2(G58), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n809), .A2(G97), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n836), .B2(new_n799), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n423), .B(new_n1009), .C1(G303), .C2(new_n796), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n1001), .A2(G311), .B1(new_n803), .B2(G317), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1010), .B(new_n1011), .C1(new_n837), .C2(new_n805), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n820), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT46), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n791), .B2(new_n464), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1013), .B(new_n1015), .C1(new_n242), .C2(new_n811), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1007), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT47), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n782), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n998), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n995), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n994), .A2(new_n1023), .ZN(G387));
  INV_X1    g0824(.A(new_n969), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n761), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n762), .A2(new_n969), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1026), .A2(new_n1027), .A3(new_n713), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n703), .A2(new_n829), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n233), .A2(new_n288), .A3(new_n289), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n715), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n1030), .A2(new_n774), .B1(new_n1031), .B2(new_n771), .ZN(new_n1032));
  AOI21_X1  g0832(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n393), .A2(new_n209), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n715), .B(new_n1033), .C1(new_n1034), .C2(KEYINPUT50), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(KEYINPUT50), .B2(new_n1034), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1032), .A2(new_n1036), .B1(G107), .B2(new_n219), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n768), .B1(new_n1037), .B2(new_n783), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n806), .A2(new_n393), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n820), .A2(G77), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1039), .A2(new_n1040), .A3(new_n1008), .A4(new_n423), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n396), .A2(new_n811), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n795), .A2(new_n209), .B1(new_n802), .B2(new_n846), .ZN(new_n1043));
  INV_X1    g0843(.A(G159), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n788), .A2(new_n1044), .B1(new_n799), .B2(new_n254), .ZN(new_n1045));
  NOR4_X1   g0845(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .A4(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n1001), .A2(G322), .B1(new_n800), .B2(G303), .ZN(new_n1047));
  INV_X1    g0847(.A(G311), .ZN(new_n1048));
  INV_X1    g0848(.A(G317), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1047), .B1(new_n1048), .B2(new_n805), .C1(new_n1049), .C2(new_n795), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT112), .Z(new_n1051));
  OR2_X1    g0851(.A1(new_n1051), .A2(KEYINPUT48), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(KEYINPUT48), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n820), .A2(G294), .B1(new_n812), .B2(G283), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT49), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n345), .B1(new_n802), .B2(new_n789), .C1(new_n464), .C2(new_n808), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1046), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1038), .B1(new_n1060), .B2(new_n1020), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1028), .B1(new_n765), .B2(new_n1025), .C1(new_n1029), .C2(new_n1061), .ZN(G393));
  INV_X1    g0862(.A(new_n1027), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n966), .A2(new_n967), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n962), .A2(new_n704), .A3(new_n965), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n966), .A2(new_n1063), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n713), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1064), .A2(new_n766), .A3(new_n1065), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n248), .A2(new_n775), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n783), .B1(new_n244), .B2(new_n219), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n767), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n788), .A2(new_n1049), .B1(new_n795), .B2(new_n1048), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT52), .Z(new_n1075));
  AOI211_X1 g0875(.A(new_n423), .B(new_n819), .C1(G116), .C2(new_n812), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G294), .A2(new_n800), .B1(new_n803), .B2(G322), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(G283), .A2(new_n820), .B1(new_n806), .B2(G303), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n811), .A2(new_n257), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n345), .B(new_n1080), .C1(G87), .C2(new_n809), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G68), .A2(new_n820), .B1(new_n803), .B2(G143), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n806), .A2(new_n202), .B1(new_n800), .B2(new_n393), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n788), .A2(new_n846), .B1(new_n795), .B2(new_n1044), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT51), .Z(new_n1086));
  OAI22_X1  g0886(.A1(new_n1075), .A2(new_n1079), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1073), .B1(new_n1087), .B2(new_n782), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n960), .B2(new_n829), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1070), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1069), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(G390));
  AND2_X1   g0892(.A1(new_n941), .A2(new_n942), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n929), .B1(new_n864), .B2(new_n932), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n934), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(G330), .B(new_n860), .C1(new_n757), .C2(new_n759), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1097), .A2(new_n929), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT113), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n671), .A2(KEYINPUT100), .A3(new_n672), .ZN(new_n1100));
  AOI21_X1  g0900(.A(KEYINPUT100), .B1(new_n671), .B2(new_n672), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT26), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n668), .A2(new_n1102), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n1100), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n677), .A2(new_n724), .A3(new_n725), .A4(new_n640), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n729), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n681), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n694), .B(new_n860), .C1(new_n1104), .C2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n932), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n912), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n905), .A2(new_n1095), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1099), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n929), .B1(new_n1108), .B2(new_n932), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n939), .A2(new_n902), .ZN(new_n1114));
  AOI21_X1  g0914(.A(KEYINPUT38), .B1(new_n1114), .B2(new_n890), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n934), .B1(new_n1115), .B2(new_n887), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n1113), .A2(new_n1116), .A3(KEYINPUT113), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1096), .B(new_n1098), .C1(new_n1112), .C2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1110), .A2(new_n1099), .A3(new_n1111), .ZN(new_n1119));
  OAI21_X1  g0919(.A(KEYINPUT113), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n864), .A2(new_n932), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n912), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n934), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1119), .A2(new_n1120), .B1(new_n1123), .B2(new_n1093), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n918), .A2(G330), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1118), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1093), .A2(new_n779), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n855), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n767), .B1(new_n1129), .B2(new_n393), .ZN(new_n1130));
  INV_X1    g0930(.A(G128), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n788), .A2(new_n1131), .B1(new_n795), .B2(new_n841), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT117), .ZN(new_n1133));
  XOR2_X1   g0933(.A(KEYINPUT54), .B(G143), .Z(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n1135), .A2(new_n799), .B1(new_n845), .B2(new_n805), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G159), .B2(new_n812), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n791), .A2(new_n846), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT53), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1133), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(G125), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n423), .B1(new_n802), .B2(new_n1141), .C1(new_n201), .C2(new_n808), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT116), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n345), .B1(new_n791), .B2(new_n211), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT118), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n254), .A2(new_n808), .B1(new_n799), .B2(new_n244), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1146), .A2(new_n1080), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n806), .A2(G107), .B1(new_n803), .B2(G294), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(G283), .A2(new_n1001), .B1(new_n796), .B2(G116), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n1140), .A2(new_n1143), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1130), .B1(new_n1151), .B2(new_n782), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1127), .A2(new_n766), .B1(new_n1128), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT115), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1097), .A2(new_n929), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1125), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n1121), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1109), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n757), .A2(new_n878), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n860), .A2(G330), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n929), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1098), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1157), .A2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n461), .B(G330), .C1(new_n757), .C2(new_n878), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n947), .A2(new_n658), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(KEYINPUT114), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1165), .B1(new_n1157), .B2(new_n1162), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT114), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n714), .B1(new_n1172), .B2(new_n1126), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1118), .B(new_n1169), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1154), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1176));
  AOI211_X1 g0976(.A(KEYINPUT114), .B(new_n1165), .C1(new_n1157), .C2(new_n1162), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1126), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AND4_X1   g0978(.A1(new_n1154), .A2(new_n1178), .A3(new_n713), .A4(new_n1174), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1153), .B1(new_n1175), .B2(new_n1179), .ZN(G378));
  INV_X1    g0980(.A(KEYINPUT57), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1174), .A2(new_n1166), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n944), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(new_n1122), .B2(new_n931), .C1(new_n1093), .C2(new_n934), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n377), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n692), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n384), .A2(new_n1187), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n368), .B(new_n1186), .C1(new_n382), .C2(new_n383), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1190), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n926), .B2(G330), .ZN(new_n1195));
  INV_X1    g0995(.A(G330), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1196), .B(new_n1193), .C1(new_n911), .C2(new_n925), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1184), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT40), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n923), .B1(new_n940), .B2(KEYINPUT38), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n918), .B2(new_n1200), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n910), .A2(new_n931), .A3(KEYINPUT40), .ZN(new_n1202));
  OAI21_X1  g1002(.A(G330), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n1193), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n926), .A2(G330), .A3(new_n1194), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(new_n945), .A3(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1198), .A2(new_n1206), .A3(KEYINPUT119), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT119), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1184), .B(new_n1208), .C1(new_n1195), .C2(new_n1197), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1181), .B1(new_n1182), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT120), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1174), .A2(new_n1166), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1214), .A2(new_n1209), .A3(new_n1207), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1215), .A2(KEYINPUT120), .A3(new_n1181), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1198), .A2(new_n1206), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1217), .A2(new_n1181), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n714), .B1(new_n1218), .B2(new_n1214), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1213), .A2(new_n1216), .A3(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1210), .A2(new_n765), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1193), .A2(new_n779), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n767), .B1(new_n1129), .B2(new_n202), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n1131), .A2(new_n795), .B1(new_n805), .B2(new_n841), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n820), .A2(new_n1134), .B1(new_n800), .B2(G137), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n1141), .B2(new_n788), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1224), .B(new_n1226), .C1(G150), .C2(new_n812), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT59), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n809), .A2(G159), .ZN(new_n1231));
  AOI211_X1 g1031(.A(G33), .B(G41), .C1(new_n803), .C2(G124), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(G116), .A2(new_n1001), .B1(new_n806), .B2(G97), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n242), .B2(new_n795), .C1(new_n396), .C2(new_n799), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1040), .A2(new_n291), .A3(new_n345), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n808), .A2(new_n428), .B1(new_n802), .B2(new_n836), .ZN(new_n1237));
  NOR4_X1   g1037(.A1(new_n1235), .A2(new_n1003), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1238), .A2(KEYINPUT58), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(KEYINPUT58), .ZN(new_n1240));
  AOI21_X1  g1040(.A(G50), .B1(new_n259), .B2(new_n291), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n423), .B2(G41), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1233), .A2(new_n1239), .A3(new_n1240), .A4(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1223), .B1(new_n1243), .B2(new_n782), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1221), .B1(new_n1222), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1220), .A2(new_n1245), .ZN(G375));
  NOR2_X1   g1046(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1247), .A2(new_n971), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1172), .A2(new_n1248), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n1135), .A2(new_n805), .B1(new_n1044), .B2(new_n791), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n795), .A2(new_n845), .B1(new_n802), .B2(new_n1131), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n423), .B1(new_n808), .B2(new_n428), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n788), .A2(new_n841), .B1(new_n799), .B2(new_n846), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1253), .B(new_n1254), .C1(G50), .C2(new_n812), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n244), .A2(new_n791), .B1(new_n805), .B2(new_n464), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n788), .A2(new_n837), .B1(new_n795), .B2(new_n836), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n799), .A2(new_n242), .B1(new_n802), .B2(new_n792), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n345), .B1(new_n808), .B2(new_n257), .ZN(new_n1259));
  NOR4_X1   g1059(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1042), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1252), .A2(new_n1255), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n767), .B1(G68), .B2(new_n1129), .C1(new_n1262), .C2(new_n1020), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n929), .B2(new_n779), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n1163), .B2(new_n766), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1249), .A2(new_n1265), .ZN(G381));
  INV_X1    g1066(.A(G375), .ZN(new_n1267));
  OR2_X1    g1067(.A1(new_n1267), .A2(KEYINPUT121), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(KEYINPUT121), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1270), .A2(new_n1153), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1268), .A2(new_n1269), .A3(new_n1271), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n994), .A2(new_n1023), .ZN(new_n1273));
  INV_X1    g1073(.A(G384), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(G393), .A2(G396), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1273), .A2(new_n1091), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  OR3_X1    g1076(.A1(new_n1272), .A2(G381), .A3(new_n1276), .ZN(G407));
  OAI211_X1 g1077(.A(G407), .B(G213), .C1(new_n693), .C2(new_n1272), .ZN(G409));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n693), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(G213), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1220), .A2(G378), .A3(new_n1245), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1222), .A2(new_n1244), .ZN(new_n1284));
  OAI221_X1 g1084(.A(new_n1284), .B1(new_n765), .B2(new_n1217), .C1(new_n1215), .C2(new_n971), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1271), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1282), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1157), .A2(new_n1165), .A3(new_n1162), .A4(KEYINPUT60), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT122), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1288), .B(new_n1289), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n713), .B(new_n1167), .C1(new_n1247), .C2(KEYINPUT60), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1265), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1274), .ZN(new_n1293));
  OAI211_X1 g1093(.A(G384), .B(new_n1265), .C1(new_n1290), .C2(new_n1291), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1293), .A2(KEYINPUT123), .A3(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT123), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(KEYINPUT125), .B(G2897), .ZN(new_n1297));
  OAI22_X1  g1097(.A1(new_n1295), .A2(new_n1296), .B1(new_n1281), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(G2897), .A3(new_n1282), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1279), .B1(new_n1287), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT127), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  OAI211_X1 g1104(.A(KEYINPUT127), .B(new_n1279), .C1(new_n1287), .C2(new_n1301), .ZN(new_n1305));
  OR2_X1    g1105(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1287), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(KEYINPUT62), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT62), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1287), .A2(new_n1309), .A3(new_n1306), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1304), .A2(new_n1305), .A3(new_n1308), .A4(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1273), .A2(G390), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(G387), .A2(new_n1091), .ZN(new_n1313));
  XOR2_X1   g1113(.A(G393), .B(G396), .Z(new_n1314));
  AND4_X1   g1114(.A1(KEYINPUT126), .A2(new_n1312), .A3(new_n1313), .A4(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT126), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1313), .A2(new_n1316), .ZN(new_n1317));
  AOI22_X1  g1117(.A1(new_n1317), .A2(new_n1314), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1315), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1311), .A2(new_n1320), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1319), .B(new_n1279), .C1(new_n1287), .C2(new_n1301), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1307), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT124), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1287), .A2(KEYINPUT63), .A3(new_n1306), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1307), .A2(KEYINPUT124), .A3(new_n1324), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1323), .A2(new_n1327), .A3(new_n1328), .A4(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1321), .A2(new_n1330), .ZN(G405));
  NAND2_X1  g1131(.A1(G375), .A2(new_n1271), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1283), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1306), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1332), .A2(new_n1283), .A3(new_n1299), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(new_n1336), .B(new_n1320), .ZN(G402));
endmodule


