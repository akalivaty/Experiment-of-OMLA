//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1221, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  XOR2_X1   g0018(.A(KEYINPUT64), .B(G238), .Z(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT65), .B(G77), .Z(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT66), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT68), .ZN(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  AOI21_X1  g0047(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT70), .ZN(new_n249));
  AND2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(KEYINPUT70), .A3(G1698), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n257), .A2(G223), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(new_n253), .ZN(new_n259));
  INV_X1    g0059(.A(G222), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n259), .A2(new_n260), .B1(new_n222), .B2(new_n255), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n248), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  OAI211_X1 g0064(.A(G1), .B(G13), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G45), .ZN(new_n266));
  AOI21_X1  g0066(.A(G1), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AND3_X1   g0067(.A1(new_n265), .A2(G274), .A3(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n248), .A2(new_n267), .ZN(new_n269));
  XOR2_X1   g0069(.A(KEYINPUT69), .B(G226), .Z(new_n270));
  AOI21_X1  g0070(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n262), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G190), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n206), .A2(G20), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G50), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT71), .ZN(new_n277));
  INV_X1    g0077(.A(G13), .ZN(new_n278));
  NOR3_X1   g0078(.A1(new_n278), .A2(new_n207), .A3(G1), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n215), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n279), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n277), .A2(new_n283), .B1(G50), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n281), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n263), .A2(G20), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n288), .A2(new_n289), .B1(G150), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n286), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n285), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT9), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n294), .B(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT74), .B(G200), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n272), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n274), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT10), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT10), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n274), .A2(new_n296), .A3(new_n302), .A4(new_n299), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n273), .A2(G169), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(new_n294), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(G179), .B2(new_n272), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n279), .A2(new_n220), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT12), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n289), .A2(G77), .B1(G20), .B2(new_n220), .ZN(new_n311));
  INV_X1    g0111(.A(new_n290), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n311), .B1(new_n201), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n313), .A2(KEYINPUT11), .A3(new_n281), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n282), .A2(G68), .A3(new_n275), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n310), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT11), .B1(new_n313), .B2(new_n281), .ZN(new_n317));
  OR3_X1    g0117(.A1(new_n316), .A2(KEYINPUT75), .A3(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT75), .B1(new_n316), .B2(new_n317), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n255), .A2(G232), .A3(G1698), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G33), .A2(G97), .ZN(new_n322));
  INV_X1    g0122(.A(G226), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n321), .B(new_n322), .C1(new_n259), .C2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n248), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT13), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n268), .B1(G238), .B2(new_n269), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n326), .B1(new_n325), .B2(new_n327), .ZN(new_n329));
  OAI21_X1  g0129(.A(G169), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n325), .A2(new_n327), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT13), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G179), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n330), .A2(KEYINPUT14), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT14), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(new_n334), .B2(G169), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n320), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n334), .A2(G200), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n316), .A2(new_n317), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n332), .A2(G190), .A3(new_n333), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n222), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT15), .B(G87), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n345), .A2(G20), .B1(new_n347), .B2(new_n289), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n288), .A2(new_n290), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n286), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n282), .A2(G77), .A3(new_n275), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n345), .B2(new_n284), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n219), .B1(new_n254), .B2(new_n256), .ZN(new_n354));
  INV_X1    g0154(.A(G232), .ZN(new_n355));
  INV_X1    g0155(.A(G107), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n259), .A2(new_n355), .B1(new_n356), .B2(new_n255), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT73), .ZN(new_n358));
  OR3_X1    g0158(.A1(new_n354), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n358), .B1(new_n354), .B2(new_n357), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(new_n248), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n268), .B1(G244), .B2(new_n269), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT72), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n362), .B(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G190), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n353), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n297), .B1(new_n361), .B2(new_n364), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n365), .A2(G179), .ZN(new_n370));
  AOI21_X1  g0170(.A(G169), .B1(new_n361), .B2(new_n364), .ZN(new_n371));
  NOR3_X1   g0171(.A1(new_n370), .A2(new_n353), .A3(new_n371), .ZN(new_n372));
  NOR4_X1   g0172(.A1(new_n308), .A2(new_n344), .A3(new_n369), .A4(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n288), .A2(new_n275), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n283), .A2(new_n374), .B1(new_n284), .B2(new_n288), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G200), .ZN(new_n377));
  INV_X1    g0177(.A(G274), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n248), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n267), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n269), .A2(G232), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n323), .A2(G1698), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n255), .B(new_n383), .C1(G223), .C2(G1698), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G33), .A2(G87), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n265), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n377), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n384), .A2(new_n385), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n248), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n268), .B1(G232), .B2(new_n269), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n387), .B1(new_n391), .B2(G190), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT7), .B1(new_n252), .B2(new_n207), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  NOR4_X1   g0194(.A1(new_n250), .A2(new_n251), .A3(new_n394), .A4(G20), .ZN(new_n395));
  OAI21_X1  g0195(.A(G68), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G159), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n312), .A2(new_n397), .ZN(new_n398));
  AND2_X1   g0198(.A1(G58), .A2(G68), .ZN(new_n399));
  NOR2_X1   g0199(.A1(G58), .A2(G68), .ZN(new_n400));
  OAI21_X1  g0200(.A(G20), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT76), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI211_X1 g0203(.A(KEYINPUT76), .B(G20), .C1(new_n399), .C2(new_n400), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n398), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n396), .A2(new_n405), .A3(KEYINPUT16), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT16), .B1(new_n396), .B2(new_n405), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT77), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n281), .B(new_n406), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  AOI211_X1 g0209(.A(KEYINPUT77), .B(KEYINPUT16), .C1(new_n396), .C2(new_n405), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n376), .B(new_n392), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  XOR2_X1   g0211(.A(new_n411), .B(KEYINPUT17), .Z(new_n412));
  OAI21_X1  g0212(.A(new_n376), .B1(new_n409), .B2(new_n410), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT18), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n391), .A2(G169), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n335), .B2(new_n391), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n413), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n414), .B1(new_n413), .B2(new_n416), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT78), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n396), .A2(new_n405), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT16), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n408), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n406), .A2(new_n281), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n410), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n375), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n416), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT18), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT78), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n413), .A2(new_n414), .A3(new_n416), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n412), .B1(new_n419), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n373), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT24), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G33), .A2(G116), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(G20), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT23), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n207), .B2(G107), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n356), .A2(KEYINPUT23), .A3(G20), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n255), .A2(new_n207), .A3(G87), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT22), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT22), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n255), .A2(new_n445), .A3(new_n207), .A4(G87), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n442), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n435), .B1(new_n447), .B2(KEYINPUT85), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(KEYINPUT85), .B2(new_n447), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n447), .A2(KEYINPUT85), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n286), .B1(new_n450), .B2(new_n435), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n206), .A2(G33), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n282), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n279), .A2(KEYINPUT25), .A3(new_n356), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT25), .B1(new_n279), .B2(new_n356), .ZN(new_n457));
  OAI22_X1  g0257(.A1(new_n454), .A2(new_n356), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT86), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n458), .B1(new_n449), .B2(new_n451), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT86), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n255), .A2(G257), .A3(G1698), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n255), .A2(G250), .A3(new_n253), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G294), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n265), .B1(new_n468), .B2(KEYINPUT87), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT87), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n465), .A2(new_n466), .A3(new_n470), .A4(new_n467), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n266), .A2(G1), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT79), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n473), .B(new_n474), .C1(KEYINPUT5), .C2(new_n264), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n206), .B(G45), .C1(new_n264), .C2(KEYINPUT5), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT79), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n264), .A2(KEYINPUT5), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n475), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n379), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n476), .A2(KEYINPUT79), .B1(KEYINPUT5), .B2(new_n264), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n248), .B1(new_n481), .B2(new_n475), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G264), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n472), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G169), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n335), .B2(new_n484), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n461), .A2(new_n464), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(new_n377), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n469), .A2(new_n471), .B1(G264), .B2(new_n482), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(new_n366), .A3(new_n480), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n462), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT88), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(new_n462), .A3(KEYINPUT88), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n255), .A2(G264), .A3(G1698), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n255), .A2(G257), .A3(new_n253), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n252), .A2(G303), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT84), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n265), .B1(new_n500), .B2(new_n501), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n482), .A2(G270), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n480), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n284), .A2(G116), .ZN(new_n507));
  INV_X1    g0307(.A(new_n454), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(G116), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G283), .ZN(new_n510));
  INV_X1    g0310(.A(G97), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n510), .B(new_n207), .C1(G33), .C2(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n512), .B(new_n281), .C1(new_n207), .C2(G116), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT20), .ZN(new_n514));
  XNOR2_X1  g0314(.A(new_n513), .B(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n509), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n506), .A2(new_n517), .A3(new_n335), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n506), .A2(G200), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n505), .A2(new_n480), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n502), .B2(new_n503), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G190), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n520), .A2(new_n523), .A3(new_n517), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT21), .ZN(new_n525));
  INV_X1    g0325(.A(G169), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(new_n509), .B2(new_n515), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n525), .B1(new_n506), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n506), .A2(new_n525), .A3(new_n527), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n519), .B(new_n524), .C1(new_n528), .C2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(G87), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n454), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g0333(.A(new_n533), .B(KEYINPUT83), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n255), .A2(new_n207), .A3(G68), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT19), .ZN(new_n536));
  NOR2_X1   g0336(.A1(G97), .A2(G107), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n532), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n322), .A2(new_n207), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR4_X1   g0340(.A1(new_n263), .A2(new_n511), .A3(KEYINPUT19), .A4(G20), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n535), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT81), .ZN(new_n543));
  OR2_X1    g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n286), .B1(new_n542), .B2(new_n543), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n544), .A2(new_n545), .B1(new_n279), .B2(new_n346), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n534), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n255), .A2(G244), .A3(G1698), .ZN(new_n548));
  INV_X1    g0348(.A(G238), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n548), .B(new_n436), .C1(new_n259), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n248), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT80), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n206), .A2(G45), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G250), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n552), .B1(new_n248), .B2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n265), .A2(KEYINPUT80), .A3(G250), .A4(new_n553), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n555), .A2(new_n556), .B1(new_n379), .B2(new_n473), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n298), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n551), .A2(G190), .A3(new_n557), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(G169), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n335), .B2(new_n558), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n454), .A2(new_n346), .ZN(new_n564));
  XNOR2_X1  g0364(.A(new_n564), .B(KEYINPUT82), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n546), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n547), .A2(new_n561), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g0367(.A1(G257), .A2(new_n482), .B1(new_n479), .B2(new_n379), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n255), .A2(KEYINPUT4), .A3(G244), .A4(new_n253), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n252), .A2(new_n221), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n569), .B(new_n510), .C1(new_n570), .C2(KEYINPUT4), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n255), .A2(G250), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n253), .B1(new_n572), .B2(KEYINPUT4), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n248), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n356), .A2(KEYINPUT6), .A3(G97), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n511), .A2(new_n356), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(new_n537), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n576), .B1(new_n578), .B2(KEYINPUT6), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n579), .A2(G20), .B1(G77), .B2(new_n290), .ZN(new_n580));
  OAI21_X1  g0380(.A(G107), .B1(new_n393), .B2(new_n395), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n281), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n284), .A2(G97), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n508), .B2(G97), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n526), .A2(new_n575), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n568), .A2(new_n574), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n335), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n583), .A2(new_n585), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n575), .A2(G200), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n590), .B(new_n591), .C1(new_n366), .C2(new_n575), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n567), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n531), .A2(new_n593), .ZN(new_n594));
  AND4_X1   g0394(.A1(new_n434), .A2(new_n487), .A3(new_n496), .A4(new_n594), .ZN(G372));
  NAND2_X1  g0395(.A1(new_n506), .A2(new_n527), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT21), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n518), .B1(new_n597), .B2(new_n529), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n486), .A2(new_n460), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n534), .A2(new_n546), .A3(new_n559), .A4(new_n560), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n592), .A2(new_n601), .A3(new_n589), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n496), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT89), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n563), .A2(new_n566), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n605), .A2(new_n601), .A3(new_n588), .A4(new_n586), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT26), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n586), .A2(new_n588), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n610), .A2(new_n567), .A3(KEYINPUT89), .A4(KEYINPUT26), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n603), .A2(new_n612), .A3(new_n605), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n434), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n307), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n417), .A2(new_n418), .ZN(new_n616));
  INV_X1    g0416(.A(new_n339), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n372), .B2(new_n343), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n616), .B1(new_n618), .B2(new_n412), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n615), .B1(new_n619), .B2(new_n304), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n614), .A2(new_n620), .ZN(G369));
  NAND3_X1  g0421(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n622), .A2(KEYINPUT27), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(KEYINPUT27), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(G213), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g0425(.A(KEYINPUT90), .B(G343), .Z(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n517), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  MUX2_X1   g0430(.A(new_n598), .B(new_n531), .S(new_n630), .Z(new_n631));
  INV_X1    g0431(.A(G330), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT91), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n461), .A2(new_n464), .A3(new_n627), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n496), .A2(new_n487), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(new_n487), .B2(new_n628), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n633), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n634), .B1(new_n633), .B2(new_n637), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n598), .A2(new_n627), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n496), .A2(new_n643), .A3(new_n487), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n486), .A2(new_n460), .A3(new_n628), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n642), .A2(new_n646), .ZN(G399));
  INV_X1    g0447(.A(KEYINPUT92), .ZN(new_n648));
  INV_X1    g0448(.A(new_n210), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n648), .B1(new_n649), .B2(G41), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n210), .A2(KEYINPUT92), .A3(new_n264), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n538), .A2(G116), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(G1), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n213), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT28), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n613), .A2(new_n628), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(KEYINPUT29), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n487), .A2(new_n598), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n659), .A2(new_n496), .A3(new_n602), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n610), .A2(new_n567), .A3(KEYINPUT26), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n661), .A2(new_n609), .B1(new_n563), .B2(new_n566), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n627), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT29), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n658), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n594), .A2(new_n496), .A3(new_n487), .A4(new_n628), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n558), .A2(new_n335), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n522), .A2(new_n587), .A3(new_n489), .A4(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT93), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT30), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT30), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n669), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(G179), .B1(new_n551), .B2(new_n557), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n506), .A2(new_n484), .A3(new_n575), .A4(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n672), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n627), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT31), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n677), .A2(KEYINPUT31), .A3(new_n627), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n667), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n666), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n656), .B1(new_n685), .B2(G1), .ZN(G364));
  INV_X1    g0486(.A(new_n652), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n278), .A2(G20), .ZN(new_n688));
  AOI21_X1  g0488(.A(KEYINPUT94), .B1(new_n688), .B2(G45), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n206), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n688), .A2(KEYINPUT94), .A3(G45), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(G13), .A2(G33), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G20), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n631), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n215), .B1(G20), .B2(new_n526), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n210), .A2(new_n252), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n266), .B2(new_n214), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n246), .B2(new_n266), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n649), .A2(new_n252), .ZN(new_n705));
  INV_X1    g0505(.A(G116), .ZN(new_n706));
  AOI22_X1  g0506(.A1(new_n705), .A2(G355), .B1(new_n706), .B2(new_n649), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n701), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n207), .A2(G190), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n335), .A2(G200), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n255), .B1(new_n712), .B2(G311), .ZN(new_n713));
  INV_X1    g0513(.A(G322), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n207), .A2(new_n366), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n710), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n207), .A2(new_n335), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(new_n366), .A3(G200), .ZN(new_n718));
  XOR2_X1   g0518(.A(KEYINPUT33), .B(G317), .Z(new_n719));
  OAI221_X1 g0519(.A(new_n713), .B1(new_n714), .B2(new_n716), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n717), .A2(G190), .A3(G200), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT95), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n721), .A2(new_n722), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n720), .B1(G326), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(G283), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n298), .A2(new_n335), .A3(new_n709), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n298), .A2(new_n335), .A3(new_n715), .ZN(new_n731));
  INV_X1    g0531(.A(G303), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n729), .A2(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G179), .A2(G200), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT96), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n735), .A2(new_n207), .A3(G190), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n733), .B1(G329), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G294), .ZN(new_n738));
  OAI21_X1  g0538(.A(G20), .B1(new_n735), .B2(new_n366), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n728), .B(new_n737), .C1(new_n738), .C2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n736), .A2(G159), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT32), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n740), .A2(new_n511), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(G50), .B2(new_n727), .ZN(new_n745));
  OAI221_X1 g0545(.A(new_n255), .B1(new_n716), .B2(new_n202), .C1(new_n222), .C2(new_n711), .ZN(new_n746));
  INV_X1    g0546(.A(new_n718), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n746), .B1(G68), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n731), .A2(new_n532), .ZN(new_n749));
  INV_X1    g0549(.A(new_n730), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n749), .B1(G107), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n745), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n741), .B1(new_n743), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n708), .B1(new_n753), .B2(new_n699), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n694), .B1(new_n698), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n631), .B(new_n632), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n755), .B1(new_n756), .B2(new_n694), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT97), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(G396));
  NOR4_X1   g0559(.A1(new_n370), .A2(new_n371), .A3(new_n353), .A4(new_n627), .ZN(new_n760));
  INV_X1    g0560(.A(new_n372), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n367), .A2(new_n368), .B1(new_n353), .B2(new_n628), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n657), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n613), .A2(new_n628), .A3(new_n763), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n693), .B1(new_n767), .B2(new_n683), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(new_n683), .B2(new_n767), .ZN(new_n769));
  INV_X1    g0569(.A(G77), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n699), .A2(new_n695), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT98), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n694), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n699), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n712), .A2(G159), .ZN(new_n776));
  INV_X1    g0576(.A(G143), .ZN(new_n777));
  INV_X1    g0577(.A(G150), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n776), .B1(new_n777), .B2(new_n716), .C1(new_n778), .C2(new_n718), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n727), .B2(G137), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT34), .Z(new_n781));
  INV_X1    g0581(.A(new_n736), .ZN(new_n782));
  INV_X1    g0582(.A(G132), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n782), .A2(new_n783), .B1(new_n201), .B2(new_n731), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n740), .A2(new_n202), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n730), .A2(new_n220), .ZN(new_n786));
  NOR4_X1   g0586(.A1(new_n784), .A2(new_n785), .A3(new_n252), .A4(new_n786), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n532), .A2(new_n730), .B1(new_n731), .B2(new_n356), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(G311), .B2(new_n736), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n255), .B1(new_n712), .B2(G116), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n790), .B1(new_n729), .B2(new_n718), .C1(new_n738), .C2(new_n716), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n744), .B(new_n791), .C1(G303), .C2(new_n727), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n781), .A2(new_n787), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n774), .B1(new_n775), .B2(new_n793), .C1(new_n763), .C2(new_n696), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n769), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(G384));
  OR2_X1    g0596(.A1(new_n579), .A2(KEYINPUT35), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n579), .A2(KEYINPUT35), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n797), .A2(G116), .A3(new_n216), .A4(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT36), .Z(new_n800));
  OR3_X1    g0600(.A1(new_n222), .A2(new_n213), .A3(new_n399), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n201), .A2(G68), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n206), .B(G13), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT99), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n339), .A2(new_n805), .A3(new_n343), .ZN(new_n806));
  AND3_X1   g0606(.A1(new_n318), .A2(new_n319), .A3(new_n627), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n343), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n330), .A2(KEYINPUT14), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n334), .A2(new_n337), .A3(G169), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n809), .B(new_n810), .C1(new_n335), .C2(new_n334), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n806), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n339), .A2(KEYINPUT99), .A3(new_n343), .ZN(new_n814));
  INV_X1    g0614(.A(new_n807), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n760), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(new_n766), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT38), .ZN(new_n820));
  INV_X1    g0620(.A(new_n625), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT100), .ZN(new_n822));
  AOI21_X1  g0622(.A(KEYINPUT16), .B1(new_n420), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n396), .A2(new_n405), .A3(KEYINPUT100), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n423), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n821), .B1(new_n825), .B2(new_n375), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n419), .A2(new_n431), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n411), .B(KEYINPUT17), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n416), .B1(new_n825), .B2(new_n375), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n826), .A2(new_n830), .A3(new_n411), .ZN(new_n831));
  AND3_X1   g0631(.A1(new_n831), .A2(KEYINPUT101), .A3(KEYINPUT37), .ZN(new_n832));
  AOI21_X1  g0632(.A(KEYINPUT101), .B1(new_n831), .B2(KEYINPUT37), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n413), .A2(new_n416), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n413), .A2(new_n821), .ZN(new_n835));
  XOR2_X1   g0635(.A(KEYINPUT102), .B(KEYINPUT37), .Z(new_n836));
  NAND4_X1  g0636(.A1(new_n834), .A2(new_n835), .A3(new_n411), .A4(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR3_X1   g0638(.A1(new_n832), .A2(new_n833), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n820), .B1(new_n829), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n403), .A2(new_n404), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n290), .A2(G159), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n394), .B1(new_n255), .B2(G20), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n220), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n822), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n847), .A2(new_n421), .A3(new_n824), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n406), .A2(new_n281), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n375), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n411), .B1(new_n625), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n427), .A2(new_n850), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT37), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT101), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n831), .A2(KEYINPUT101), .A3(KEYINPUT37), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n855), .A2(new_n856), .A3(new_n837), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n857), .B(KEYINPUT38), .C1(new_n432), .C2(new_n826), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n840), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n819), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n616), .B2(new_n821), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT103), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n859), .A2(KEYINPUT39), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT39), .ZN(new_n864));
  XOR2_X1   g0664(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n865));
  NAND3_X1  g0665(.A1(new_n834), .A2(new_n835), .A3(new_n411), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(new_n836), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n835), .B1(new_n616), .B2(new_n828), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n865), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n858), .A2(new_n864), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n863), .A2(KEYINPUT104), .A3(new_n870), .ZN(new_n871));
  AOI211_X1 g0671(.A(KEYINPUT104), .B(new_n864), .C1(new_n840), .C2(new_n858), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n617), .A2(new_n628), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n871), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n616), .A2(new_n821), .ZN(new_n877));
  AOI211_X1 g0677(.A(KEYINPUT103), .B(new_n877), .C1(new_n819), .C2(new_n859), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n862), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n434), .B1(new_n658), .B2(new_n665), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n620), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n880), .B(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n763), .A2(new_n813), .A3(new_n816), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n677), .A2(KEYINPUT31), .A3(new_n627), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT31), .B1(new_n677), .B2(new_n627), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n884), .B1(new_n887), .B2(new_n667), .ZN(new_n888));
  INV_X1    g0688(.A(new_n858), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n417), .A2(new_n418), .A3(KEYINPUT78), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n429), .B1(new_n428), .B2(new_n430), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n828), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n826), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n894), .B2(new_n857), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n888), .B1(new_n889), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT40), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n858), .A2(new_n869), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT106), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT106), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n858), .A2(new_n901), .A3(new_n869), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n763), .A2(new_n816), .A3(new_n813), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n682), .A2(new_n903), .A3(KEYINPUT40), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n900), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n898), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n434), .A2(new_n682), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(new_n907), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n908), .A2(G330), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n883), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n206), .B2(new_n688), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n883), .A2(new_n910), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n804), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT107), .Z(G367));
  OAI211_X1 g0715(.A(new_n592), .B(new_n589), .C1(new_n590), .C2(new_n628), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n589), .B1(new_n487), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n627), .B1(new_n917), .B2(KEYINPUT108), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(KEYINPUT108), .B2(new_n917), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT42), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n610), .A2(new_n627), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n916), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n644), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n919), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n925), .A2(KEYINPUT109), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n925), .A2(KEYINPUT109), .B1(new_n920), .B2(new_n924), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n547), .A2(new_n628), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n567), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n605), .B2(new_n929), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n926), .A2(new_n927), .A3(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT110), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n926), .A2(new_n927), .A3(KEYINPUT110), .A4(new_n932), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n926), .A2(new_n927), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n931), .B(KEYINPUT43), .Z(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n642), .A2(new_n923), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n937), .A2(new_n942), .A3(new_n940), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n652), .B(KEYINPUT41), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n642), .A2(KEYINPUT113), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n644), .A2(new_n922), .A3(new_n645), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n948), .A2(KEYINPUT111), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT45), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(KEYINPUT111), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n950), .B1(new_n949), .B2(new_n951), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT44), .ZN(new_n956));
  OR3_X1    g0756(.A1(new_n646), .A2(new_n956), .A3(new_n922), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n956), .B1(new_n646), .B2(new_n922), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n957), .A2(KEYINPUT112), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(KEYINPUT112), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n947), .B1(new_n955), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n954), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n952), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n958), .A2(KEYINPUT112), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n958), .A2(KEYINPUT112), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n964), .B1(new_n965), .B2(new_n957), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n963), .B(new_n966), .C1(KEYINPUT113), .C2(new_n642), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n644), .B1(new_n637), .B2(new_n643), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(new_n633), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n970), .A2(new_n684), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n961), .A2(new_n967), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n946), .B1(new_n972), .B2(new_n685), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n944), .B(new_n945), .C1(new_n973), .C2(new_n692), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n700), .B1(new_n210), .B2(new_n346), .C1(new_n238), .C2(new_n702), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n693), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n697), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n252), .B1(new_n711), .B2(new_n729), .C1(new_n732), .C2(new_n716), .ZN(new_n978));
  INV_X1    g0778(.A(G317), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n782), .A2(new_n979), .B1(new_n511), .B2(new_n730), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n978), .B(new_n980), .C1(G294), .C2(new_n747), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n727), .A2(G311), .B1(G107), .B2(new_n739), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT46), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n731), .B2(new_n706), .ZN(new_n984));
  INV_X1    g0784(.A(new_n731), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n985), .A2(KEYINPUT46), .A3(G116), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n981), .A2(new_n982), .A3(new_n984), .A4(new_n986), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G58), .A2(new_n985), .B1(new_n750), .B2(new_n345), .ZN(new_n988));
  INV_X1    g0788(.A(G137), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n988), .B1(new_n989), .B2(new_n782), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n255), .B1(new_n711), .B2(new_n201), .C1(new_n778), .C2(new_n716), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G159), .B2(new_n747), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n739), .A2(G68), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n777), .C2(new_n726), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n987), .B1(new_n990), .B2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT47), .Z(new_n996));
  OAI221_X1 g0796(.A(new_n976), .B1(new_n977), .B2(new_n931), .C1(new_n996), .C2(new_n775), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n974), .A2(new_n997), .ZN(G387));
  NAND2_X1  g0798(.A1(new_n685), .A2(new_n969), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n970), .A2(new_n684), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n999), .A2(new_n687), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n653), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n705), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(G107), .B2(new_n210), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n235), .A2(new_n266), .ZN(new_n1005));
  AOI211_X1 g0805(.A(G45), .B(new_n1002), .C1(G68), .C2(G77), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n287), .A2(G50), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT50), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n702), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1004), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n693), .B1(new_n1010), .B2(new_n701), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n740), .A2(new_n729), .B1(new_n738), .B2(new_n731), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n712), .A2(G303), .ZN(new_n1013));
  INV_X1    g0813(.A(G311), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1013), .B1(new_n1014), .B2(new_n718), .C1(new_n979), .C2(new_n716), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n727), .B2(G322), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1012), .B1(new_n1016), .B2(KEYINPUT48), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT114), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(KEYINPUT48), .B2(new_n1016), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT49), .Z(new_n1020));
  AOI21_X1  g0820(.A(new_n255), .B1(new_n736), .B2(G326), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n706), .B2(new_n730), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n731), .A2(new_n222), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G97), .B2(new_n750), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n778), .B2(new_n782), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n255), .B1(new_n711), .B2(new_n220), .C1(new_n201), .C2(new_n716), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n288), .B2(new_n747), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n739), .A2(new_n347), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(new_n397), .C2(new_n726), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n1020), .A2(new_n1022), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1011), .B1(new_n1030), .B2(new_n699), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n637), .A2(new_n977), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n969), .A2(new_n692), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1001), .A2(new_n1033), .ZN(G393));
  NAND2_X1  g0834(.A1(new_n963), .A2(new_n966), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n999), .B1(new_n1035), .B2(new_n947), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n652), .B1(new_n1036), .B2(new_n967), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1035), .A2(new_n642), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1035), .A2(new_n642), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1039), .A2(new_n999), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n923), .A2(new_n697), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n252), .B1(new_n711), .B2(new_n738), .C1(new_n718), .C2(new_n732), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n782), .A2(new_n714), .B1(new_n729), .B2(new_n731), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1043), .B(new_n1044), .C1(G107), .C2(new_n750), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n726), .A2(new_n979), .B1(new_n1014), .B2(new_n716), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n739), .A2(G116), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1045), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n726), .A2(new_n778), .B1(new_n397), .B2(new_n716), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT51), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n739), .A2(G77), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n255), .B1(new_n711), .B2(new_n287), .C1(new_n718), .C2(new_n201), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G87), .B2(new_n750), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G143), .A2(new_n736), .B1(new_n985), .B2(G68), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n775), .B1(new_n1052), .B2(new_n1059), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n243), .A2(new_n702), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n701), .B1(G97), .B2(new_n649), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n694), .B(new_n1060), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1037), .A2(new_n1041), .B1(new_n1042), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT115), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1040), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1065), .B1(new_n1066), .B2(new_n1038), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1039), .A2(KEYINPUT115), .A3(new_n1040), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1067), .A2(new_n1068), .A3(new_n692), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1064), .A2(new_n1069), .ZN(G390));
  AOI21_X1  g0870(.A(new_n632), .B1(new_n887), .B2(new_n667), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n817), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1071), .A2(new_n763), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n819), .A2(new_n875), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n871), .B2(new_n873), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n900), .A2(new_n902), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n761), .A2(new_n762), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n760), .B1(new_n663), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n874), .B1(new_n1079), .B2(new_n817), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1074), .B1(new_n1076), .B2(new_n1081), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT104), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n859), .B2(KEYINPUT39), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n872), .B1(new_n1085), .B2(new_n870), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1083), .B(new_n1073), .C1(new_n1086), .C2(new_n1075), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1082), .A2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n881), .B(new_n620), .C1(new_n433), .C2(new_n683), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n817), .B1(new_n683), .B2(new_n764), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n1073), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n766), .A2(new_n818), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1090), .A2(new_n1073), .A3(new_n1079), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1089), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1088), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1082), .A2(new_n1095), .A3(new_n1087), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1097), .A2(new_n687), .A3(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1082), .A2(new_n692), .A3(new_n1087), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n693), .B1(new_n288), .B2(new_n772), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n749), .B(new_n786), .C1(G294), .C2(new_n736), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n727), .A2(G283), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n252), .B1(new_n711), .B2(new_n511), .C1(new_n706), .C2(new_n716), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G107), .B2(new_n747), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1102), .A2(new_n1055), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n727), .A2(G128), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n255), .B1(new_n730), .B2(new_n201), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n1108), .A2(KEYINPUT117), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n718), .A2(new_n989), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT54), .B(G143), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n716), .A2(new_n783), .B1(new_n711), .B2(new_n1111), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n1110), .B(new_n1112), .C1(new_n736), .C2(G125), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1108), .A2(KEYINPUT117), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1107), .A2(new_n1109), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  OR3_X1    g0915(.A1(new_n731), .A2(KEYINPUT53), .A3(new_n778), .ZN(new_n1116));
  OAI21_X1  g0916(.A(KEYINPUT53), .B1(new_n731), .B2(new_n778), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1116), .B(new_n1117), .C1(new_n740), .C2(new_n397), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1106), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1101), .B1(new_n1119), .B2(new_n699), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n1086), .B2(new_n696), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1099), .A2(new_n1100), .A3(new_n1121), .ZN(G378));
  NAND3_X1  g0922(.A1(new_n898), .A2(new_n905), .A3(G330), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n294), .A2(new_n625), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n308), .A2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n308), .A2(new_n1124), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  OR3_X1    g0928(.A1(new_n1125), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1128), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1123), .A2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n898), .A2(new_n905), .A3(G330), .A4(new_n1131), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n880), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n878), .B1(new_n1086), .B2(new_n875), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1137), .A2(new_n862), .A3(new_n1134), .A4(new_n1133), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n692), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n694), .B1(new_n201), .B2(new_n771), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n993), .B1(new_n726), .B2(new_n706), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT118), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n255), .A2(G41), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1144), .B1(new_n346), .B2(new_n711), .C1(new_n356), .C2(new_n716), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G97), .B2(new_n747), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n730), .A2(new_n202), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1023), .B(new_n1147), .C1(G283), .C2(new_n736), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1143), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT119), .Z(new_n1150));
  OR2_X1    g0950(.A1(new_n1150), .A2(KEYINPUT58), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(KEYINPUT58), .ZN(new_n1152));
  AOI211_X1 g0952(.A(G50), .B(new_n1144), .C1(new_n263), .C2(new_n264), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n727), .A2(G125), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n739), .A2(G150), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1111), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n985), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(G128), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n716), .A2(new_n1158), .B1(new_n711), .B2(new_n989), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G132), .B2(new_n747), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1154), .A2(new_n1155), .A3(new_n1157), .A4(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1161), .A2(KEYINPUT59), .ZN(new_n1162));
  AOI211_X1 g0962(.A(G33), .B(G41), .C1(new_n736), .C2(G124), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n397), .B2(new_n730), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1161), .A2(KEYINPUT59), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1153), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1151), .A2(new_n1152), .A3(new_n1167), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1141), .B1(new_n775), .B2(new_n1168), .C1(new_n1131), .C2(new_n696), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1140), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1089), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1098), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1176), .A2(KEYINPUT120), .A3(new_n687), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1139), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n1172), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(KEYINPUT120), .B1(new_n1176), .B2(new_n687), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1171), .B1(new_n1180), .B2(new_n1181), .ZN(G375));
  NAND3_X1  g0982(.A1(new_n1089), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n1183), .A2(KEYINPUT121), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1095), .A2(new_n946), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1183), .A2(KEYINPUT121), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n692), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n693), .B1(G68), .B2(new_n772), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n727), .A2(G294), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n718), .A2(new_n706), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n716), .A2(new_n729), .B1(new_n711), .B2(new_n356), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(new_n736), .C2(G303), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n985), .A2(G97), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1191), .A2(new_n1194), .A3(new_n1028), .A4(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n252), .B1(new_n730), .B2(new_n770), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT122), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n727), .A2(G132), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n739), .A2(G50), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n255), .B1(new_n711), .B2(new_n778), .C1(new_n989), .C2(new_n716), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n747), .B2(new_n1156), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1147), .B1(G128), .B2(new_n736), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n397), .B2(new_n731), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n1196), .A2(new_n1198), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT123), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n775), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1190), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1072), .B2(new_n696), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1189), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1187), .A2(new_n1213), .ZN(G381));
  NAND4_X1  g1014(.A1(new_n974), .A2(new_n997), .A3(new_n1064), .A4(new_n1069), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1001), .A2(new_n758), .A3(new_n1033), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1215), .A2(G384), .A3(G381), .A4(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT124), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(G375), .A2(G378), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(G407));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n626), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(G407), .A2(G213), .A3(new_n1221), .ZN(G409));
  NAND2_X1  g1022(.A1(new_n626), .A2(G213), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(G378), .B(new_n1171), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1225));
  INV_X1    g1025(.A(G378), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1178), .A2(new_n946), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1226), .B1(new_n1170), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1224), .B1(new_n1225), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT60), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1184), .B(new_n1186), .C1(new_n1230), .C2(new_n1095), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1183), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n652), .B1(new_n1232), .B2(KEYINPUT60), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(G384), .A3(new_n1213), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(G384), .B1(new_n1234), .B2(new_n1213), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1229), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT63), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(G2897), .B(new_n1224), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1237), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1224), .A2(G2897), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n1235), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1229), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1229), .A2(KEYINPUT63), .A3(new_n1238), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(G393), .A2(G396), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1216), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1215), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n974), .A2(new_n997), .B1(new_n1064), .B2(new_n1069), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1250), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G387), .A2(G390), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1250), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n1215), .A3(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT61), .B1(new_n1253), .B2(new_n1256), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1241), .A2(new_n1247), .A3(new_n1248), .A4(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT62), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1229), .A2(new_n1259), .A3(new_n1238), .ZN(new_n1260));
  XOR2_X1   g1060(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n1229), .B2(new_n1246), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1259), .B1(new_n1229), .B2(new_n1238), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(new_n1260), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(new_n1251), .A2(new_n1252), .A3(new_n1250), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1255), .B1(new_n1254), .B2(new_n1215), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT126), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT126), .B1(new_n1253), .B2(new_n1256), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1258), .B1(new_n1264), .B2(new_n1270), .ZN(G405));
  NOR2_X1   g1071(.A1(new_n1238), .A2(KEYINPUT127), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1238), .A2(KEYINPUT127), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1225), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(new_n1226), .B2(G375), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1267), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1272), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1253), .A2(KEYINPUT126), .A3(new_n1256), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1273), .A2(new_n1276), .A3(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1276), .B1(new_n1273), .B2(new_n1280), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(G402));
endmodule


