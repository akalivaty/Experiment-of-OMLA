//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND3_X1  g0005(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  AOI21_X1  g0007(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G1), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n210), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT0), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n217), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n214), .B(new_n220), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  INV_X1    g0043(.A(G107), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G97), .ZN(new_n245));
  INV_X1    g0045(.A(G97), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G107), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n243), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  AOI21_X1  g0053(.A(G1), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  AND3_X1   g0056(.A1(new_n254), .A2(new_n256), .A3(G274), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT67), .B(G1), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G41), .A2(G45), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(G1), .A2(G13), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n258), .A2(new_n260), .B1(new_n261), .B2(new_n255), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n257), .B1(new_n262), .B2(G226), .ZN(new_n263));
  OR2_X1    g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G223), .A3(G1698), .ZN(new_n267));
  AND2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G77), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n266), .A2(G222), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(KEYINPUT68), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n274), .A2(new_n267), .A3(KEYINPUT68), .A4(new_n271), .ZN(new_n276));
  INV_X1    g0076(.A(new_n208), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n277), .A2(new_n206), .B1(G33), .B2(G41), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n263), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  OR2_X1    g0080(.A1(new_n280), .A2(G179), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT69), .ZN(new_n284));
  INV_X1    g0084(.A(G58), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n284), .B1(new_n285), .B2(KEYINPUT70), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT8), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n285), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT69), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n284), .B(KEYINPUT8), .C1(new_n285), .C2(KEYINPUT70), .ZN(new_n291));
  AND3_X1   g0091(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n210), .A2(G33), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n283), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n277), .A2(new_n206), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n215), .A2(KEYINPUT67), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT67), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G1), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n298), .A2(new_n300), .A3(G13), .A4(G20), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(G50), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n296), .B1(G20), .B2(new_n258), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n302), .B1(new_n303), .B2(G50), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n297), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n280), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n281), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n308), .A2(KEYINPUT71), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(KEYINPUT71), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G33), .ZN(new_n312));
  INV_X1    g0112(.A(G87), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G226), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G1698), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(G223), .B2(G1698), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n315), .B1(new_n318), .B2(new_n270), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n278), .ZN(new_n320));
  INV_X1    g0120(.A(G274), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n261), .B2(new_n255), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n254), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n298), .A2(new_n300), .ZN(new_n324));
  OAI211_X1 g0124(.A(G232), .B(new_n256), .C1(new_n324), .C2(new_n259), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n320), .A2(KEYINPUT76), .A3(new_n323), .A4(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n257), .B1(new_n319), .B2(new_n278), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT76), .B1(new_n328), .B2(new_n325), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n306), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(G223), .A2(G1698), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n316), .B2(G1698), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n314), .B1(new_n332), .B2(new_n266), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n255), .B1(new_n207), .B2(new_n208), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n323), .B(new_n325), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(G179), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n330), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n303), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n301), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n292), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT7), .B1(new_n270), .B2(new_n210), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n264), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n265), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(G68), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n282), .A2(G159), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AND3_X1   g0149(.A1(KEYINPUT75), .A2(G58), .A3(G68), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT75), .B1(G58), .B2(G68), .ZN(new_n351));
  OR3_X1    g0151(.A1(new_n350), .A2(new_n351), .A3(new_n201), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n349), .B1(new_n352), .B2(G20), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT16), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n347), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G68), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n264), .A2(new_n210), .A3(new_n265), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT7), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n356), .B1(new_n359), .B2(new_n345), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n350), .A2(new_n351), .A3(new_n201), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n348), .B1(new_n361), .B2(new_n210), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT16), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n355), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n343), .B1(new_n364), .B2(new_n296), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT18), .B1(new_n338), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT17), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n354), .B1(new_n347), .B2(new_n353), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n360), .A2(new_n362), .A3(KEYINPUT16), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n296), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n343), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n335), .A2(G190), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT76), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n335), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n326), .ZN(new_n376));
  INV_X1    g0176(.A(G200), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n373), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n367), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n336), .B1(new_n376), .B2(new_n306), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT18), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n372), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(G200), .B1(new_n375), .B2(new_n326), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n365), .B(KEYINPUT17), .C1(new_n383), .C2(new_n373), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n366), .A2(new_n379), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  XOR2_X1   g0186(.A(KEYINPUT8), .B(G58), .Z(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(new_n282), .B1(G20), .B2(G77), .ZN(new_n388));
  XNOR2_X1  g0188(.A(KEYINPUT15), .B(G87), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n388), .B1(new_n293), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G77), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n390), .A2(new_n296), .B1(new_n391), .B2(new_n341), .ZN(new_n392));
  INV_X1    g0192(.A(new_n303), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n392), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n262), .A2(G244), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n266), .A2(G238), .A3(G1698), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n266), .A2(G232), .A3(new_n273), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n396), .B(new_n397), .C1(new_n244), .C2(new_n266), .ZN(new_n398));
  AOI211_X1 g0198(.A(new_n257), .B(new_n395), .C1(new_n398), .C2(new_n278), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n394), .B1(new_n399), .B2(G190), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(new_n377), .B2(new_n399), .ZN(new_n401));
  OR2_X1    g0201(.A1(new_n399), .A2(G169), .ZN(new_n402));
  INV_X1    g0202(.A(G179), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n394), .A3(new_n404), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n280), .A2(G200), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT9), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n305), .A2(new_n408), .ZN(new_n409));
  OAI211_X1 g0209(.A(G190), .B(new_n263), .C1(new_n275), .C2(new_n279), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n297), .A2(KEYINPUT9), .A3(new_n304), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n407), .A2(new_n409), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  OR2_X1    g0212(.A1(new_n412), .A2(KEYINPUT10), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(KEYINPUT10), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n311), .A2(new_n386), .A3(new_n406), .A4(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n257), .B1(new_n262), .B2(G238), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n316), .A2(new_n273), .ZN(new_n418));
  INV_X1    g0218(.A(G232), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G1698), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n418), .B(new_n420), .C1(new_n268), .C2(new_n269), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT72), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G33), .A2(G97), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n278), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n422), .B1(new_n421), .B2(new_n423), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n417), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT13), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT73), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT13), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n417), .B(new_n430), .C1(new_n425), .C2(new_n426), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n428), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n427), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(G169), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT14), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT14), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n432), .A2(new_n436), .A3(G169), .A4(new_n433), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n428), .A2(G179), .A3(new_n431), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT74), .B1(new_n301), .B2(G68), .ZN(new_n440));
  XOR2_X1   g0240(.A(new_n440), .B(KEYINPUT12), .Z(new_n441));
  INV_X1    g0241(.A(new_n282), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(new_n202), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n293), .A2(new_n391), .B1(new_n210), .B2(G68), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n296), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT11), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n441), .B(new_n446), .C1(new_n356), .C2(new_n393), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n439), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G190), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n449), .B1(new_n427), .B2(KEYINPUT13), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n447), .B1(new_n450), .B2(new_n431), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n432), .A2(G200), .A3(new_n433), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n416), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n298), .A2(new_n300), .A3(G45), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT5), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G41), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(G270), .B(new_n256), .C1(new_n456), .C2(new_n460), .ZN(new_n461));
  XNOR2_X1  g0261(.A(KEYINPUT5), .B(G41), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n322), .A2(new_n258), .A3(new_n462), .A4(G45), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT80), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT80), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n461), .A2(new_n466), .A3(new_n463), .ZN(new_n467));
  AND2_X1   g0267(.A1(KEYINPUT81), .A2(G303), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT81), .A2(G303), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n264), .B(new_n265), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(G264), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n471));
  OAI211_X1 g0271(.A(G257), .B(new_n273), .C1(new_n268), .C2(new_n269), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n278), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n465), .A2(new_n467), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(KEYINPUT82), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT82), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n464), .A2(KEYINPUT80), .B1(new_n278), .B2(new_n473), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n477), .B1(new_n478), .B2(new_n467), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT20), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G283), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n482), .B(new_n210), .C1(G33), .C2(new_n246), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT83), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n483), .B(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n296), .B1(new_n210), .B2(G116), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n481), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g0287(.A(new_n483), .B(KEYINPUT83), .ZN(new_n488));
  INV_X1    g0288(.A(G116), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n209), .A2(new_n295), .B1(G20), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n490), .A3(KEYINPUT20), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n301), .A2(G116), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n298), .A2(new_n300), .A3(G33), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n301), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(new_n296), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n493), .B1(new_n496), .B2(G116), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n306), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT21), .B1(new_n480), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n475), .A2(KEYINPUT82), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n478), .A2(new_n477), .A3(new_n467), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n498), .A2(new_n500), .A3(KEYINPUT21), .A4(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n478), .A2(G179), .A3(new_n467), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n492), .A2(new_n497), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n499), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n480), .A2(G200), .ZN(new_n509));
  INV_X1    g0309(.A(new_n505), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n509), .B(new_n510), .C1(new_n449), .C2(new_n480), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n244), .A2(KEYINPUT23), .A3(G20), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT23), .B1(new_n244), .B2(G20), .ZN(new_n513));
  OAI22_X1  g0313(.A1(new_n512), .A2(new_n513), .B1(new_n489), .B2(new_n293), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n210), .B(G87), .C1(new_n268), .C2(new_n269), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT22), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT22), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n266), .A2(new_n517), .A3(new_n210), .A4(G87), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n514), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n519), .A2(KEYINPUT24), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n296), .B1(new_n519), .B2(KEYINPUT24), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT77), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n495), .B2(new_n296), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n277), .A2(new_n206), .A3(new_n295), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n525), .A2(KEYINPUT77), .A3(new_n301), .A4(new_n494), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n526), .A3(G107), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT85), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n301), .B2(G107), .ZN(new_n529));
  XNOR2_X1  g0329(.A(KEYINPUT84), .B(KEYINPUT25), .ZN(new_n530));
  OR2_X1    g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n341), .A2(KEYINPUT85), .A3(new_n244), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n532), .A2(new_n529), .A3(new_n530), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n527), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n522), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(G257), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n536));
  OAI211_X1 g0336(.A(G250), .B(new_n273), .C1(new_n268), .C2(new_n269), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G294), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n278), .ZN(new_n540));
  OAI211_X1 g0340(.A(G264), .B(new_n256), .C1(new_n456), .C2(new_n460), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n463), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT86), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT86), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n540), .A2(new_n544), .A3(new_n463), .A4(new_n541), .ZN(new_n545));
  AOI21_X1  g0345(.A(G190), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n542), .A2(new_n377), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n535), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n543), .A2(G169), .A3(new_n545), .ZN(new_n549));
  OR2_X1    g0349(.A1(new_n542), .A2(new_n403), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n533), .A2(new_n531), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n552), .B(new_n527), .C1(new_n521), .C2(new_n520), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n548), .A2(new_n554), .ZN(new_n555));
  OR2_X1    g0355(.A1(KEYINPUT79), .A2(G87), .ZN(new_n556));
  NAND2_X1  g0356(.A1(KEYINPUT79), .A2(G87), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n556), .A2(new_n246), .A3(new_n244), .A4(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT19), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n210), .B1(new_n423), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n266), .A2(new_n210), .A3(G68), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n559), .B1(new_n293), .B2(new_n246), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n564), .A2(new_n296), .B1(new_n341), .B2(new_n389), .ZN(new_n565));
  INV_X1    g0365(.A(new_n389), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n524), .A2(new_n526), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n456), .A2(G250), .A3(new_n256), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n322), .A2(G45), .A3(new_n258), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(G238), .B(new_n273), .C1(new_n268), .C2(new_n269), .ZN(new_n572));
  OAI211_X1 g0372(.A(G244), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G33), .A2(G116), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n278), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n306), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n571), .A2(new_n576), .A3(new_n403), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n568), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n577), .A2(G200), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n524), .A2(new_n526), .A3(G87), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n571), .A2(new_n576), .A3(G190), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n581), .A2(new_n565), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(G250), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n482), .ZN(new_n587));
  OAI211_X1 g0387(.A(G244), .B(new_n273), .C1(new_n268), .C2(new_n269), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT78), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n587), .B1(KEYINPUT4), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT4), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n588), .A2(KEYINPUT78), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n334), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(G257), .B(new_n256), .C1(new_n456), .C2(new_n460), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n463), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n306), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n589), .A2(KEYINPUT4), .ZN(new_n597));
  INV_X1    g0397(.A(new_n587), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n592), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n595), .B1(new_n599), .B2(new_n278), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n403), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT6), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n245), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g0403(.A(G97), .B(G107), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n603), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  OAI22_X1  g0405(.A1(new_n605), .A2(new_n210), .B1(new_n391), .B2(new_n442), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n244), .B1(new_n359), .B2(new_n345), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n296), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n524), .A2(new_n526), .A3(G97), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n341), .A2(new_n246), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n596), .A2(new_n601), .A3(new_n611), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n600), .A2(G190), .ZN(new_n614));
  OAI21_X1  g0414(.A(G200), .B1(new_n593), .B2(new_n595), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n585), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n555), .A2(new_n617), .ZN(new_n618));
  AND4_X1   g0418(.A1(new_n455), .A2(new_n508), .A3(new_n511), .A4(new_n618), .ZN(G372));
  INV_X1    g0419(.A(KEYINPUT90), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n415), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT90), .B1(new_n413), .B2(new_n414), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n372), .A2(new_n380), .A3(new_n381), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n381), .B1(new_n372), .B2(new_n380), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT88), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT88), .B1(new_n366), .B2(new_n382), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n405), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n439), .A2(new_n447), .B1(new_n630), .B2(new_n453), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n379), .A2(new_n384), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n623), .B1(KEYINPUT89), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT89), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n635), .B(new_n629), .C1(new_n631), .C2(new_n632), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n634), .A2(new_n636), .B1(new_n310), .B2(new_n309), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n596), .A2(new_n601), .A3(new_n611), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n585), .A2(new_n638), .A3(KEYINPUT26), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n580), .A2(new_n584), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n640), .B1(new_n641), .B2(new_n612), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n639), .A2(new_n642), .A3(KEYINPUT87), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT87), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n644), .B(new_n640), .C1(new_n641), .C2(new_n612), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n643), .A2(new_n580), .A3(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n548), .A2(new_n612), .A3(new_n585), .A4(new_n616), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n647), .B1(new_n508), .B2(new_n554), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n455), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n637), .A2(new_n650), .ZN(G369));
  AND2_X1   g0451(.A1(new_n210), .A2(G13), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n258), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT91), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n657));
  INV_X1    g0457(.A(G213), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G343), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n505), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n508), .A2(new_n511), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n508), .B2(new_n664), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n548), .B(new_n554), .C1(new_n535), .C2(new_n662), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n663), .A2(new_n551), .A3(new_n553), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n554), .A2(new_n663), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n662), .B1(new_n499), .B2(new_n507), .ZN(new_n675));
  XOR2_X1   g0475(.A(new_n675), .B(KEYINPUT92), .Z(new_n676));
  AOI21_X1  g0476(.A(new_n674), .B1(new_n676), .B2(new_n670), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n673), .A2(new_n677), .ZN(G399));
  INV_X1    g0478(.A(new_n218), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(G41), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n558), .A2(G116), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G1), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n212), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  INV_X1    g0485(.A(G330), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT94), .ZN(new_n687));
  INV_X1    g0487(.A(new_n467), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n473), .A2(new_n278), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n466), .B1(new_n461), .B2(new_n463), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AND4_X1   g0491(.A1(new_n541), .A2(new_n571), .A3(new_n540), .A4(new_n576), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n691), .A2(G179), .A3(new_n692), .A4(new_n600), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n687), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n692), .A2(new_n600), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(new_n504), .A3(KEYINPUT94), .A4(KEYINPUT30), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n692), .A2(new_n600), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n694), .B1(new_n699), .B2(new_n503), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n542), .A2(new_n577), .A3(new_n403), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n599), .A2(new_n278), .ZN(new_n702));
  INV_X1    g0502(.A(new_n595), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n500), .A2(new_n701), .A3(new_n501), .A4(new_n704), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n698), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n663), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT31), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n700), .A2(new_n705), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT93), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n700), .A2(new_n705), .A3(KEYINPUT93), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(new_n698), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n662), .A2(new_n709), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n708), .A2(new_n709), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n618), .A2(new_n508), .A3(new_n511), .A4(new_n662), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n686), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT21), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n721), .A2(new_n554), .A3(new_n506), .A4(new_n502), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT95), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n502), .A2(new_n506), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(KEYINPUT95), .A3(new_n721), .A4(new_n554), .ZN(new_n726));
  INV_X1    g0526(.A(new_n617), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n724), .A2(new_n726), .A3(new_n548), .A4(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n580), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n639), .B2(new_n642), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n663), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT29), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n662), .B1(new_n646), .B2(new_n648), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT29), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n718), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n685), .B1(new_n736), .B2(G1), .ZN(G364));
  AOI21_X1  g0537(.A(new_n215), .B1(new_n652), .B2(G45), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n680), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n218), .A2(new_n266), .ZN(new_n741));
  INV_X1    g0541(.A(G355), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n741), .A2(new_n742), .B1(G116), .B2(new_n218), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n679), .A2(new_n266), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n745), .B1(new_n253), .B2(new_n213), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n243), .A2(new_n253), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n743), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n209), .B1(G20), .B2(new_n306), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n740), .B1(new_n748), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n210), .A2(new_n403), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n757), .A2(new_n377), .A3(G190), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n757), .A2(new_n449), .A3(new_n377), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n759), .A2(new_n356), .B1(new_n761), .B2(new_n202), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G190), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n756), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n270), .B(new_n762), .C1(G77), .C2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n210), .A2(G179), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n767), .A2(new_n449), .A3(G200), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G107), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n767), .A2(new_n763), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G159), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n770), .B1(new_n773), .B2(KEYINPUT32), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n767), .A2(G190), .A3(G200), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(new_n556), .B2(new_n557), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n449), .A2(G200), .ZN(new_n778));
  AND3_X1   g0578(.A1(new_n756), .A2(KEYINPUT96), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(KEYINPUT96), .B1(new_n756), .B2(new_n778), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G58), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n778), .A2(new_n403), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n246), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(KEYINPUT32), .B2(new_n773), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n766), .A2(new_n777), .A3(new_n783), .A4(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n760), .B(KEYINPUT97), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n791), .A2(G326), .B1(G294), .B2(new_n785), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(KEYINPUT98), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n782), .A2(G322), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n772), .A2(G329), .ZN(new_n796));
  XOR2_X1   g0596(.A(KEYINPUT33), .B(G317), .Z(new_n797));
  OAI21_X1  g0597(.A(new_n796), .B1(new_n759), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G311), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n270), .B1(new_n764), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G283), .ZN(new_n801));
  INV_X1    g0601(.A(G303), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n801), .A2(new_n768), .B1(new_n775), .B2(new_n802), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n798), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT98), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n795), .B(new_n804), .C1(new_n792), .C2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n789), .B1(new_n794), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n755), .B1(new_n807), .B2(new_n749), .ZN(new_n808));
  INV_X1    g0608(.A(new_n752), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n666), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n740), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n667), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n666), .A2(G330), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT99), .Z(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G396));
  NOR2_X1   g0616(.A1(new_n405), .A2(new_n663), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n663), .A2(new_n394), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n401), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n817), .B1(new_n819), .B2(new_n405), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n733), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n662), .B(new_n820), .C1(new_n646), .C2(new_n648), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n718), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n811), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n718), .B1(new_n822), .B2(new_n823), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n825), .B1(KEYINPUT100), .B2(new_n826), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n826), .A2(KEYINPUT100), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n760), .A2(G137), .B1(G159), .B2(new_n765), .ZN(new_n830));
  INV_X1    g0630(.A(G143), .ZN(new_n831));
  INV_X1    g0631(.A(G150), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n830), .B1(new_n831), .B2(new_n781), .C1(new_n832), .C2(new_n759), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT34), .Z(new_n834));
  NOR2_X1   g0634(.A1(new_n786), .A2(new_n285), .ZN(new_n835));
  INV_X1    g0635(.A(G132), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n266), .B1(new_n771), .B2(new_n836), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n202), .A2(new_n775), .B1(new_n768), .B2(new_n356), .ZN(new_n838));
  NOR4_X1   g0638(.A1(new_n834), .A2(new_n835), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n266), .B(new_n787), .C1(G116), .C2(new_n765), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n759), .A2(new_n801), .B1(new_n771), .B2(new_n799), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(G303), .B2(new_n760), .ZN(new_n842));
  INV_X1    g0642(.A(new_n775), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n843), .A2(G107), .B1(new_n769), .B2(G87), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n782), .A2(G294), .ZN(new_n845));
  AND4_X1   g0645(.A1(new_n840), .A2(new_n842), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n749), .B1(new_n839), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n749), .A2(new_n750), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n811), .B1(new_n848), .B2(new_n391), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n847), .B(new_n849), .C1(new_n820), .C2(new_n751), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n829), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(G384));
  INV_X1    g0652(.A(new_n605), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n853), .A2(KEYINPUT35), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(KEYINPUT35), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n854), .A2(G116), .A3(new_n211), .A4(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT36), .Z(new_n857));
  OR4_X1    g0657(.A1(new_n391), .A2(new_n350), .A3(new_n351), .A4(new_n212), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n202), .A2(G68), .ZN(new_n859));
  AOI211_X1 g0659(.A(G13), .B(new_n258), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n817), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n823), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n525), .B1(new_n355), .B2(new_n363), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n661), .B1(new_n864), .B2(new_n343), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n385), .A2(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n330), .B(new_n337), .C1(new_n864), .C2(new_n343), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n370), .B(new_n371), .C1(new_n383), .C2(new_n373), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n868), .A2(new_n869), .A3(new_n865), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT37), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n868), .A2(new_n869), .A3(new_n865), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT38), .B1(new_n867), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n867), .A2(new_n874), .A3(KEYINPUT38), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n663), .A2(new_n447), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n448), .A2(new_n453), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n453), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n447), .B(new_n663), .C1(new_n881), .C2(new_n439), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n863), .A2(new_n878), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n660), .B1(new_n627), .B2(new_n628), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT101), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n867), .A2(new_n874), .A3(KEYINPUT38), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT39), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n889), .A2(new_n875), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n871), .A2(new_n873), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n869), .A2(new_n367), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n377), .B1(new_n327), .B2(new_n329), .ZN(new_n894));
  INV_X1    g0694(.A(new_n373), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT17), .B1(new_n896), .B2(new_n365), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT103), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n626), .B1(new_n624), .B2(new_n625), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n366), .A2(KEYINPUT88), .A3(new_n382), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT103), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n379), .A2(new_n384), .A3(new_n901), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n898), .A2(new_n899), .A3(new_n900), .A4(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n892), .B1(new_n903), .B2(new_n866), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n877), .B1(new_n904), .B2(KEYINPUT38), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n891), .B1(new_n905), .B2(new_n890), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n448), .A2(new_n663), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT102), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n907), .B(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n884), .A2(KEYINPUT101), .A3(new_n885), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n888), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n732), .A2(new_n455), .A3(new_n735), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n637), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n912), .B(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT31), .B1(new_n707), .B2(new_n663), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n709), .B(new_n662), .C1(new_n698), .C2(new_n706), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n821), .B1(new_n918), .B2(new_n717), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n905), .A2(new_n919), .A3(KEYINPUT40), .A4(new_n883), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT40), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n710), .B1(new_n695), .B2(new_n697), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n709), .B1(new_n922), .B2(new_n662), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n717), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(new_n883), .A3(new_n820), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n889), .A2(new_n875), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n921), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n920), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n455), .A2(new_n925), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n929), .A2(new_n930), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n931), .A2(G330), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n915), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n258), .B2(new_n652), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n915), .A2(new_n933), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n861), .B1(new_n935), .B2(new_n936), .ZN(G367));
  OAI221_X1 g0737(.A(new_n753), .B1(new_n218), .B2(new_n389), .C1(new_n745), .C2(new_n239), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT106), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n811), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n939), .B2(new_n938), .ZN(new_n941));
  INV_X1    g0741(.A(G159), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n759), .A2(new_n942), .B1(new_n764), .B2(new_n202), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n270), .B(new_n943), .C1(G137), .C2(new_n772), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n768), .A2(new_n391), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n786), .A2(new_n356), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n945), .B(new_n946), .C1(G58), .C2(new_n843), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n791), .A2(G143), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n782), .A2(G150), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n944), .A2(new_n947), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n843), .A2(G116), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT46), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n468), .A2(new_n469), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n952), .B1(new_n953), .B2(new_n781), .C1(new_n799), .C2(new_n790), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n758), .A2(G294), .B1(G317), .B2(new_n772), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n266), .B1(new_n765), .B2(G283), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n769), .A2(G97), .B1(new_n785), .B2(G107), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n950), .B1(new_n954), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT47), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n941), .B1(new_n960), .B2(new_n749), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n662), .B1(new_n565), .B2(new_n582), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n729), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n641), .B2(new_n962), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(new_n809), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n670), .B1(new_n666), .B2(G330), .ZN(new_n967));
  OR3_X1    g0767(.A1(new_n672), .A2(new_n676), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n676), .B1(new_n672), .B2(new_n967), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n736), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT45), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n676), .A2(new_n670), .ZN(new_n975));
  INV_X1    g0775(.A(new_n674), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n616), .B(new_n612), .C1(new_n613), .C2(new_n662), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n638), .A2(new_n663), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n974), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n677), .A2(KEYINPUT45), .A3(new_n980), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n977), .A2(KEYINPUT44), .A3(new_n981), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT44), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n677), .B2(new_n980), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n984), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n672), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n984), .A2(new_n673), .A3(new_n988), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n973), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n992), .A2(new_n736), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n680), .B(KEYINPUT41), .Z(new_n994));
  OAI21_X1  g0794(.A(KEYINPUT105), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n994), .B1(new_n992), .B2(new_n736), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT105), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n739), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n672), .A2(new_n980), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT104), .Z(new_n1001));
  NOR2_X1   g0801(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n676), .A2(new_n670), .A3(new_n980), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1004), .A2(KEYINPUT42), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n612), .B1(new_n978), .B2(new_n554), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n1004), .A2(KEYINPUT42), .B1(new_n662), .B2(new_n1006), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n1005), .A2(new_n1007), .B1(KEYINPUT43), .B2(new_n964), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1003), .B(new_n1008), .Z(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n966), .B1(new_n999), .B2(new_n1010), .ZN(G387));
  INV_X1    g0811(.A(new_n973), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n971), .A2(new_n972), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(new_n680), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n266), .B1(new_n764), .B2(new_n356), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n786), .A2(new_n389), .B1(new_n768), .B2(new_n246), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(G159), .C2(new_n760), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n843), .A2(G77), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n832), .B2(new_n771), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT108), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n758), .A2(new_n339), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n782), .A2(G50), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1017), .A2(new_n1020), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n764), .A2(new_n953), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(new_n782), .B2(G317), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1026), .A2(KEYINPUT109), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(KEYINPUT109), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n791), .A2(G322), .B1(G311), .B2(new_n758), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT48), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(G294), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n786), .A2(new_n801), .B1(new_n775), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1032), .A2(KEYINPUT49), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n266), .B1(new_n772), .B2(G326), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(new_n489), .C2(new_n768), .ZN(new_n1038));
  AOI21_X1  g0838(.A(KEYINPUT49), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1023), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n749), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n682), .B(KEYINPUT107), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n253), .B1(new_n356), .B2(new_n391), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n387), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1044), .A2(G50), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT50), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1042), .B(new_n1047), .C1(new_n1046), .C2(new_n1045), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1048), .B(new_n744), .C1(new_n236), .C2(new_n253), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(G107), .B2(new_n218), .C1(new_n682), .C2(new_n741), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n811), .B1(new_n1050), .B2(new_n753), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1041), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n671), .B2(new_n752), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n970), .B2(new_n739), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1014), .A2(new_n1054), .ZN(G393));
  AND2_X1   g0855(.A1(new_n992), .A2(new_n680), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n990), .A2(new_n991), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n1012), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n990), .A2(new_n739), .A3(new_n991), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT112), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n745), .A2(new_n250), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n753), .B1(new_n246), .B2(new_n218), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n740), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT110), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n782), .A2(G159), .B1(G150), .B2(new_n760), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT51), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n758), .A2(G50), .B1(new_n387), .B2(new_n765), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT111), .Z(new_n1069));
  OAI221_X1 g0869(.A(new_n266), .B1(new_n771), .B2(new_n831), .C1(new_n313), .C2(new_n768), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n786), .A2(new_n391), .B1(new_n775), .B2(new_n356), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n1067), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n782), .A2(G311), .B1(G317), .B2(new_n760), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT52), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G294), .A2(new_n765), .B1(new_n772), .B2(G322), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1075), .B(new_n270), .C1(new_n953), .C2(new_n759), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n770), .B1(new_n801), .B2(new_n775), .C1(new_n786), .C2(new_n489), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n1074), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1072), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1065), .B1(new_n1079), .B2(new_n749), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n981), .A2(new_n752), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n1060), .A2(new_n1061), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1061), .B1(new_n1060), .B2(new_n1082), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1059), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(G390));
  INV_X1    g0887(.A(new_n848), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n740), .B1(new_n1088), .B2(new_n339), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n759), .A2(new_n244), .B1(new_n761), .B2(new_n801), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G97), .B2(new_n765), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n270), .B1(new_n771), .B2(new_n1033), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G68), .B2(new_n769), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n843), .A2(G87), .B1(new_n785), .B2(G77), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n782), .A2(G116), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1091), .A2(new_n1093), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n758), .A2(G137), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT54), .B(G143), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1097), .B1(new_n942), .B2(new_n786), .C1(new_n764), .C2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT114), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n270), .B1(new_n772), .B2(G125), .ZN(new_n1101));
  INV_X1    g0901(.A(G128), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1101), .B1(new_n761), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(G50), .B2(new_n769), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n775), .A2(new_n832), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT53), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1104), .B(new_n1106), .C1(new_n836), .C2(new_n781), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1096), .B1(new_n1100), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1089), .B1(new_n1108), .B2(new_n749), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n906), .B2(new_n751), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n909), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n819), .A2(new_n405), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n817), .B1(new_n731), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n883), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1111), .B(new_n905), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n909), .B1(new_n883), .B2(new_n863), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1115), .B1(new_n906), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n925), .A2(G330), .A3(new_n820), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1118), .A2(new_n1114), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n718), .A2(new_n820), .A3(new_n883), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1115), .B(new_n1121), .C1(new_n906), .C2(new_n1116), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n633), .A2(KEYINPUT89), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1124), .B(new_n636), .C1(new_n621), .C2(new_n622), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n455), .A2(G330), .A3(new_n925), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n913), .A2(new_n1125), .A3(new_n311), .A4(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n883), .B1(new_n718), .B2(new_n820), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n863), .B1(new_n1128), .B2(new_n1119), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1118), .A2(new_n1114), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1121), .A2(new_n1130), .A3(new_n1113), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1127), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT113), .Z(new_n1133));
  INV_X1    g0933(.A(new_n1123), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1120), .A2(new_n1132), .A3(new_n1122), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n680), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1110), .B1(new_n738), .B2(new_n1123), .C1(new_n1135), .C2(new_n1137), .ZN(G378));
  INV_X1    g0938(.A(KEYINPUT57), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT118), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1127), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1136), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n920), .A2(new_n928), .A3(G330), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n308), .B1(new_n621), .B2(new_n622), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n661), .A2(new_n305), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n308), .B(new_n1145), .C1(new_n621), .C2(new_n622), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT116), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1143), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT38), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n379), .A2(new_n901), .A3(new_n384), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n901), .B1(new_n379), .B2(new_n384), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n865), .B1(new_n629), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1157), .B1(new_n1161), .B2(new_n892), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n921), .B1(new_n1162), .B2(new_n877), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n926), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n686), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(KEYINPUT116), .B1(new_n1165), .B2(new_n928), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n920), .A2(new_n928), .A3(KEYINPUT116), .A4(G330), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1150), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n912), .B(new_n1156), .C1(new_n1166), .C2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1143), .A2(new_n1155), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1174), .A2(new_n1167), .A3(new_n1170), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n912), .B1(new_n1175), .B2(new_n1156), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1142), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1140), .B1(new_n1136), .B2(new_n1141), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1139), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1178), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1156), .B1(new_n1166), .B2(new_n1171), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n912), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n1172), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1180), .A2(KEYINPUT57), .A3(new_n1184), .A4(new_n1142), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1179), .A2(new_n1185), .A3(new_n680), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n738), .B1(new_n1183), .B2(new_n1172), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT117), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n740), .B1(new_n1088), .B2(G50), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT115), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n758), .A2(G97), .B1(G283), .B2(new_n772), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n389), .B2(new_n764), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n782), .B2(G107), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n270), .A2(new_n252), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1195), .B(new_n946), .C1(G116), .C2(new_n760), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n769), .A2(G58), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1194), .A2(new_n1196), .A3(new_n1018), .A4(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT58), .ZN(new_n1199));
  AOI21_X1  g0999(.A(G50), .B1(new_n312), .B2(new_n252), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1198), .A2(new_n1199), .B1(new_n1195), .B2(new_n1200), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n786), .A2(new_n832), .B1(new_n775), .B2(new_n1098), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n758), .A2(G132), .B1(new_n760), .B2(G125), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n765), .A2(G137), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1202), .B(new_n1205), .C1(G128), .C2(new_n782), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(KEYINPUT59), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n769), .A2(G159), .ZN(new_n1209));
  AOI211_X1 g1009(.A(G33), .B(G41), .C1(new_n772), .C2(G124), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1207), .A2(KEYINPUT59), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1201), .B1(new_n1199), .B2(new_n1198), .C1(new_n1211), .C2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1191), .B1(new_n1213), .B2(new_n749), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n1154), .B2(new_n751), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1188), .A2(new_n1189), .A3(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1215), .ZN(new_n1217));
  OAI21_X1  g1017(.A(KEYINPUT117), .B1(new_n1187), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1186), .A2(new_n1219), .ZN(G375));
  INV_X1    g1020(.A(new_n1129), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1131), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n739), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n811), .B1(new_n848), .B2(new_n356), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n761), .A2(new_n1033), .B1(new_n771), .B2(new_n802), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G116), .B2(new_n758), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n266), .B(new_n945), .C1(G107), .C2(new_n765), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(G97), .A2(new_n843), .B1(new_n785), .B2(new_n566), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n782), .A2(G283), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n266), .B1(new_n771), .B2(new_n1102), .C1(new_n832), .C2(new_n764), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1197), .B1(new_n942), .B2(new_n775), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1231), .B(new_n1232), .C1(G50), .C2(new_n785), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(KEYINPUT119), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n759), .A2(new_n1098), .B1(new_n761), .B2(new_n836), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n782), .B2(G137), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT119), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1237), .B1(new_n1233), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1230), .B1(new_n1235), .B2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1240), .A2(KEYINPUT120), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(KEYINPUT120), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n749), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1224), .B1(new_n1241), .B2(new_n1243), .C1(new_n883), .C2(new_n751), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1223), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1129), .A2(new_n1127), .A3(new_n1131), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n994), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1246), .B1(new_n1133), .B2(new_n1249), .ZN(G381));
  INV_X1    g1050(.A(G378), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1251), .A2(new_n1186), .A3(new_n1219), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1086), .B(new_n966), .C1(new_n999), .C2(new_n1010), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1014), .A2(new_n815), .A3(new_n1054), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n851), .ZN(new_n1256));
  OR4_X1    g1056(.A1(G381), .A2(new_n1252), .A3(new_n1253), .A4(new_n1256), .ZN(G407));
  OAI211_X1 g1057(.A(G407), .B(G213), .C1(G343), .C2(new_n1252), .ZN(G409));
  NOR2_X1   g1058(.A1(new_n658), .A2(G343), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1177), .A2(new_n994), .A3(new_n1178), .ZN(new_n1261));
  OAI21_X1  g1061(.A(KEYINPUT121), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT121), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1183), .A2(new_n1263), .A3(new_n1172), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1262), .A2(new_n739), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1215), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1261), .B1(new_n1266), .B2(KEYINPUT122), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT122), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1265), .A2(new_n1268), .A3(new_n1215), .ZN(new_n1269));
  AOI21_X1  g1069(.A(G378), .B1(new_n1267), .B2(new_n1269), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1186), .A2(new_n1219), .A3(G378), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1260), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1259), .A2(G2897), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1132), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT60), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1247), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1274), .A2(new_n1276), .A3(KEYINPUT123), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT123), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n680), .B1(new_n1247), .B2(new_n1275), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(new_n1278), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n851), .B1(new_n1281), .B2(new_n1245), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1277), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1284), .A2(G384), .A3(new_n1246), .ZN(new_n1285));
  AOI211_X1 g1085(.A(KEYINPUT124), .B(new_n1273), .C1(new_n1282), .C2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1282), .A2(new_n1285), .A3(KEYINPUT124), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1287), .A2(G2897), .A3(new_n1259), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT124), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1282), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1285), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1289), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1286), .B1(new_n1288), .B2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT61), .B1(new_n1272), .B2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1186), .A2(new_n1219), .A3(G378), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1269), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1268), .B1(new_n1265), .B2(new_n1215), .ZN(new_n1297));
  NOR3_X1   g1097(.A1(new_n1296), .A2(new_n1297), .A3(new_n1261), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1295), .B1(new_n1298), .B2(G378), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT62), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1299), .A2(new_n1300), .A3(new_n1260), .A4(new_n1301), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1260), .B(new_n1301), .C1(new_n1270), .C2(new_n1271), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(KEYINPUT62), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1294), .A2(new_n1302), .A3(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT125), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n815), .B1(new_n1014), .B2(new_n1054), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1255), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1306), .B1(new_n1255), .B2(new_n1307), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1253), .A2(new_n1309), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n996), .A2(new_n997), .ZN(new_n1311));
  AOI211_X1 g1111(.A(KEYINPUT105), .B(new_n994), .C1(new_n992), .C2(new_n736), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n738), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(new_n1313), .A2(new_n1009), .B1(new_n965), .B2(new_n961), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1314), .A2(new_n1086), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1308), .B1(new_n1310), .B2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(G387), .A2(G390), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1308), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1317), .A2(new_n1253), .A3(new_n1318), .A4(new_n1309), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1316), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1305), .A2(new_n1320), .ZN(new_n1321));
  AND2_X1   g1121(.A1(new_n1316), .A2(new_n1319), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT63), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1303), .A2(new_n1323), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1299), .A2(KEYINPUT63), .A3(new_n1260), .A4(new_n1301), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1322), .A2(new_n1324), .A3(new_n1294), .A4(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1321), .A2(new_n1326), .ZN(G405));
  NAND2_X1  g1127(.A1(G375), .A2(new_n1251), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1328), .B1(new_n1271), .B2(KEYINPUT126), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT126), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(G375), .A2(new_n1330), .A3(new_n1251), .ZN(new_n1331));
  NOR3_X1   g1131(.A1(new_n1290), .A2(new_n1291), .A3(KEYINPUT127), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT127), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1301), .A2(new_n1333), .ZN(new_n1334));
  OAI211_X1 g1134(.A(new_n1329), .B(new_n1331), .C1(new_n1332), .C2(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(G378), .B1(new_n1186), .B2(new_n1219), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1336), .B1(new_n1330), .B2(new_n1295), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1331), .ZN(new_n1338));
  OAI22_X1  g1138(.A1(new_n1337), .A2(new_n1338), .B1(new_n1333), .B2(new_n1301), .ZN(new_n1339));
  AND3_X1   g1139(.A1(new_n1320), .A2(new_n1335), .A3(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1320), .B1(new_n1335), .B2(new_n1339), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1340), .A2(new_n1341), .ZN(G402));
endmodule


