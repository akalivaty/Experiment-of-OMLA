//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1248,
    new_n1249, new_n1250, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n206), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n206), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  NOR2_X1   g0017(.A1(G58), .A2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT64), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n220), .A2(G50), .A3(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n214), .A2(new_n217), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n213), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  XOR2_X1   g0045(.A(KEYINPUT8), .B(G58), .Z(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n225), .A2(G1), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G13), .A3(G20), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n224), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n249), .A2(new_n255), .B1(new_n252), .B2(new_n247), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT16), .ZN(new_n258));
  INV_X1    g0058(.A(G68), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT80), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n264));
  AOI21_X1  g0064(.A(G20), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n260), .B1(new_n265), .B2(KEYINPUT7), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT7), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  OAI211_X1 g0068(.A(KEYINPUT80), .B(new_n267), .C1(new_n268), .C2(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT81), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT81), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n262), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(new_n264), .A3(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n267), .A2(G20), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n259), .B1(new_n270), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G58), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(new_n259), .ZN(new_n280));
  OAI21_X1  g0080(.A(G20), .B1(new_n280), .B2(new_n218), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G159), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n258), .B1(new_n278), .B2(new_n284), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n253), .A2(new_n224), .ZN(new_n286));
  INV_X1    g0086(.A(new_n276), .ZN(new_n287));
  OAI22_X1  g0087(.A1(new_n265), .A2(KEYINPUT7), .B1(new_n287), .B2(new_n268), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n284), .B1(new_n288), .B2(G68), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n286), .B1(new_n289), .B2(KEYINPUT16), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n257), .B1(new_n285), .B2(new_n290), .ZN(new_n291));
  AND2_X1   g0091(.A1(G33), .A2(G41), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT65), .B1(new_n292), .B2(new_n224), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n250), .B1(G41), .B2(G45), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G41), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT65), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n296), .A2(new_n297), .A3(G1), .A4(G13), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n293), .A2(new_n295), .A3(G274), .A4(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n293), .A2(G232), .A3(new_n294), .A4(new_n298), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT83), .ZN(new_n301));
  AND3_X1   g0101(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(new_n299), .B2(new_n300), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n296), .A2(G1), .A3(G13), .ZN(new_n304));
  OR2_X1    g0104(.A1(G223), .A2(G1698), .ZN(new_n305));
  INV_X1    g0105(.A(G226), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G1698), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n262), .A2(new_n305), .A3(new_n264), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(G33), .A2(G87), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n304), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NOR3_X1   g0110(.A1(new_n302), .A2(new_n303), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n299), .A2(new_n300), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT83), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT82), .ZN(new_n316));
  NOR2_X1   g0116(.A1(G223), .A2(G1698), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(new_n306), .B2(G1698), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n318), .A2(new_n268), .B1(G33), .B2(G87), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n316), .B1(new_n319), .B2(new_n304), .ZN(new_n320));
  INV_X1    g0120(.A(G179), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n310), .A2(KEYINPUT82), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n311), .A2(G169), .B1(new_n315), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT18), .B1(new_n291), .B2(new_n324), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n313), .B(new_n314), .C1(new_n304), .C2(new_n319), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n302), .A2(new_n303), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n326), .A2(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT18), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n288), .A2(G68), .ZN(new_n332));
  INV_X1    g0132(.A(new_n284), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(KEYINPUT16), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n254), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n266), .A2(new_n269), .B1(new_n276), .B2(new_n275), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n333), .B1(new_n336), .B2(new_n259), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n335), .B1(new_n258), .B2(new_n337), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n330), .B(new_n331), .C1(new_n338), .C2(new_n257), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n325), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G190), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n320), .A2(new_n341), .A3(new_n322), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n311), .A2(G200), .B1(new_n315), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n261), .A2(G33), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n225), .B1(new_n271), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT80), .B1(new_n345), .B2(new_n267), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n265), .A2(new_n260), .A3(KEYINPUT7), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n277), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n284), .B1(new_n348), .B2(G68), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n290), .B1(new_n349), .B2(KEYINPUT16), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT17), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n256), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n343), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT84), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n343), .A2(new_n350), .A3(new_n256), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT17), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n343), .A2(new_n350), .A3(KEYINPUT84), .A4(new_n353), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT85), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AND4_X1   g0162(.A1(KEYINPUT84), .A2(new_n343), .A3(new_n350), .A4(new_n353), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n351), .B1(new_n291), .B2(new_n343), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n365), .A2(KEYINPUT85), .A3(new_n356), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n340), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n293), .A2(new_n298), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(G244), .A3(new_n294), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n369), .A2(new_n299), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n268), .A2(G238), .A3(G1698), .ZN(new_n371));
  INV_X1    g0171(.A(G1698), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n268), .A2(G232), .A3(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n371), .B(new_n373), .C1(new_n203), .C2(new_n268), .ZN(new_n374));
  INV_X1    g0174(.A(new_n304), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n370), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n321), .ZN(new_n379));
  INV_X1    g0179(.A(G77), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n248), .A2(new_n380), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n255), .A2(new_n381), .B1(new_n380), .B2(new_n252), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT15), .B(G87), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n225), .A2(G33), .ZN(new_n384));
  OR3_X1    g0184(.A1(new_n383), .A2(KEYINPUT69), .A3(new_n384), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n246), .A2(new_n282), .B1(G20), .B2(G77), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT69), .B1(new_n383), .B2(new_n384), .ZN(new_n387));
  AND3_X1   g0187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n382), .B1(new_n388), .B2(new_n286), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n377), .A2(new_n327), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n379), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AOI22_X1  g0191(.A1(G200), .A2(new_n377), .B1(new_n389), .B2(KEYINPUT70), .ZN(new_n392));
  OR2_X1    g0192(.A1(new_n389), .A2(KEYINPUT70), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(KEYINPUT71), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n378), .A2(G190), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT71), .B1(new_n392), .B2(new_n393), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n391), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G150), .ZN(new_n399));
  INV_X1    g0199(.A(new_n282), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n247), .A2(new_n384), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G50), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n225), .B1(new_n218), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n254), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n250), .A2(G20), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT67), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(G50), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT67), .B1(new_n248), .B2(new_n402), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n255), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(G50), .B2(new_n251), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n410), .A2(KEYINPUT68), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(KEYINPUT68), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n404), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(G222), .A2(G1698), .ZN(new_n414));
  XOR2_X1   g0214(.A(KEYINPUT66), .B(G223), .Z(new_n415));
  AOI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(G1698), .ZN(new_n416));
  INV_X1    g0216(.A(new_n268), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n375), .B1(new_n268), .B2(G77), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n368), .A2(new_n294), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n299), .B1(new_n421), .B2(new_n306), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n321), .ZN(new_n424));
  OAI221_X1 g0224(.A(new_n299), .B1(new_n421), .B2(new_n306), .C1(new_n418), .C2(new_n419), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n327), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n413), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n413), .A2(KEYINPUT9), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT9), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n404), .C1(new_n411), .C2(new_n412), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT10), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n423), .A2(G190), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n425), .A2(G200), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n433), .A2(new_n434), .A3(KEYINPUT72), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n431), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n432), .B1(new_n431), .B2(new_n435), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n427), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n398), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n252), .A2(new_n259), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT12), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n282), .A2(G50), .B1(G20), .B2(new_n259), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(new_n380), .B2(new_n384), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(KEYINPUT11), .A3(new_n254), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n255), .A2(G68), .A3(new_n405), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n441), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT11), .B1(new_n443), .B2(new_n254), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  XOR2_X1   g0248(.A(new_n448), .B(KEYINPUT77), .Z(new_n449));
  NAND4_X1  g0249(.A1(new_n293), .A2(G238), .A3(new_n294), .A4(new_n298), .ZN(new_n450));
  NOR2_X1   g0250(.A1(G226), .A2(G1698), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n451), .B1(new_n231), .B2(G1698), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n452), .A2(new_n268), .B1(G33), .B2(G97), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n299), .B(new_n450), .C1(new_n453), .C2(new_n304), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT76), .B1(new_n454), .B2(KEYINPUT13), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(KEYINPUT13), .B2(new_n454), .ZN(new_n456));
  INV_X1    g0256(.A(new_n454), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT13), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(KEYINPUT76), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n449), .B1(G190), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT73), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n457), .A2(new_n462), .A3(new_n458), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT73), .B1(new_n454), .B2(KEYINPUT13), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT74), .B1(new_n457), .B2(new_n458), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT74), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n454), .A2(new_n467), .A3(KEYINPUT13), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n465), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT75), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n469), .A2(new_n470), .A3(G200), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n470), .B1(new_n469), .B2(G200), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n461), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g0273(.A1(KEYINPUT78), .A2(G169), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n463), .A2(new_n464), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n466), .A2(new_n468), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT14), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n460), .A2(G179), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT79), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT14), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n469), .A2(new_n482), .A3(new_n474), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n460), .A2(KEYINPUT79), .A3(G179), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n478), .A2(new_n481), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n449), .ZN(new_n486));
  AND4_X1   g0286(.A1(new_n367), .A2(new_n439), .A3(new_n473), .A4(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT5), .ZN(new_n488));
  INV_X1    g0288(.A(G41), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(KEYINPUT5), .A2(G41), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(new_n250), .A3(G45), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n368), .A2(G257), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n250), .A2(G45), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n490), .B2(new_n491), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n496), .A2(G274), .A3(new_n293), .A4(new_n298), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n268), .A2(G250), .A3(G1698), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G283), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n262), .A2(new_n264), .A3(G244), .A4(new_n372), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n499), .B(new_n500), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT86), .B1(new_n502), .B2(new_n501), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n502), .A2(KEYINPUT86), .A3(new_n501), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n498), .B(new_n321), .C1(new_n507), .C2(new_n304), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT87), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n506), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(new_n504), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n375), .B1(new_n512), .B2(new_n503), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n513), .A2(KEYINPUT87), .A3(new_n321), .A4(new_n498), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n336), .A2(new_n203), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G97), .A2(G107), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT6), .B1(new_n204), .B2(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n203), .A2(KEYINPUT6), .A3(G97), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI22_X1  g0320(.A1(new_n520), .A2(new_n225), .B1(new_n380), .B2(new_n400), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n254), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n251), .A2(G97), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n250), .A2(G33), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n286), .A2(new_n251), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n523), .B1(new_n526), .B2(G97), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n498), .B1(new_n507), .B2(new_n304), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n522), .A2(new_n527), .B1(new_n528), .B2(new_n327), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n515), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n522), .A2(new_n527), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n528), .A2(G200), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n498), .B(G190), .C1(new_n507), .C2(new_n304), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n268), .A2(new_n225), .A3(G87), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT22), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT22), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n268), .A2(new_n537), .A3(new_n225), .A4(G87), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT24), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G116), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n541), .A2(G20), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT23), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n225), .B2(G107), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n539), .A2(new_n540), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n540), .B1(new_n539), .B2(new_n546), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n254), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n268), .A2(G257), .A3(G1698), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n268), .A2(G250), .A3(new_n372), .ZN(new_n552));
  NAND2_X1  g0352(.A1(G33), .A2(G294), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n375), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n368), .A2(G264), .A3(new_n493), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n557), .A2(G190), .A3(new_n497), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n252), .A2(KEYINPUT25), .A3(new_n203), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT25), .B1(new_n252), .B2(new_n203), .ZN(new_n561));
  OAI22_X1  g0361(.A1(new_n560), .A2(new_n561), .B1(new_n525), .B2(new_n203), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n555), .A2(new_n497), .A3(new_n556), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G200), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n550), .A2(new_n558), .A3(new_n563), .A4(new_n565), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n530), .A2(new_n534), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT90), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n268), .A2(G244), .A3(G1698), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n262), .A2(new_n264), .A3(G238), .A4(new_n372), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n541), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n375), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n495), .A2(KEYINPUT88), .A3(G250), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT88), .ZN(new_n574));
  AOI21_X1  g0374(.A(G274), .B1(new_n574), .B2(G250), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n573), .B1(new_n495), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n368), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n572), .A2(new_n321), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n225), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(G87), .B2(new_n204), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n262), .A2(new_n264), .A3(new_n225), .A4(G68), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT19), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n384), .B2(new_n202), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n254), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT89), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n525), .B2(new_n383), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n383), .A2(new_n252), .ZN(new_n589));
  INV_X1    g0389(.A(new_n383), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n255), .A2(KEYINPUT89), .A3(new_n590), .A4(new_n524), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n586), .A2(new_n588), .A3(new_n589), .A4(new_n591), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n571), .A2(new_n375), .B1(new_n368), .B2(new_n576), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n578), .B(new_n592), .C1(G169), .C2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n572), .A2(G190), .A3(new_n577), .ZN(new_n596));
  INV_X1    g0396(.A(G200), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n572), .B2(new_n577), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n585), .A2(new_n254), .B1(new_n252), .B2(new_n383), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n526), .A2(G87), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR3_X1   g0401(.A1(new_n596), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n568), .B1(new_n595), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n550), .A2(new_n563), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n564), .A2(new_n327), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n555), .A2(new_n321), .A3(new_n497), .A4(new_n556), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n593), .A2(G190), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(new_n599), .A3(new_n600), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n594), .B(KEYINPUT90), .C1(new_n610), .C2(new_n598), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n603), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n493), .A2(G270), .A3(new_n293), .A4(new_n298), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n613), .A2(new_n497), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n268), .A2(G264), .A3(G1698), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n268), .A2(G257), .A3(new_n372), .ZN(new_n616));
  INV_X1    g0416(.A(G303), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n615), .B(new_n616), .C1(new_n617), .C2(new_n268), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n375), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G200), .ZN(new_n621));
  INV_X1    g0421(.A(G116), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n252), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n525), .B2(new_n622), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n500), .B(new_n225), .C1(G33), .C2(new_n202), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n622), .A2(G20), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n254), .A2(KEYINPUT91), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT91), .B1(new_n254), .B2(new_n626), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT20), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI211_X1 g0431(.A(KEYINPUT20), .B(new_n625), .C1(new_n627), .C2(new_n628), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n624), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n621), .B(new_n633), .C1(new_n341), .C2(new_n620), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT21), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n618), .A2(new_n375), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n613), .A2(new_n497), .ZN(new_n637));
  OAI21_X1  g0437(.A(G169), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n635), .B1(new_n638), .B2(new_n633), .ZN(new_n639));
  INV_X1    g0439(.A(new_n633), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n640), .A2(KEYINPUT21), .A3(G169), .A4(new_n620), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n637), .B1(new_n375), .B2(new_n618), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n640), .A2(G179), .A3(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n634), .A2(new_n639), .A3(new_n641), .A4(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n612), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n487), .A2(new_n567), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g0446(.A(new_n646), .B(KEYINPUT92), .Z(G372));
  INV_X1    g0447(.A(KEYINPUT93), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n368), .A2(new_n648), .A3(new_n576), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n648), .B1(new_n368), .B2(new_n576), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n572), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n327), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n588), .A2(new_n591), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n653), .A2(new_n599), .B1(new_n593), .B2(new_n321), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n530), .A2(new_n534), .A3(new_n566), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n596), .A2(new_n601), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n651), .A2(G200), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n641), .A2(new_n639), .A3(new_n643), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n605), .A2(new_n606), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n550), .B2(new_n563), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n659), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n655), .B1(new_n656), .B2(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n603), .A2(new_n515), .A3(new_n529), .A4(new_n611), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n657), .A2(new_n658), .B1(new_n652), .B2(new_n654), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n515), .A2(new_n666), .A3(new_n529), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  MUX2_X1   g0468(.A(new_n665), .B(new_n667), .S(new_n668), .Z(new_n669));
  OAI21_X1  g0469(.A(new_n487), .B1(new_n664), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n427), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n325), .A2(new_n339), .ZN(new_n672));
  INV_X1    g0472(.A(new_n391), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n473), .A2(new_n673), .B1(new_n449), .B2(new_n485), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT85), .B1(new_n365), .B2(new_n356), .ZN(new_n675));
  AND4_X1   g0475(.A1(KEYINPUT85), .A2(new_n356), .A3(new_n358), .A4(new_n359), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n672), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n436), .A2(new_n437), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n671), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n670), .A2(new_n681), .ZN(G369));
  NAND3_X1  g0482(.A1(new_n250), .A2(new_n225), .A3(G13), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(KEYINPUT27), .ZN(new_n684));
  XOR2_X1   g0484(.A(new_n684), .B(KEYINPUT94), .Z(new_n685));
  INV_X1    g0485(.A(G213), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n683), .B2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G343), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(new_n633), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n660), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n644), .B2(new_n692), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G330), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n566), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n691), .B1(new_n550), .B2(new_n563), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n608), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n662), .A2(new_n691), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n696), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n660), .A2(new_n691), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n701), .B1(new_n700), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n704), .A2(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n215), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G1), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n222), .B2(new_n711), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT28), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n645), .A2(new_n567), .A3(new_n691), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n642), .A2(new_n557), .A3(G179), .A4(new_n593), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n717), .B1(new_n718), .B2(new_n528), .ZN(new_n719));
  INV_X1    g0519(.A(new_n528), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n620), .A2(new_n321), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n593), .A2(new_n556), .A3(new_n555), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n720), .A2(new_n721), .A3(KEYINPUT30), .A4(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(G179), .B1(new_n614), .B2(new_n619), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n528), .A2(new_n564), .A3(new_n724), .A4(new_n651), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n719), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n690), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT31), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n726), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n716), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G330), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT96), .ZN(new_n734));
  AND3_X1   g0534(.A1(new_n641), .A2(new_n639), .A3(new_n643), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n608), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n522), .A2(new_n533), .A3(new_n527), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n515), .A2(new_n529), .B1(new_n737), .B2(new_n532), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n736), .A2(new_n738), .A3(new_n566), .A4(new_n659), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n665), .A2(new_n668), .ZN(new_n740));
  AND4_X1   g0540(.A1(KEYINPUT26), .A2(new_n515), .A3(new_n666), .A4(new_n529), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n739), .B(new_n655), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n734), .B1(new_n742), .B2(new_n691), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n741), .B1(new_n668), .B2(new_n665), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n734), .B(new_n691), .C1(new_n744), .C2(new_n664), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(KEYINPUT29), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n691), .B1(new_n669), .B2(new_n664), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(KEYINPUT95), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT29), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT95), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n751), .B(new_n691), .C1(new_n669), .C2(new_n664), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n733), .B1(new_n747), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n715), .B1(new_n754), .B2(G1), .ZN(G364));
  INV_X1    g0555(.A(G13), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n250), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n710), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n268), .A2(new_n215), .ZN(new_n761));
  INV_X1    g0561(.A(G355), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n761), .A2(new_n762), .B1(G116), .B2(new_n215), .ZN(new_n763));
  INV_X1    g0563(.A(G45), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n241), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n709), .A2(new_n268), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(new_n223), .B2(new_n764), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n763), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(G20), .B1(KEYINPUT97), .B2(G169), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(KEYINPUT97), .A2(G169), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n224), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G20), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n760), .B1(new_n769), .B2(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n341), .A2(G179), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n225), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n225), .A2(new_n321), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n341), .ZN(new_n785));
  AOI22_X1  g0585(.A1(G97), .A2(new_n782), .B1(new_n785), .B2(G50), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G190), .A2(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n268), .B1(new_n788), .B2(new_n380), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n783), .A2(G190), .A3(new_n597), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n789), .B1(G58), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n225), .A2(G179), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n793), .A2(G190), .A3(G200), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G87), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n793), .A2(new_n787), .ZN(new_n797));
  INV_X1    g0597(.A(G159), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT32), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n786), .A2(new_n792), .A3(new_n796), .A4(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n784), .A2(G190), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n793), .A2(new_n341), .A3(G200), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n803), .A2(G68), .B1(new_n805), .B2(G107), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n800), .B2(new_n799), .ZN(new_n807));
  INV_X1    g0607(.A(G317), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(KEYINPUT33), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n808), .A2(KEYINPUT33), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n803), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G294), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n811), .B1(new_n812), .B2(new_n781), .C1(new_n617), .C2(new_n794), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n785), .A2(G326), .B1(new_n805), .B2(G283), .ZN(new_n814));
  INV_X1    g0614(.A(new_n797), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n791), .A2(G322), .B1(new_n815), .B2(G329), .ZN(new_n816));
  INV_X1    g0616(.A(new_n788), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n268), .B1(new_n817), .B2(G311), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n814), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n802), .A2(new_n807), .B1(new_n813), .B2(new_n819), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n820), .A2(KEYINPUT98), .ZN(new_n821));
  INV_X1    g0621(.A(new_n773), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n820), .B2(KEYINPUT98), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n779), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n776), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n694), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n760), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n695), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n694), .A2(G330), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n826), .B1(new_n828), .B2(new_n829), .ZN(G396));
  NAND2_X1  g0630(.A1(new_n690), .A2(new_n389), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n396), .B2(new_n397), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n391), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n391), .A2(new_n690), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n749), .A2(new_n752), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n834), .B1(new_n832), .B2(new_n391), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n838), .B(new_n691), .C1(new_n669), .C2(new_n664), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n733), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT100), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n837), .A2(new_n733), .A3(new_n839), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n842), .A2(new_n827), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n773), .A2(new_n774), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n827), .B1(new_n846), .B2(new_n380), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G116), .A2(new_n817), .B1(new_n815), .B2(G311), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n848), .B(new_n417), .C1(new_n812), .C2(new_n790), .ZN(new_n849));
  INV_X1    g0649(.A(new_n785), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n850), .A2(new_n617), .B1(new_n794), .B2(new_n203), .ZN(new_n851));
  INV_X1    g0651(.A(new_n803), .ZN(new_n852));
  INV_X1    g0652(.A(G283), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n852), .A2(new_n853), .B1(new_n202), .B2(new_n781), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n805), .A2(G87), .ZN(new_n855));
  NOR4_X1   g0655(.A1(new_n849), .A2(new_n851), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n791), .A2(G143), .B1(new_n817), .B2(G159), .ZN(new_n857));
  INV_X1    g0657(.A(G137), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n857), .B1(new_n852), .B2(new_n399), .C1(new_n858), .C2(new_n850), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT34), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n805), .A2(G68), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n402), .B2(new_n794), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n862), .A2(KEYINPUT99), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n862), .A2(KEYINPUT99), .ZN(new_n864));
  INV_X1    g0664(.A(G132), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n268), .B1(new_n797), .B2(new_n865), .C1(new_n781), .C2(new_n279), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n856), .B1(new_n860), .B2(new_n867), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n847), .B1(new_n822), .B2(new_n868), .C1(new_n838), .C2(new_n775), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n845), .A2(new_n869), .ZN(G384));
  NOR2_X1   g0670(.A1(new_n757), .A2(new_n250), .ZN(new_n871));
  INV_X1    g0671(.A(G330), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT40), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n289), .A2(KEYINPUT16), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n256), .B1(new_n335), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n330), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n688), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n357), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n330), .B1(new_n338), .B2(new_n257), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n877), .B1(new_n338), .B2(new_n257), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n881), .A2(new_n882), .A3(new_n357), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n367), .B2(new_n878), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n672), .B1(new_n675), .B2(new_n676), .ZN(new_n888));
  INV_X1    g0688(.A(new_n878), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n885), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n891), .A2(new_n887), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n886), .A2(new_n887), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n449), .A2(new_n690), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n486), .A2(new_n473), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n485), .A2(new_n449), .A3(new_n690), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n836), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT105), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n727), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n726), .A2(KEYINPUT105), .A3(new_n690), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(new_n728), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(new_n730), .A3(new_n716), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n873), .B1(new_n893), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n897), .A2(KEYINPUT40), .A3(new_n902), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n892), .B1(new_n367), .B2(new_n878), .ZN(new_n906));
  XOR2_X1   g0706(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n907));
  NAND3_X1  g0707(.A1(new_n881), .A2(new_n882), .A3(new_n357), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n909), .A2(new_n884), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n882), .B1(new_n360), .B2(new_n672), .ZN(new_n911));
  OAI211_X1 g0711(.A(KEYINPUT103), .B(new_n907), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n909), .A2(new_n884), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n340), .B1(new_n365), .B2(new_n356), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n914), .B1(new_n915), .B2(new_n882), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT103), .B1(new_n916), .B2(new_n907), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n906), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n905), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n904), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT106), .Z(new_n921));
  AND2_X1   g0721(.A1(new_n487), .A2(new_n902), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n872), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n922), .B2(new_n921), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n891), .B1(new_n888), .B2(new_n889), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n906), .B1(new_n925), .B2(KEYINPUT38), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n839), .A2(new_n835), .B1(new_n895), .B2(new_n896), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n672), .A2(new_n877), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT101), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT101), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n932), .B(new_n929), .C1(new_n926), .C2(new_n927), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT104), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n913), .A2(new_n917), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT39), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n906), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n935), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n926), .A2(KEYINPUT39), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT103), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n912), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT39), .B1(new_n890), .B2(new_n892), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n944), .A2(new_n945), .A3(KEYINPUT104), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n939), .A2(new_n940), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n485), .A2(new_n449), .A3(new_n691), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n934), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n747), .A2(new_n487), .A3(new_n753), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n681), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n951), .B(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n871), .B1(new_n924), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n954), .B2(new_n924), .ZN(new_n956));
  INV_X1    g0756(.A(new_n520), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n957), .A2(KEYINPUT35), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(KEYINPUT35), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n958), .A2(G116), .A3(new_n226), .A4(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT36), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n222), .A2(new_n380), .A3(new_n280), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n259), .A2(G50), .ZN(new_n963));
  OAI211_X1 g0763(.A(G1), .B(new_n756), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n956), .A2(new_n961), .A3(new_n964), .ZN(G367));
  NOR2_X1   g0765(.A1(new_n237), .A2(new_n767), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n777), .B1(new_n215), .B2(new_n383), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n760), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n852), .A2(new_n798), .B1(new_n804), .B2(new_n380), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(G58), .B2(new_n795), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n790), .A2(new_n399), .B1(new_n788), .B2(new_n402), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n417), .B(new_n971), .C1(G137), .C2(new_n815), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n781), .A2(new_n259), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(G143), .B2(new_n785), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n970), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(G311), .A2(new_n785), .B1(new_n791), .B2(G303), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT113), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n417), .B1(new_n797), .B2(new_n808), .C1(new_n202), .C2(new_n804), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(KEYINPUT114), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(KEYINPUT114), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n977), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n782), .A2(G107), .B1(new_n817), .B2(G283), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n803), .A2(G294), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT46), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n794), .B2(new_n622), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n795), .A2(KEYINPUT46), .A3(G116), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n983), .A2(new_n984), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n975), .B1(new_n982), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT47), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n968), .B1(new_n990), .B2(new_n773), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n690), .A2(new_n601), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT107), .Z(new_n993));
  NAND3_X1  g0793(.A1(new_n993), .A2(new_n654), .A3(new_n652), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT108), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n666), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n994), .B(new_n995), .C1(new_n997), .C2(new_n993), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n991), .B1(new_n1000), .B2(new_n825), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n738), .B1(new_n531), .B2(new_n691), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n515), .A2(new_n529), .A3(new_n690), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1005), .A2(new_n706), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT45), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT111), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT44), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1004), .B(new_n707), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1008), .B(new_n1009), .C1(new_n707), .C2(new_n1004), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1007), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(new_n704), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n703), .B(new_n705), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n695), .A2(KEYINPUT112), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1015), .B(new_n1016), .Z(new_n1017));
  NAND3_X1  g0817(.A1(new_n1014), .A2(new_n754), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n754), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n710), .B(KEYINPUT41), .Z(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n759), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n534), .A2(new_n662), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n690), .B1(new_n1023), .B2(new_n530), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n700), .A2(new_n702), .A3(new_n705), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT42), .B1(new_n1025), .B2(new_n1004), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1025), .A2(new_n1004), .A3(KEYINPUT42), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1024), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1000), .A2(KEYINPUT43), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1000), .A2(KEYINPUT43), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT110), .Z(new_n1033));
  NAND2_X1  g0833(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT109), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n704), .A2(new_n1005), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1033), .A2(new_n1037), .A3(new_n1035), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1001), .B1(new_n1022), .B2(new_n1041), .ZN(G387));
  NAND2_X1  g0842(.A1(new_n1017), .A2(new_n759), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n761), .A2(new_n712), .B1(G107), .B2(new_n215), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n234), .A2(new_n764), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n246), .A2(new_n402), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT50), .Z(new_n1047));
  INV_X1    g0847(.A(new_n712), .ZN(new_n1048));
  AOI211_X1 g0848(.A(G45), .B(new_n1048), .C1(G68), .C2(G77), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n767), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1044), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n760), .B1(new_n1051), .B2(new_n778), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n788), .A2(new_n259), .B1(new_n797), .B2(new_n399), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n417), .B(new_n1053), .C1(G50), .C2(new_n791), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n795), .A2(G77), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n590), .A2(new_n782), .B1(new_n803), .B2(new_n246), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n785), .A2(G159), .B1(new_n805), .B2(G97), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n268), .B1(new_n815), .B2(G326), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n781), .A2(new_n853), .B1(new_n794), .B2(new_n812), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n791), .A2(G317), .B1(new_n817), .B2(G303), .ZN(new_n1061));
  INV_X1    g0861(.A(G311), .ZN(new_n1062));
  INV_X1    g0862(.A(G322), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1061), .B1(new_n852), .B2(new_n1062), .C1(new_n1063), .C2(new_n850), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT48), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1060), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n1065), .B2(new_n1064), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT49), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1059), .B1(new_n622), .B2(new_n804), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1058), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1052), .B1(new_n1071), .B2(new_n773), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n703), .B2(new_n825), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1017), .A2(new_n754), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n710), .B(KEYINPUT115), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1017), .A2(new_n754), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1043), .B(new_n1073), .C1(new_n1076), .C2(new_n1077), .ZN(G393));
  INV_X1    g0878(.A(new_n1014), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n1074), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1080), .A2(new_n1018), .A3(new_n1075), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(KEYINPUT116), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT116), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1080), .A2(new_n1083), .A3(new_n1018), .A4(new_n1075), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n244), .A2(new_n766), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n777), .B1(new_n202), .B2(new_n215), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n850), .A2(new_n399), .B1(new_n798), .B2(new_n790), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT51), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n817), .A2(new_n246), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n855), .B1(G50), .B2(new_n803), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n417), .B1(new_n815), .B2(G143), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n781), .A2(new_n380), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G68), .B2(new_n795), .ZN(new_n1094));
  AND4_X1   g0894(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .A4(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n850), .A2(new_n808), .B1(new_n1062), .B2(new_n790), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT52), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n852), .A2(new_n617), .B1(new_n622), .B2(new_n781), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n417), .B1(new_n797), .B2(new_n1063), .C1(new_n812), .C2(new_n788), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n203), .A2(new_n804), .B1(new_n794), .B2(new_n853), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1089), .A2(new_n1095), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n760), .B1(new_n1086), .B2(new_n1087), .C1(new_n1102), .C2(new_n822), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n1005), .B2(new_n776), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n1014), .B2(new_n759), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1085), .A2(new_n1105), .ZN(G390));
  AND2_X1   g0906(.A1(new_n839), .A2(new_n835), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n895), .A2(new_n896), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n948), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n939), .A2(new_n940), .A3(new_n946), .A4(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n691), .B1(new_n744), .B2(new_n664), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(KEYINPUT96), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1113), .A2(new_n745), .A3(new_n835), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n833), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n948), .B(new_n918), .C1(new_n1115), .C2(new_n1109), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1108), .A2(G330), .A3(new_n731), .A4(new_n838), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1111), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1108), .A2(G330), .A3(new_n838), .A4(new_n902), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n1111), .B2(new_n1116), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n902), .A2(G330), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n487), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n952), .A2(new_n681), .A3(new_n1122), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1114), .A2(new_n833), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n902), .A2(G330), .A3(new_n838), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n1109), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n1117), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n731), .A2(G330), .A3(new_n838), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1121), .A2(new_n897), .B1(new_n1109), .B2(new_n1128), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n1124), .A2(new_n1127), .B1(new_n1129), .B2(new_n1107), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1123), .A2(new_n1130), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n1118), .A2(new_n1120), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1075), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1109), .A2(new_n1128), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1107), .B1(new_n1136), .B2(new_n1119), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n1126), .A2(new_n1117), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1137), .B1(new_n1138), .B2(new_n1115), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n952), .A2(new_n681), .A3(new_n1122), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1134), .B1(new_n1135), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1135), .A2(new_n759), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n852), .A2(new_n203), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1093), .B(new_n1144), .C1(G283), .C2(new_n785), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n790), .A2(new_n622), .B1(new_n797), .B2(new_n812), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n268), .B(new_n1146), .C1(G97), .C2(new_n817), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1145), .A2(new_n796), .A3(new_n861), .A4(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT54), .B(G143), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n790), .A2(new_n865), .B1(new_n788), .B2(new_n1149), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n417), .B(new_n1150), .C1(G125), .C2(new_n815), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n794), .A2(new_n399), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT53), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n803), .A2(G137), .B1(new_n805), .B2(G50), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(G159), .A2(new_n782), .B1(new_n785), .B2(G128), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1151), .A2(new_n1153), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n822), .B1(new_n1148), .B2(new_n1156), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n827), .B(new_n1157), .C1(new_n247), .C2(new_n846), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n947), .B2(new_n775), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1142), .A2(new_n1143), .A3(new_n1159), .ZN(G378));
  INV_X1    g0960(.A(KEYINPUT120), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1111), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1162), .B(new_n1141), .C1(new_n1163), .C2(new_n1119), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n904), .A2(new_n919), .A3(G330), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n413), .A2(new_n877), .ZN(new_n1166));
  XOR2_X1   g0966(.A(new_n438), .B(new_n1166), .Z(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1167), .B(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1165), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1169), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1171), .A2(new_n904), .A3(new_n919), .A4(G330), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n951), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1170), .A2(new_n934), .A3(new_n950), .A4(new_n1172), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n1164), .A2(new_n1123), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1161), .B1(new_n1176), .B2(KEYINPUT57), .ZN(new_n1177));
  AND4_X1   g0977(.A1(new_n950), .A2(new_n1170), .A3(new_n934), .A4(new_n1172), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1172), .A2(new_n1170), .B1(new_n934), .B2(new_n950), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n1132), .A2(new_n1140), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT57), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(KEYINPUT120), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1181), .B1(new_n1164), .B2(new_n1123), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT119), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1179), .A2(KEYINPUT119), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1183), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1177), .A2(new_n1182), .A3(new_n1075), .A4(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n758), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1169), .A2(new_n774), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n268), .A2(G41), .ZN(new_n1191));
  AOI211_X1 g0991(.A(G50), .B(new_n1191), .C1(new_n263), .C2(new_n489), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n790), .A2(new_n203), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1193), .A2(KEYINPUT118), .B1(new_n803), .B2(G97), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1194), .B1(KEYINPUT118), .B2(new_n1193), .C1(new_n622), .C2(new_n850), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n973), .B(new_n1195), .C1(new_n590), .C2(new_n817), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n805), .A2(G58), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n815), .A2(G283), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1055), .A2(new_n1197), .A3(new_n1191), .A4(new_n1198), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT117), .Z(new_n1200));
  AND2_X1   g1000(.A1(new_n1196), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1192), .B1(new_n1201), .B2(KEYINPUT58), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n785), .A2(G125), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n852), .B2(new_n865), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n791), .A2(G128), .B1(new_n817), .B2(G137), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n794), .B2(new_n1149), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(G150), .C2(new_n782), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n805), .A2(G159), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G33), .B(G41), .C1(new_n815), .C2(G124), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1202), .B1(KEYINPUT58), .B2(new_n1201), .C1(new_n1209), .C2(new_n1213), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n1214), .A2(new_n773), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n827), .B(new_n1215), .C1(new_n402), .C2(new_n846), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1189), .B1(new_n1190), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1188), .A2(new_n1217), .ZN(G375));
  INV_X1    g1018(.A(KEYINPUT121), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1123), .A2(new_n1130), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT121), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1222), .A2(new_n1021), .A3(new_n1131), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n622), .A2(new_n852), .B1(new_n850), .B2(new_n812), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G97), .B2(new_n795), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n790), .A2(new_n853), .B1(new_n788), .B2(new_n203), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n268), .B(new_n1226), .C1(G303), .C2(new_n815), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n782), .A2(new_n590), .B1(new_n805), .B2(G77), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1225), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT123), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n850), .A2(new_n865), .B1(new_n402), .B2(new_n781), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G159), .B2(new_n795), .ZN(new_n1232));
  INV_X1    g1032(.A(G128), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n788), .A2(new_n399), .B1(new_n797), .B2(new_n1233), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n417), .B(new_n1234), .C1(G137), .C2(new_n791), .ZN(new_n1235));
  OR2_X1    g1035(.A1(new_n852), .A2(new_n1149), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1232), .A2(new_n1197), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1230), .A2(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1229), .A2(KEYINPUT123), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n773), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n827), .B1(new_n846), .B2(new_n259), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1240), .B(new_n1241), .C1(new_n1108), .C2(new_n775), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n758), .B(KEYINPUT122), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1243), .B1(new_n1130), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1223), .A2(new_n1246), .ZN(G381));
  OR4_X1    g1047(.A1(G396), .A2(G387), .A3(G384), .A4(G393), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1142), .A2(new_n1143), .A3(new_n1159), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1188), .A2(new_n1249), .A3(new_n1217), .ZN(new_n1250));
  OR4_X1    g1050(.A1(G390), .A2(new_n1248), .A3(G381), .A4(new_n1250), .ZN(G407));
  OAI211_X1 g1051(.A(G407), .B(G213), .C1(G343), .C2(new_n1250), .ZN(G409));
  NAND3_X1  g1052(.A1(new_n1188), .A2(G378), .A3(new_n1217), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1245), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1190), .A2(new_n1216), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1254), .B(new_n1255), .C1(new_n1020), .C2(new_n1180), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1249), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1253), .A2(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n686), .A2(G343), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(G384), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT60), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1075), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1131), .A2(KEYINPUT60), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1264), .B1(new_n1222), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1246), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1261), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1262), .A2(new_n1219), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1139), .A2(KEYINPUT121), .A3(new_n1140), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1265), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1264), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(G384), .A3(new_n1246), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1268), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1258), .A2(new_n1260), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1259), .A2(KEYINPUT124), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1268), .A2(new_n1274), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1259), .A2(G2897), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1268), .A2(new_n1274), .A3(new_n1282), .A4(new_n1280), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1284), .A2(KEYINPUT125), .A3(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT125), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  XOR2_X1   g1090(.A(G393), .B(G396), .Z(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(G387), .A2(new_n1085), .A3(new_n1105), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G387), .B1(new_n1085), .B2(new_n1105), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1292), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(G387), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G390), .A2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1298), .A2(new_n1291), .A3(new_n1293), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT61), .ZN(new_n1300));
  AND3_X1   g1100(.A1(new_n1296), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1259), .B1(new_n1253), .B2(new_n1257), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1302), .A2(KEYINPUT63), .A3(new_n1276), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1279), .A2(new_n1290), .A3(new_n1301), .A4(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1300), .B1(new_n1302), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT62), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1277), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1302), .A2(KEYINPUT62), .A3(new_n1276), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1306), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1296), .A2(new_n1299), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT126), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1296), .A2(new_n1299), .A3(KEYINPUT126), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1304), .B1(new_n1310), .B2(new_n1315), .ZN(G405));
  NAND2_X1  g1116(.A1(G375), .A2(new_n1249), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1275), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT127), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1253), .A2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(G375), .A2(new_n1276), .A3(new_n1249), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1318), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1320), .B1(new_n1318), .B2(new_n1321), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1311), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1318), .A2(new_n1321), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1320), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1311), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1328), .A2(new_n1322), .A3(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1325), .A2(new_n1330), .ZN(G402));
endmodule


