//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n823, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939;
  NOR2_X1   g000(.A1(G127gat), .A2(G134gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT70), .B(G127gat), .ZN(new_n204));
  INV_X1    g003(.A(G134gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G113gat), .B(G120gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n208));
  INV_X1    g007(.A(G120gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(G113gat), .ZN(new_n210));
  INV_X1    g009(.A(G113gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(G120gat), .ZN(new_n212));
  NOR3_X1   g011(.A1(new_n210), .A2(new_n212), .A3(KEYINPUT71), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(KEYINPUT71), .A3(G120gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n215));
  AND2_X1   g014(.A1(G127gat), .A2(G134gat), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n214), .B(new_n215), .C1(new_n202), .C2(new_n216), .ZN(new_n217));
  OAI22_X1  g016(.A1(new_n206), .A2(new_n208), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G169gat), .ZN(new_n220));
  INV_X1    g019(.A(G176gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(KEYINPUT66), .B2(KEYINPUT23), .ZN(new_n224));
  AND2_X1   g023(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n222), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G190gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(G183gat), .ZN(new_n228));
  INV_X1    g027(.A(G183gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(G190gat), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT24), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G183gat), .A2(G190gat), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n232), .A2(KEYINPUT24), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n220), .A2(KEYINPUT23), .ZN(new_n234));
  OR2_X1    g033(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n226), .A2(new_n231), .A3(new_n233), .A4(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n239));
  AND3_X1   g038(.A1(new_n238), .A2(KEYINPUT67), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT67), .B1(new_n238), .B2(new_n239), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT25), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n242), .B1(new_n234), .B2(new_n221), .ZN(new_n243));
  AND4_X1   g042(.A1(new_n226), .A2(new_n243), .A3(new_n231), .A4(new_n233), .ZN(new_n244));
  NOR3_X1   g043(.A1(new_n240), .A2(new_n241), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT26), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n222), .A2(new_n246), .A3(new_n223), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n247), .B(new_n232), .C1(new_n246), .C2(new_n222), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n249), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT27), .B(G183gat), .ZN(new_n252));
  OR2_X1    g051(.A1(new_n252), .A2(KEYINPUT68), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(KEYINPUT68), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n253), .A2(KEYINPUT28), .A3(new_n227), .A4(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT28), .ZN(new_n256));
  INV_X1    g055(.A(new_n252), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n256), .B1(new_n257), .B2(G190gat), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n250), .A2(new_n251), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n219), .B1(new_n245), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G227gat), .ZN(new_n261));
  INV_X1    g060(.A(G233gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n238), .A2(new_n239), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n244), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n238), .A2(KEYINPUT67), .A3(new_n239), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n250), .A2(new_n251), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n255), .A2(new_n258), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n268), .A2(new_n218), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n260), .A2(new_n263), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT32), .ZN(new_n274));
  XNOR2_X1  g073(.A(G15gat), .B(G43gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(G71gat), .B(G99gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(KEYINPUT72), .B(KEYINPUT33), .Z(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n277), .B1(new_n273), .B2(KEYINPUT32), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n273), .A2(new_n278), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n283), .B1(new_n282), .B2(new_n284), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n281), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(KEYINPUT74), .B(KEYINPUT34), .Z(new_n288));
  NOR3_X1   g087(.A1(new_n245), .A2(new_n219), .A3(new_n259), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n218), .B1(new_n268), .B2(new_n271), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n288), .B1(new_n291), .B2(new_n263), .ZN(new_n292));
  INV_X1    g091(.A(new_n288), .ZN(new_n293));
  OAI221_X1 g092(.A(new_n293), .B1(new_n261), .B2(new_n262), .C1(new_n289), .C2(new_n290), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n287), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n277), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n274), .A2(new_n284), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT73), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n295), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n281), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n296), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305));
  XNOR2_X1  g104(.A(G197gat), .B(G204gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(G211gat), .A2(G218gat), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(KEYINPUT76), .B2(KEYINPUT22), .ZN(new_n308));
  AND2_X1   g107(.A1(KEYINPUT76), .A2(KEYINPUT22), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n306), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n305), .B1(new_n312), .B2(KEYINPUT29), .ZN(new_n313));
  INV_X1    g112(.A(G141gat), .ZN(new_n314));
  INV_X1    g113(.A(G148gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT2), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT78), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT78), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT2), .ZN(new_n320));
  NAND2_X1  g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n316), .A2(new_n318), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  AND2_X1   g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G155gat), .B(G162gat), .ZN(new_n327));
  INV_X1    g126(.A(G155gat), .ZN(new_n328));
  INV_X1    g127(.A(G162gat), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT2), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n327), .A2(new_n316), .A3(new_n330), .A4(new_n321), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n313), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n326), .A2(new_n305), .A3(new_n331), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n312), .B1(new_n335), .B2(KEYINPUT29), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G228gat), .A2(G233gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n333), .A2(G228gat), .A3(G233gat), .A4(new_n336), .ZN(new_n340));
  NAND2_X1  g139(.A1(KEYINPUT85), .A2(G22gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G78gat), .B(G106gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT31), .B(G50gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n341), .B1(new_n339), .B2(new_n340), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT86), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n347), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT86), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n349), .A2(new_n350), .A3(new_n345), .A4(new_n342), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n339), .A2(new_n340), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT84), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n354), .A2(G22gat), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n354), .A2(G22gat), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n353), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI211_X1 g156(.A(new_n354), .B(G22gat), .C1(new_n339), .C2(new_n340), .ZN(new_n358));
  OR2_X1    g157(.A1(new_n358), .A2(new_n345), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n352), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n304), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G226gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n362), .A2(new_n262), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(KEYINPUT29), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n364), .B1(new_n268), .B2(new_n271), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n312), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n268), .B(new_n271), .C1(new_n362), .C2(new_n262), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NOR3_X1   g168(.A1(new_n245), .A2(new_n259), .A3(new_n363), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n312), .B1(new_n370), .B2(new_n365), .ZN(new_n371));
  XOR2_X1   g170(.A(G8gat), .B(G36gat), .Z(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(KEYINPUT77), .ZN(new_n373));
  XNOR2_X1  g172(.A(G64gat), .B(G92gat), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n373), .B(new_n374), .Z(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n369), .A2(new_n371), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT30), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n369), .A2(new_n371), .A3(KEYINPUT30), .A4(new_n376), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n369), .A2(new_n371), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n375), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT83), .ZN(new_n385));
  XNOR2_X1  g184(.A(G1gat), .B(G29gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT0), .ZN(new_n387));
  XNOR2_X1  g186(.A(G57gat), .B(G85gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n387), .B(new_n388), .Z(new_n389));
  AND2_X1   g188(.A1(new_n218), .A2(new_n334), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT79), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n391), .B1(new_n332), .B2(KEYINPUT3), .ZN(new_n392));
  AOI211_X1 g191(.A(KEYINPUT79), .B(new_n305), .C1(new_n326), .C2(new_n331), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n390), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT4), .B1(new_n218), .B2(new_n332), .ZN(new_n395));
  XNOR2_X1  g194(.A(G141gat), .B(G148gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n325), .A2(new_n396), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n397), .A2(new_n330), .B1(new_n325), .B2(new_n322), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT71), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n207), .A2(new_n400), .ZN(new_n401));
  OR2_X1    g200(.A1(new_n216), .A2(new_n202), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n401), .A2(new_n215), .A3(new_n402), .A4(new_n214), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n215), .B1(new_n210), .B2(new_n212), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n404), .B(new_n203), .C1(new_n205), .C2(new_n204), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n398), .A2(new_n399), .A3(new_n403), .A4(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n395), .A2(new_n406), .A3(KEYINPUT80), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n408), .B(KEYINPUT4), .C1(new_n218), .C2(new_n332), .ZN(new_n409));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n394), .A2(new_n407), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT5), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n218), .B(new_n332), .ZN(new_n413));
  INV_X1    g212(.A(new_n410), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT79), .B1(new_n398), .B2(new_n305), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n332), .A2(new_n391), .A3(KEYINPUT3), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n414), .B1(new_n419), .B2(new_n390), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT5), .B1(new_n395), .B2(new_n406), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n389), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n385), .B1(new_n423), .B2(KEYINPUT6), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n411), .A2(new_n415), .B1(new_n420), .B2(new_n421), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n426));
  NOR4_X1   g225(.A1(new_n425), .A2(KEYINPUT83), .A3(new_n426), .A4(new_n389), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n416), .A2(new_n389), .A3(new_n422), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n426), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT81), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n431), .B1(new_n425), .B2(new_n389), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n422), .ZN(new_n433));
  INV_X1    g232(.A(new_n389), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(KEYINPUT81), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n430), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n428), .B1(new_n436), .B2(KEYINPUT82), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n432), .ZN(new_n438));
  INV_X1    g237(.A(new_n430), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(KEYINPUT82), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n384), .B1(new_n437), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT35), .B1(new_n361), .B2(new_n442), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n357), .A2(new_n358), .A3(new_n345), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n444), .B1(new_n348), .B2(new_n351), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n445), .B1(new_n296), .B2(new_n303), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n383), .A2(KEYINPUT88), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT88), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n379), .A2(new_n382), .A3(new_n448), .A4(new_n380), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n434), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n439), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT35), .B1(new_n428), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n446), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n443), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g254(.A(KEYINPUT89), .B(new_n312), .C1(new_n370), .C2(new_n365), .ZN(new_n456));
  OAI211_X1 g255(.A(KEYINPUT37), .B(new_n456), .C1(new_n381), .C2(KEYINPUT89), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT38), .ZN(new_n458));
  XNOR2_X1  g257(.A(KEYINPUT90), .B(KEYINPUT37), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n369), .A2(new_n371), .A3(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n457), .A2(new_n458), .A3(new_n375), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n375), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT37), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n463), .B1(new_n369), .B2(new_n371), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT38), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n428), .A2(new_n452), .A3(new_n377), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n360), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT40), .ZN(new_n469));
  INV_X1    g268(.A(new_n394), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n395), .A2(new_n406), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n414), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n413), .A2(new_n414), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n472), .A2(KEYINPUT39), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n389), .B1(new_n472), .B2(KEYINPUT39), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n469), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n451), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n474), .A2(new_n475), .A3(new_n469), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n447), .A2(new_n479), .A3(new_n449), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n468), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n302), .B1(new_n301), .B2(new_n281), .ZN(new_n482));
  AOI211_X1 g281(.A(new_n280), .B(new_n295), .C1(new_n299), .C2(new_n300), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT36), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  XOR2_X1   g283(.A(KEYINPUT75), .B(KEYINPUT36), .Z(new_n485));
  NAND3_X1  g284(.A1(new_n296), .A2(new_n303), .A3(new_n485), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n484), .A2(new_n486), .B1(new_n442), .B2(new_n445), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n481), .B1(new_n487), .B2(KEYINPUT87), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n442), .A2(new_n445), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n296), .A2(new_n303), .A3(new_n485), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT36), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n296), .B2(new_n303), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n489), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT87), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n455), .B1(new_n488), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT97), .ZN(new_n497));
  AOI21_X1  g296(.A(G64gat), .B1(new_n497), .B2(G57gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(KEYINPUT96), .A3(G57gat), .ZN(new_n499));
  OR2_X1    g298(.A1(KEYINPUT96), .A2(G57gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n498), .B1(new_n501), .B2(G64gat), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n502), .A2(KEYINPUT98), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(KEYINPUT98), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G71gat), .ZN(new_n506));
  INV_X1    g305(.A(G78gat), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(G71gat), .A2(G78gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT9), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n514), .B1(G57gat), .B2(G64gat), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n515), .A2(new_n508), .A3(new_n510), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT21), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(G127gat), .B(G155gat), .Z(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT93), .ZN(new_n524));
  INV_X1    g323(.A(G1gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n523), .A2(KEYINPUT93), .A3(G1gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT16), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n523), .A2(new_n528), .B1(KEYINPUT94), .B2(G8gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(new_n518), .B2(new_n519), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n522), .B(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(G231gat), .A2(G233gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT99), .ZN(new_n536));
  XOR2_X1   g335(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G183gat), .B(G211gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n534), .B(new_n540), .Z(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G50gat), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT15), .B1(new_n543), .B2(G43gat), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n544), .B1(G43gat), .B2(new_n543), .ZN(new_n545));
  XOR2_X1   g344(.A(KEYINPUT14), .B(G29gat), .Z(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(G36gat), .ZN(new_n547));
  INV_X1    g346(.A(G29gat), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n548), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n545), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n547), .A2(new_n549), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT91), .B(G43gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(G50gat), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT92), .B1(new_n543), .B2(G43gat), .ZN(new_n554));
  OR2_X1    g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT92), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT15), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n551), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n550), .B1(new_n558), .B2(new_n545), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n559), .A2(KEYINPUT17), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(KEYINPUT17), .ZN(new_n561));
  NAND2_X1  g360(.A1(G85gat), .A2(G92gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n562), .B(new_n563), .Z(new_n564));
  NAND2_X1  g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565));
  INV_X1    g364(.A(G85gat), .ZN(new_n566));
  INV_X1    g365(.A(G92gat), .ZN(new_n567));
  AOI22_X1  g366(.A1(KEYINPUT8), .A2(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G99gat), .B(G106gat), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n569), .B(new_n570), .Z(new_n571));
  NAND3_X1  g370(.A1(new_n560), .A2(new_n561), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n559), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n569), .B(new_n570), .ZN(new_n574));
  AND2_X1   g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575));
  AOI22_X1  g374(.A1(new_n573), .A2(new_n574), .B1(KEYINPUT41), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(G190gat), .B(G218gat), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n575), .A2(KEYINPUT41), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT100), .ZN(new_n581));
  XNOR2_X1  g380(.A(G134gat), .B(G162gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n579), .A2(new_n584), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G230gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(new_n262), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n503), .A2(new_n504), .B1(new_n509), .B2(new_n511), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n571), .B1(new_n591), .B2(new_n516), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n513), .A2(new_n517), .A3(new_n574), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT10), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n513), .A2(new_n574), .A3(KEYINPUT10), .A4(new_n517), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n590), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n592), .A2(new_n593), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n590), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G120gat), .B(G148gat), .Z(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT102), .ZN(new_n603));
  XNOR2_X1  g402(.A(G176gat), .B(G204gat), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n603), .B(new_n604), .Z(new_n605));
  NAND2_X1  g404(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n605), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n598), .A2(new_n600), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n542), .A2(new_n588), .A3(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n559), .A2(new_n532), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT95), .ZN(new_n613));
  INV_X1    g412(.A(new_n532), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n613), .B1(new_n573), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G229gat), .A2(G233gat), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n616), .B(KEYINPUT13), .Z(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n560), .A2(new_n532), .A3(new_n561), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n613), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT18), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n613), .A2(KEYINPUT18), .A3(new_n616), .A4(new_n619), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n618), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G113gat), .B(G141gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(G197gat), .ZN(new_n626));
  XOR2_X1   g425(.A(KEYINPUT11), .B(G169gat), .Z(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n628), .B(KEYINPUT12), .Z(new_n629));
  NAND2_X1  g428(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n629), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n618), .A2(new_n622), .A3(new_n631), .A4(new_n623), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n611), .A2(new_n634), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n496), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n437), .A2(new_n441), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(G1gat), .ZN(G1324gat));
  INV_X1    g438(.A(KEYINPUT42), .ZN(new_n640));
  INV_X1    g439(.A(new_n450), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n636), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT103), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT16), .B(G8gat), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n640), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(G8gat), .ZN(new_n646));
  OR3_X1    g445(.A1(new_n642), .A2(new_n640), .A3(new_n644), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(G1325gat));
  INV_X1    g447(.A(new_n636), .ZN(new_n649));
  INV_X1    g448(.A(new_n304), .ZN(new_n650));
  OR3_X1    g449(.A1(new_n649), .A2(G15gat), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n490), .A2(new_n492), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(G15gat), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(G1326gat));
  NAND2_X1  g454(.A1(new_n636), .A2(new_n445), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT43), .B(G22gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(G1327gat));
  NAND2_X1  g457(.A1(new_n496), .A2(new_n587), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n542), .A2(new_n634), .A3(new_n609), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n663), .A2(new_n548), .A3(new_n637), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT35), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT82), .B1(new_n438), .B2(new_n439), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT83), .B1(new_n451), .B2(new_n426), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n423), .A2(new_n385), .A3(KEYINPUT6), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n383), .B1(new_n672), .B2(new_n440), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n667), .B1(new_n446), .B2(new_n673), .ZN(new_n674));
  AND4_X1   g473(.A1(new_n304), .A2(new_n453), .A3(new_n360), .A4(new_n450), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n468), .A2(new_n480), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n677), .B1(new_n493), .B2(new_n494), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n487), .A2(KEYINPUT87), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n676), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI211_X1 g479(.A(KEYINPUT105), .B(KEYINPUT44), .C1(new_n680), .C2(new_n588), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  OAI22_X1  g481(.A1(new_n455), .A2(KEYINPUT106), .B1(new_n493), .B2(new_n677), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n676), .A2(new_n684), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n682), .B(new_n587), .C1(new_n683), .C2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT105), .B1(new_n659), .B2(KEYINPUT44), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n661), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT107), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n691), .B(new_n661), .C1(new_n687), .C2(new_n688), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n690), .A2(new_n637), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n666), .B1(new_n693), .B2(new_n548), .ZN(G1328gat));
  NOR3_X1   g493(.A1(new_n662), .A2(G36gat), .A3(new_n450), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT46), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n690), .A2(new_n641), .A3(new_n692), .ZN(new_n697));
  INV_X1    g496(.A(G36gat), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(G1329gat));
  INV_X1    g498(.A(new_n552), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n700), .B1(new_n689), .B2(new_n653), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n650), .A2(new_n700), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n663), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n701), .A2(KEYINPUT47), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n690), .A2(new_n652), .A3(new_n692), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n705), .A2(new_n700), .B1(new_n663), .B2(new_n702), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n706), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g506(.A(G50gat), .B1(new_n689), .B2(new_n360), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n663), .A2(new_n543), .A3(new_n445), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(KEYINPUT48), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n690), .A2(new_n445), .A3(new_n692), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n712), .A3(G50gat), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT48), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n709), .A2(KEYINPUT108), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n711), .B2(G50gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n710), .B1(new_n715), .B2(new_n717), .ZN(G1331gat));
  OR2_X1    g517(.A1(new_n683), .A2(new_n685), .ZN(new_n719));
  NOR4_X1   g518(.A1(new_n633), .A2(new_n541), .A3(new_n587), .A4(new_n610), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n637), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT109), .ZN(new_n724));
  XOR2_X1   g523(.A(KEYINPUT96), .B(G57gat), .Z(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1332gat));
  INV_X1    g525(.A(KEYINPUT49), .ZN(new_n727));
  INV_X1    g526(.A(G64gat), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n722), .B(new_n641), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT110), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n727), .A2(new_n728), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1333gat));
  NAND3_X1  g531(.A1(new_n722), .A2(G71gat), .A3(new_n652), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT111), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n506), .B1(new_n721), .B2(new_n650), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT50), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT50), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n734), .A2(new_n738), .A3(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1334gat));
  NOR2_X1   g539(.A1(new_n721), .A2(new_n360), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(new_n507), .ZN(G1335gat));
  NOR2_X1   g541(.A1(new_n542), .A2(new_n633), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n587), .B(new_n743), .C1(new_n683), .C2(new_n685), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT51), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n746), .A2(new_n566), .A3(new_n637), .A4(new_n609), .ZN(new_n747));
  OR2_X1    g546(.A1(new_n687), .A2(new_n688), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n542), .A2(new_n633), .A3(new_n610), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n748), .A2(new_n637), .A3(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n747), .B1(new_n751), .B2(new_n566), .ZN(G1336gat));
  NAND3_X1  g551(.A1(new_n748), .A2(new_n641), .A3(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G92gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n744), .A2(KEYINPUT112), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n744), .A2(KEYINPUT112), .A3(KEYINPUT51), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n450), .A2(G92gat), .A3(new_n610), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n760), .A2(KEYINPUT113), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(KEYINPUT113), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n754), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT52), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT52), .B1(new_n746), .B2(new_n759), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n754), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(G1337gat));
  XOR2_X1   g566(.A(KEYINPUT114), .B(G99gat), .Z(new_n768));
  NAND4_X1  g567(.A1(new_n746), .A2(new_n304), .A3(new_n609), .A4(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n748), .A2(new_n652), .A3(new_n749), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n771), .B2(new_n768), .ZN(G1338gat));
  NAND3_X1  g571(.A1(new_n748), .A2(new_n445), .A3(new_n749), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G106gat), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n360), .A2(new_n610), .A3(G106gat), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT53), .B1(new_n746), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n757), .A2(new_n758), .A3(new_n775), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n777), .B1(new_n779), .B2(new_n780), .ZN(G1339gat));
  NOR2_X1   g580(.A1(new_n615), .A2(new_n617), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n616), .B1(new_n613), .B2(new_n619), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n628), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n784), .A2(new_n632), .A3(new_n609), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT117), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n595), .A2(new_n596), .A3(new_n590), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n598), .A2(KEYINPUT54), .A3(new_n788), .ZN(new_n789));
  AOI211_X1 g588(.A(KEYINPUT54), .B(new_n590), .C1(new_n595), .C2(new_n596), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n790), .A2(new_n791), .A3(new_n607), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n597), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT115), .B1(new_n794), .B2(new_n605), .ZN(new_n795));
  OAI211_X1 g594(.A(KEYINPUT55), .B(new_n789), .C1(new_n792), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n608), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n791), .B1(new_n790), .B2(new_n607), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n794), .A2(KEYINPUT115), .A3(new_n605), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT55), .B1(new_n800), .B2(new_n789), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n633), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n587), .B1(new_n787), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n784), .A2(new_n632), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n587), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n805), .B1(new_n784), .B2(new_n632), .ZN(new_n808));
  NOR4_X1   g607(.A1(new_n807), .A2(new_n801), .A3(new_n808), .A4(new_n797), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n541), .B1(new_n804), .B2(new_n809), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n611), .A2(new_n633), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n812), .A2(new_n637), .A3(new_n446), .A4(new_n450), .ZN(new_n813));
  OAI21_X1  g612(.A(G113gat), .B1(new_n813), .B2(new_n634), .ZN(new_n814));
  XOR2_X1   g613(.A(new_n814), .B(KEYINPUT118), .Z(new_n815));
  AND2_X1   g614(.A1(new_n812), .A2(new_n637), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n816), .A2(new_n446), .A3(new_n450), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(new_n211), .A3(new_n633), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n818), .ZN(G1340gat));
  NOR3_X1   g618(.A1(new_n813), .A2(new_n209), .A3(new_n610), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n817), .A2(new_n609), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n820), .B1(new_n821), .B2(new_n209), .ZN(G1341gat));
  NAND3_X1  g621(.A1(new_n817), .A2(new_n204), .A3(new_n542), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n813), .A2(new_n541), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n823), .B1(new_n204), .B2(new_n824), .ZN(G1342gat));
  NOR3_X1   g624(.A1(new_n588), .A2(new_n641), .A3(G134gat), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n816), .A2(new_n446), .A3(new_n826), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n827), .A2(KEYINPUT56), .ZN(new_n828));
  OAI21_X1  g627(.A(G134gat), .B1(new_n813), .B2(new_n588), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(KEYINPUT56), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(G1343gat));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n637), .A2(new_n450), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n652), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n360), .B1(new_n810), .B2(new_n811), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT119), .B1(new_n797), .B2(new_n801), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n800), .A2(new_n789), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n842), .A2(new_n843), .A3(new_n608), .A4(new_n796), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n839), .A2(new_n844), .A3(new_n633), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n785), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n809), .B1(new_n846), .B2(new_n588), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n811), .B1(new_n847), .B2(new_n542), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(new_n445), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n838), .B(new_n633), .C1(new_n849), .C2(new_n837), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(G141gat), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n652), .A2(new_n360), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n816), .A2(new_n852), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n853), .A2(KEYINPUT121), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(KEYINPUT121), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(new_n450), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n633), .A2(new_n314), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n832), .B(new_n851), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n853), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n857), .A2(new_n641), .ZN(new_n860));
  AOI22_X1  g659(.A1(new_n850), .A2(G141gat), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n832), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(KEYINPUT120), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n861), .A2(new_n864), .A3(new_n832), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n858), .B1(new_n863), .B2(new_n865), .ZN(G1344gat));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n848), .A2(new_n868), .ZN(new_n869));
  OAI211_X1 g668(.A(KEYINPUT122), .B(new_n811), .C1(new_n847), .C2(new_n542), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n360), .A2(KEYINPUT57), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n836), .A2(new_n837), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n609), .A3(new_n834), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n867), .B1(new_n875), .B2(G148gat), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n838), .B1(new_n849), .B2(new_n837), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n610), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n878), .A2(KEYINPUT59), .A3(new_n315), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n609), .A2(new_n315), .ZN(new_n880));
  OAI22_X1  g679(.A1(new_n876), .A2(new_n879), .B1(new_n856), .B2(new_n880), .ZN(G1345gat));
  OAI21_X1  g680(.A(G155gat), .B1(new_n877), .B2(new_n541), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n542), .A2(new_n328), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n856), .B2(new_n883), .ZN(G1346gat));
  OAI21_X1  g683(.A(G162gat), .B1(new_n877), .B2(new_n588), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n587), .A2(new_n329), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n856), .B2(new_n886), .ZN(G1347gat));
  NOR2_X1   g686(.A1(new_n637), .A2(new_n450), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n889), .B1(new_n810), .B2(new_n811), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n446), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n634), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(new_n220), .ZN(G1348gat));
  INV_X1    g692(.A(new_n891), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n609), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(G176gat), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n235), .A2(new_n236), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(new_n895), .ZN(G1349gat));
  NAND4_X1  g697(.A1(new_n894), .A2(new_n253), .A3(new_n254), .A4(new_n542), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900));
  OAI21_X1  g699(.A(G183gat), .B1(new_n891), .B2(new_n541), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g702(.A1(new_n894), .A2(new_n587), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n904), .A2(G190gat), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(G190gat), .ZN(new_n906));
  XNOR2_X1  g705(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n908), .B1(new_n906), .B2(new_n907), .ZN(G1351gat));
  AND2_X1   g708(.A1(new_n890), .A2(new_n852), .ZN(new_n910));
  AOI21_X1  g709(.A(G197gat), .B1(new_n910), .B2(new_n633), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n652), .A2(new_n889), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n874), .A2(new_n912), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n633), .A2(G197gat), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(G1352gat));
  NAND3_X1  g714(.A1(new_n874), .A2(new_n609), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(G204gat), .ZN(new_n917));
  INV_X1    g716(.A(G204gat), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n910), .A2(new_n918), .A3(new_n609), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n919), .B(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT125), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n917), .A2(KEYINPUT125), .A3(new_n921), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1353gat));
  INV_X1    g725(.A(G211gat), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n910), .A2(new_n927), .A3(new_n542), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n872), .A2(new_n873), .A3(new_n542), .A4(new_n912), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n929), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT63), .B1(new_n929), .B2(G211gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT126), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n934), .B(new_n928), .C1(new_n930), .C2(new_n931), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1354gat));
  AOI21_X1  g735(.A(G218gat), .B1(new_n910), .B2(new_n587), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n587), .A2(G218gat), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT127), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n937), .B1(new_n913), .B2(new_n939), .ZN(G1355gat));
endmodule


