

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U552 ( .A(n773), .ZN(n753) );
  AND2_X1 U553 ( .A1(n779), .A2(n777), .ZN(n769) );
  AND2_X1 U554 ( .A1(n753), .A2(G1996), .ZN(n723) );
  AND2_X1 U555 ( .A1(G2104), .A2(n522), .ZN(n519) );
  XNOR2_X1 U556 ( .A(n518), .B(KEYINPUT102), .ZN(n809) );
  NAND2_X1 U557 ( .A1(n799), .A2(n790), .ZN(n518) );
  AND2_X1 U558 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U559 ( .A1(n770), .A2(n769), .ZN(n771) );
  AND2_X1 U560 ( .A1(n725), .A2(n724), .ZN(n732) );
  INV_X1 U561 ( .A(KEYINPUT96), .ZN(n737) );
  INV_X1 U562 ( .A(KEYINPUT101), .ZN(n806) );
  XNOR2_X1 U563 ( .A(n807), .B(n806), .ZN(n808) );
  NOR2_X1 U564 ( .A1(G164), .A2(G1384), .ZN(n718) );
  NOR2_X1 U565 ( .A1(G651), .A2(n639), .ZN(n657) );
  INV_X1 U566 ( .A(G2105), .ZN(n522) );
  XNOR2_X2 U567 ( .A(n519), .B(KEYINPUT64), .ZN(n883) );
  AND2_X1 U568 ( .A1(n883), .A2(G102), .ZN(n520) );
  XNOR2_X1 U569 ( .A(n520), .B(KEYINPUT82), .ZN(n526) );
  AND2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n886) );
  NAND2_X1 U571 ( .A1(G114), .A2(n886), .ZN(n521) );
  XNOR2_X1 U572 ( .A(KEYINPUT81), .B(n521), .ZN(n524) );
  NOR2_X1 U573 ( .A1(G2104), .A2(n522), .ZN(n887) );
  AND2_X1 U574 ( .A1(n887), .A2(G126), .ZN(n523) );
  OR2_X1 U575 ( .A1(n524), .A2(n523), .ZN(n525) );
  OR2_X1 U576 ( .A1(n526), .A2(n525), .ZN(n530) );
  NOR2_X1 U577 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  XOR2_X2 U578 ( .A(KEYINPUT17), .B(n527), .Z(n882) );
  NAND2_X1 U579 ( .A1(G138), .A2(n882), .ZN(n528) );
  XNOR2_X1 U580 ( .A(KEYINPUT83), .B(n528), .ZN(n529) );
  NOR2_X2 U581 ( .A1(n530), .A2(n529), .ZN(G164) );
  NAND2_X1 U582 ( .A1(G113), .A2(n886), .ZN(n532) );
  NAND2_X1 U583 ( .A1(G125), .A2(n887), .ZN(n531) );
  NAND2_X1 U584 ( .A1(n532), .A2(n531), .ZN(n537) );
  NAND2_X1 U585 ( .A1(n883), .A2(G101), .ZN(n533) );
  XOR2_X1 U586 ( .A(KEYINPUT23), .B(n533), .Z(n535) );
  NAND2_X1 U587 ( .A1(n882), .A2(G137), .ZN(n534) );
  NAND2_X1 U588 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U589 ( .A1(n537), .A2(n536), .ZN(G160) );
  NOR2_X1 U590 ( .A1(G651), .A2(G543), .ZN(n649) );
  NAND2_X1 U591 ( .A1(G85), .A2(n649), .ZN(n539) );
  XOR2_X1 U592 ( .A(KEYINPUT0), .B(G543), .Z(n639) );
  INV_X1 U593 ( .A(G651), .ZN(n540) );
  NOR2_X1 U594 ( .A1(n639), .A2(n540), .ZN(n653) );
  NAND2_X1 U595 ( .A1(G72), .A2(n653), .ZN(n538) );
  NAND2_X1 U596 ( .A1(n539), .A2(n538), .ZN(n545) );
  NOR2_X1 U597 ( .A1(G543), .A2(n540), .ZN(n541) );
  XOR2_X1 U598 ( .A(KEYINPUT1), .B(n541), .Z(n650) );
  NAND2_X1 U599 ( .A1(G60), .A2(n650), .ZN(n543) );
  NAND2_X1 U600 ( .A1(G47), .A2(n657), .ZN(n542) );
  NAND2_X1 U601 ( .A1(n543), .A2(n542), .ZN(n544) );
  OR2_X1 U602 ( .A1(n545), .A2(n544), .ZN(G290) );
  XNOR2_X1 U603 ( .A(G2451), .B(G2443), .ZN(n555) );
  XOR2_X1 U604 ( .A(G2446), .B(KEYINPUT105), .Z(n547) );
  XNOR2_X1 U605 ( .A(G2438), .B(G2435), .ZN(n546) );
  XNOR2_X1 U606 ( .A(n547), .B(n546), .ZN(n551) );
  XOR2_X1 U607 ( .A(KEYINPUT106), .B(G2454), .Z(n549) );
  XNOR2_X1 U608 ( .A(G1341), .B(G1348), .ZN(n548) );
  XNOR2_X1 U609 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U610 ( .A(n551), .B(n550), .Z(n553) );
  XNOR2_X1 U611 ( .A(G2430), .B(G2427), .ZN(n552) );
  XNOR2_X1 U612 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U613 ( .A(n555), .B(n554), .ZN(n556) );
  AND2_X1 U614 ( .A1(n556), .A2(G14), .ZN(G401) );
  NAND2_X1 U615 ( .A1(G64), .A2(n650), .ZN(n558) );
  NAND2_X1 U616 ( .A1(G52), .A2(n657), .ZN(n557) );
  NAND2_X1 U617 ( .A1(n558), .A2(n557), .ZN(n565) );
  XNOR2_X1 U618 ( .A(KEYINPUT66), .B(KEYINPUT9), .ZN(n563) );
  NAND2_X1 U619 ( .A1(n653), .A2(G77), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n649), .A2(G90), .ZN(n559) );
  XOR2_X1 U621 ( .A(KEYINPUT65), .B(n559), .Z(n560) );
  NAND2_X1 U622 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U623 ( .A(n563), .B(n562), .Z(n564) );
  NOR2_X1 U624 ( .A1(n565), .A2(n564), .ZN(G171) );
  AND2_X1 U625 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U626 ( .A(G57), .ZN(G237) );
  INV_X1 U627 ( .A(G132), .ZN(G219) );
  INV_X1 U628 ( .A(G82), .ZN(G220) );
  NAND2_X1 U629 ( .A1(G89), .A2(n649), .ZN(n566) );
  XNOR2_X1 U630 ( .A(n566), .B(KEYINPUT72), .ZN(n567) );
  XNOR2_X1 U631 ( .A(KEYINPUT4), .B(n567), .ZN(n570) );
  NAND2_X1 U632 ( .A1(n653), .A2(G76), .ZN(n568) );
  XOR2_X1 U633 ( .A(KEYINPUT73), .B(n568), .Z(n569) );
  NAND2_X1 U634 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U635 ( .A(KEYINPUT5), .B(n571), .ZN(n577) );
  NAND2_X1 U636 ( .A1(G63), .A2(n650), .ZN(n573) );
  NAND2_X1 U637 ( .A1(G51), .A2(n657), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n575) );
  XOR2_X1 U639 ( .A(KEYINPUT74), .B(KEYINPUT6), .Z(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U642 ( .A(KEYINPUT7), .B(n578), .ZN(G168) );
  XOR2_X1 U643 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U644 ( .A1(G7), .A2(G661), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n579), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U646 ( .A(G223), .B(KEYINPUT68), .Z(n833) );
  NAND2_X1 U647 ( .A1(n833), .A2(G567), .ZN(n580) );
  XOR2_X1 U648 ( .A(KEYINPUT11), .B(n580), .Z(G234) );
  XNOR2_X1 U649 ( .A(KEYINPUT13), .B(KEYINPUT69), .ZN(n585) );
  NAND2_X1 U650 ( .A1(n649), .A2(G81), .ZN(n581) );
  XNOR2_X1 U651 ( .A(n581), .B(KEYINPUT12), .ZN(n583) );
  NAND2_X1 U652 ( .A1(G68), .A2(n653), .ZN(n582) );
  NAND2_X1 U653 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U654 ( .A(n585), .B(n584), .ZN(n588) );
  NAND2_X1 U655 ( .A1(n650), .A2(G56), .ZN(n586) );
  XOR2_X1 U656 ( .A(KEYINPUT14), .B(n586), .Z(n587) );
  NOR2_X1 U657 ( .A1(n588), .A2(n587), .ZN(n590) );
  NAND2_X1 U658 ( .A1(n657), .A2(G43), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n930) );
  INV_X1 U660 ( .A(G860), .ZN(n628) );
  OR2_X1 U661 ( .A1(n930), .A2(n628), .ZN(G153) );
  XOR2_X1 U662 ( .A(G171), .B(KEYINPUT70), .Z(G301) );
  NAND2_X1 U663 ( .A1(G868), .A2(G301), .ZN(n591) );
  XOR2_X1 U664 ( .A(KEYINPUT71), .B(n591), .Z(n600) );
  NAND2_X1 U665 ( .A1(G92), .A2(n649), .ZN(n593) );
  NAND2_X1 U666 ( .A1(G79), .A2(n653), .ZN(n592) );
  NAND2_X1 U667 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U668 ( .A1(G66), .A2(n650), .ZN(n595) );
  NAND2_X1 U669 ( .A1(G54), .A2(n657), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U672 ( .A(KEYINPUT15), .B(n598), .Z(n919) );
  INV_X1 U673 ( .A(n919), .ZN(n613) );
  INV_X1 U674 ( .A(G868), .ZN(n612) );
  NAND2_X1 U675 ( .A1(n613), .A2(n612), .ZN(n599) );
  NAND2_X1 U676 ( .A1(n600), .A2(n599), .ZN(G284) );
  NAND2_X1 U677 ( .A1(G91), .A2(n649), .ZN(n602) );
  NAND2_X1 U678 ( .A1(G78), .A2(n653), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n602), .A2(n601), .ZN(n605) );
  NAND2_X1 U680 ( .A1(G65), .A2(n650), .ZN(n603) );
  XNOR2_X1 U681 ( .A(KEYINPUT67), .B(n603), .ZN(n604) );
  NOR2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n657), .A2(G53), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n607), .A2(n606), .ZN(G299) );
  NOR2_X1 U685 ( .A1(G286), .A2(n612), .ZN(n609) );
  NOR2_X1 U686 ( .A1(G868), .A2(G299), .ZN(n608) );
  NOR2_X1 U687 ( .A1(n609), .A2(n608), .ZN(G297) );
  NAND2_X1 U688 ( .A1(n628), .A2(G559), .ZN(n610) );
  NAND2_X1 U689 ( .A1(n610), .A2(n919), .ZN(n611) );
  XNOR2_X1 U690 ( .A(n611), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U691 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U692 ( .A(n614), .B(KEYINPUT75), .ZN(n615) );
  NOR2_X1 U693 ( .A1(G559), .A2(n615), .ZN(n617) );
  NOR2_X1 U694 ( .A1(G868), .A2(n930), .ZN(n616) );
  NOR2_X1 U695 ( .A1(n617), .A2(n616), .ZN(G282) );
  NAND2_X1 U696 ( .A1(G123), .A2(n887), .ZN(n618) );
  XNOR2_X1 U697 ( .A(n618), .B(KEYINPUT18), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n886), .A2(G111), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n882), .A2(G135), .ZN(n622) );
  NAND2_X1 U701 ( .A1(G99), .A2(n883), .ZN(n621) );
  NAND2_X1 U702 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U703 ( .A1(n624), .A2(n623), .ZN(n970) );
  XNOR2_X1 U704 ( .A(n970), .B(G2096), .ZN(n626) );
  INV_X1 U705 ( .A(G2100), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(G156) );
  NAND2_X1 U707 ( .A1(G559), .A2(n919), .ZN(n627) );
  XOR2_X1 U708 ( .A(n930), .B(n627), .Z(n665) );
  NAND2_X1 U709 ( .A1(n628), .A2(n665), .ZN(n635) );
  NAND2_X1 U710 ( .A1(G67), .A2(n650), .ZN(n630) );
  NAND2_X1 U711 ( .A1(G55), .A2(n657), .ZN(n629) );
  NAND2_X1 U712 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U713 ( .A1(G93), .A2(n649), .ZN(n632) );
  NAND2_X1 U714 ( .A1(G80), .A2(n653), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U716 ( .A1(n634), .A2(n633), .ZN(n667) );
  XOR2_X1 U717 ( .A(n635), .B(n667), .Z(G145) );
  NAND2_X1 U718 ( .A1(G49), .A2(n657), .ZN(n637) );
  NAND2_X1 U719 ( .A1(G74), .A2(G651), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U721 ( .A1(n650), .A2(n638), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n639), .A2(G87), .ZN(n640) );
  NAND2_X1 U723 ( .A1(n641), .A2(n640), .ZN(G288) );
  NAND2_X1 U724 ( .A1(G88), .A2(n649), .ZN(n643) );
  NAND2_X1 U725 ( .A1(G62), .A2(n650), .ZN(n642) );
  NAND2_X1 U726 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U727 ( .A1(n653), .A2(G75), .ZN(n644) );
  XOR2_X1 U728 ( .A(KEYINPUT76), .B(n644), .Z(n645) );
  NOR2_X1 U729 ( .A1(n646), .A2(n645), .ZN(n648) );
  NAND2_X1 U730 ( .A1(n657), .A2(G50), .ZN(n647) );
  NAND2_X1 U731 ( .A1(n648), .A2(n647), .ZN(G303) );
  INV_X1 U732 ( .A(G303), .ZN(G166) );
  NAND2_X1 U733 ( .A1(G86), .A2(n649), .ZN(n652) );
  NAND2_X1 U734 ( .A1(G61), .A2(n650), .ZN(n651) );
  NAND2_X1 U735 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U736 ( .A1(n653), .A2(G73), .ZN(n654) );
  XOR2_X1 U737 ( .A(KEYINPUT2), .B(n654), .Z(n655) );
  NOR2_X1 U738 ( .A1(n656), .A2(n655), .ZN(n659) );
  NAND2_X1 U739 ( .A1(n657), .A2(G48), .ZN(n658) );
  NAND2_X1 U740 ( .A1(n659), .A2(n658), .ZN(G305) );
  XNOR2_X1 U741 ( .A(G166), .B(KEYINPUT19), .ZN(n661) );
  INV_X1 U742 ( .A(G299), .ZN(n746) );
  XNOR2_X1 U743 ( .A(G290), .B(n746), .ZN(n660) );
  XNOR2_X1 U744 ( .A(n661), .B(n660), .ZN(n662) );
  XOR2_X1 U745 ( .A(n667), .B(n662), .Z(n663) );
  XNOR2_X1 U746 ( .A(G288), .B(n663), .ZN(n664) );
  XNOR2_X1 U747 ( .A(n664), .B(G305), .ZN(n843) );
  XNOR2_X1 U748 ( .A(n665), .B(n843), .ZN(n666) );
  NAND2_X1 U749 ( .A1(n666), .A2(G868), .ZN(n669) );
  OR2_X1 U750 ( .A1(G868), .A2(n667), .ZN(n668) );
  NAND2_X1 U751 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2078), .A2(G2084), .ZN(n670) );
  XNOR2_X1 U753 ( .A(n670), .B(KEYINPUT77), .ZN(n671) );
  XNOR2_X1 U754 ( .A(n671), .B(KEYINPUT20), .ZN(n672) );
  NAND2_X1 U755 ( .A1(n672), .A2(G2090), .ZN(n673) );
  XNOR2_X1 U756 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U757 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U759 ( .A1(G220), .A2(G219), .ZN(n675) );
  XNOR2_X1 U760 ( .A(KEYINPUT22), .B(n675), .ZN(n676) );
  NAND2_X1 U761 ( .A1(n676), .A2(G96), .ZN(n677) );
  NOR2_X1 U762 ( .A1(G218), .A2(n677), .ZN(n678) );
  XOR2_X1 U763 ( .A(KEYINPUT78), .B(n678), .Z(n840) );
  NAND2_X1 U764 ( .A1(n840), .A2(G2106), .ZN(n682) );
  NAND2_X1 U765 ( .A1(G69), .A2(G120), .ZN(n679) );
  NOR2_X1 U766 ( .A1(G237), .A2(n679), .ZN(n680) );
  NAND2_X1 U767 ( .A1(G108), .A2(n680), .ZN(n839) );
  NAND2_X1 U768 ( .A1(G567), .A2(n839), .ZN(n681) );
  NAND2_X1 U769 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U770 ( .A(KEYINPUT79), .B(n683), .ZN(G319) );
  INV_X1 U771 ( .A(G319), .ZN(n910) );
  NAND2_X1 U772 ( .A1(G661), .A2(G483), .ZN(n684) );
  NOR2_X1 U773 ( .A1(n910), .A2(n684), .ZN(n838) );
  NAND2_X1 U774 ( .A1(G36), .A2(n838), .ZN(n685) );
  XNOR2_X1 U775 ( .A(n685), .B(KEYINPUT80), .ZN(G176) );
  XNOR2_X1 U776 ( .A(G1986), .B(KEYINPUT84), .ZN(n686) );
  XNOR2_X1 U777 ( .A(n686), .B(G290), .ZN(n927) );
  NAND2_X1 U778 ( .A1(G160), .A2(G40), .ZN(n716) );
  NOR2_X1 U779 ( .A1(n718), .A2(n716), .ZN(n827) );
  NAND2_X1 U780 ( .A1(n927), .A2(n827), .ZN(n815) );
  NAND2_X1 U781 ( .A1(n882), .A2(G140), .ZN(n688) );
  NAND2_X1 U782 ( .A1(G104), .A2(n883), .ZN(n687) );
  NAND2_X1 U783 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U784 ( .A(KEYINPUT34), .B(n689), .ZN(n695) );
  NAND2_X1 U785 ( .A1(G116), .A2(n886), .ZN(n691) );
  NAND2_X1 U786 ( .A1(G128), .A2(n887), .ZN(n690) );
  NAND2_X1 U787 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U788 ( .A(KEYINPUT35), .B(n692), .ZN(n693) );
  XNOR2_X1 U789 ( .A(KEYINPUT85), .B(n693), .ZN(n694) );
  NOR2_X1 U790 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U791 ( .A(KEYINPUT36), .B(n696), .ZN(n905) );
  XNOR2_X1 U792 ( .A(G2067), .B(KEYINPUT37), .ZN(n825) );
  NOR2_X1 U793 ( .A1(n905), .A2(n825), .ZN(n975) );
  NAND2_X1 U794 ( .A1(n827), .A2(n975), .ZN(n823) );
  NAND2_X1 U795 ( .A1(G131), .A2(n882), .ZN(n698) );
  NAND2_X1 U796 ( .A1(G119), .A2(n887), .ZN(n697) );
  NAND2_X1 U797 ( .A1(n698), .A2(n697), .ZN(n702) );
  NAND2_X1 U798 ( .A1(n886), .A2(G107), .ZN(n700) );
  NAND2_X1 U799 ( .A1(G95), .A2(n883), .ZN(n699) );
  NAND2_X1 U800 ( .A1(n700), .A2(n699), .ZN(n701) );
  OR2_X1 U801 ( .A1(n702), .A2(n701), .ZN(n880) );
  NAND2_X1 U802 ( .A1(G1991), .A2(n880), .ZN(n712) );
  NAND2_X1 U803 ( .A1(G117), .A2(n886), .ZN(n704) );
  NAND2_X1 U804 ( .A1(G129), .A2(n887), .ZN(n703) );
  NAND2_X1 U805 ( .A1(n704), .A2(n703), .ZN(n707) );
  NAND2_X1 U806 ( .A1(G105), .A2(n883), .ZN(n705) );
  XOR2_X1 U807 ( .A(KEYINPUT38), .B(n705), .Z(n706) );
  NOR2_X1 U808 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U809 ( .A(n708), .B(KEYINPUT86), .ZN(n710) );
  NAND2_X1 U810 ( .A1(G141), .A2(n882), .ZN(n709) );
  NAND2_X1 U811 ( .A1(n710), .A2(n709), .ZN(n902) );
  NAND2_X1 U812 ( .A1(G1996), .A2(n902), .ZN(n711) );
  NAND2_X1 U813 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U814 ( .A(KEYINPUT87), .B(n713), .ZN(n990) );
  INV_X1 U815 ( .A(n990), .ZN(n714) );
  NAND2_X1 U816 ( .A1(n714), .A2(n827), .ZN(n816) );
  NAND2_X1 U817 ( .A1(n823), .A2(n816), .ZN(n715) );
  XNOR2_X1 U818 ( .A(n715), .B(KEYINPUT88), .ZN(n813) );
  INV_X1 U819 ( .A(n716), .ZN(n717) );
  NAND2_X2 U820 ( .A1(n718), .A2(n717), .ZN(n773) );
  NAND2_X1 U821 ( .A1(G8), .A2(n773), .ZN(n799) );
  NOR2_X1 U822 ( .A1(G1981), .A2(G305), .ZN(n719) );
  XNOR2_X1 U823 ( .A(n719), .B(KEYINPUT24), .ZN(n720) );
  XNOR2_X1 U824 ( .A(n720), .B(KEYINPUT89), .ZN(n721) );
  NOR2_X1 U825 ( .A1(n799), .A2(n721), .ZN(n722) );
  XNOR2_X1 U826 ( .A(n722), .B(KEYINPUT90), .ZN(n811) );
  NOR2_X1 U827 ( .A1(G2084), .A2(n773), .ZN(n758) );
  NAND2_X1 U828 ( .A1(G8), .A2(n758), .ZN(n772) );
  NOR2_X1 U829 ( .A1(G1966), .A2(n799), .ZN(n770) );
  XOR2_X1 U830 ( .A(n723), .B(KEYINPUT26), .Z(n725) );
  NAND2_X1 U831 ( .A1(n773), .A2(G1341), .ZN(n724) );
  INV_X1 U832 ( .A(n930), .ZN(n733) );
  AND2_X1 U833 ( .A1(n733), .A2(n919), .ZN(n726) );
  NAND2_X1 U834 ( .A1(n732), .A2(n726), .ZN(n730) );
  NOR2_X1 U835 ( .A1(n753), .A2(G1348), .ZN(n728) );
  NOR2_X1 U836 ( .A1(G2067), .A2(n773), .ZN(n727) );
  NOR2_X1 U837 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U838 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U839 ( .A(n731), .B(KEYINPUT95), .ZN(n736) );
  NOR2_X1 U840 ( .A1(n919), .A2(n734), .ZN(n735) );
  NOR2_X1 U841 ( .A1(n736), .A2(n735), .ZN(n738) );
  XNOR2_X1 U842 ( .A(n738), .B(n737), .ZN(n745) );
  NAND2_X1 U843 ( .A1(G1956), .A2(n773), .ZN(n739) );
  XNOR2_X1 U844 ( .A(KEYINPUT93), .B(n739), .ZN(n743) );
  XOR2_X1 U845 ( .A(KEYINPUT92), .B(KEYINPUT27), .Z(n741) );
  NAND2_X1 U846 ( .A1(n753), .A2(G2072), .ZN(n740) );
  XOR2_X1 U847 ( .A(n741), .B(n740), .Z(n742) );
  NOR2_X1 U848 ( .A1(n743), .A2(n742), .ZN(n747) );
  NAND2_X1 U849 ( .A1(n747), .A2(n746), .ZN(n744) );
  NAND2_X1 U850 ( .A1(n745), .A2(n744), .ZN(n751) );
  NOR2_X1 U851 ( .A1(n747), .A2(n746), .ZN(n749) );
  XOR2_X1 U852 ( .A(KEYINPUT94), .B(KEYINPUT28), .Z(n748) );
  XNOR2_X1 U853 ( .A(n749), .B(n748), .ZN(n750) );
  NAND2_X1 U854 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U855 ( .A(n752), .B(KEYINPUT29), .Z(n757) );
  XNOR2_X1 U856 ( .A(KEYINPUT91), .B(G1961), .ZN(n943) );
  NAND2_X1 U857 ( .A1(n773), .A2(n943), .ZN(n755) );
  XNOR2_X1 U858 ( .A(G2078), .B(KEYINPUT25), .ZN(n1001) );
  NAND2_X1 U859 ( .A1(n753), .A2(n1001), .ZN(n754) );
  NAND2_X1 U860 ( .A1(n755), .A2(n754), .ZN(n764) );
  NAND2_X1 U861 ( .A1(n764), .A2(G171), .ZN(n756) );
  NAND2_X1 U862 ( .A1(n757), .A2(n756), .ZN(n779) );
  NOR2_X1 U863 ( .A1(n770), .A2(n758), .ZN(n759) );
  NAND2_X1 U864 ( .A1(G8), .A2(n759), .ZN(n760) );
  XNOR2_X1 U865 ( .A(KEYINPUT98), .B(n760), .ZN(n762) );
  XOR2_X1 U866 ( .A(KEYINPUT30), .B(KEYINPUT97), .Z(n761) );
  XNOR2_X1 U867 ( .A(n762), .B(n761), .ZN(n763) );
  NOR2_X1 U868 ( .A1(G168), .A2(n763), .ZN(n767) );
  NOR2_X1 U869 ( .A1(G171), .A2(n764), .ZN(n765) );
  XOR2_X1 U870 ( .A(KEYINPUT99), .B(n765), .Z(n766) );
  NOR2_X1 U871 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U872 ( .A(KEYINPUT31), .B(n768), .Z(n777) );
  NAND2_X1 U873 ( .A1(n772), .A2(n771), .ZN(n787) );
  NOR2_X1 U874 ( .A1(G1971), .A2(n799), .ZN(n775) );
  NOR2_X1 U875 ( .A1(G2090), .A2(n773), .ZN(n774) );
  NOR2_X1 U876 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U877 ( .A1(n776), .A2(G303), .ZN(n780) );
  AND2_X1 U878 ( .A1(n777), .A2(n780), .ZN(n778) );
  NAND2_X1 U879 ( .A1(n779), .A2(n778), .ZN(n784) );
  INV_X1 U880 ( .A(n780), .ZN(n781) );
  OR2_X1 U881 ( .A1(n781), .A2(G286), .ZN(n782) );
  AND2_X1 U882 ( .A1(G8), .A2(n782), .ZN(n783) );
  NAND2_X1 U883 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U884 ( .A(KEYINPUT32), .B(n785), .ZN(n786) );
  NAND2_X1 U885 ( .A1(n787), .A2(n786), .ZN(n794) );
  NAND2_X1 U886 ( .A1(G166), .A2(G8), .ZN(n788) );
  OR2_X1 U887 ( .A1(G2090), .A2(n788), .ZN(n789) );
  NAND2_X1 U888 ( .A1(n794), .A2(n789), .ZN(n790) );
  NOR2_X1 U889 ( .A1(G1976), .A2(G288), .ZN(n797) );
  NOR2_X1 U890 ( .A1(G1971), .A2(G303), .ZN(n791) );
  NOR2_X1 U891 ( .A1(n797), .A2(n791), .ZN(n926) );
  INV_X1 U892 ( .A(KEYINPUT33), .ZN(n792) );
  AND2_X1 U893 ( .A1(n926), .A2(n792), .ZN(n793) );
  NAND2_X1 U894 ( .A1(n794), .A2(n793), .ZN(n805) );
  NAND2_X1 U895 ( .A1(G1976), .A2(G288), .ZN(n922) );
  INV_X1 U896 ( .A(n922), .ZN(n795) );
  NOR2_X1 U897 ( .A1(n795), .A2(n799), .ZN(n796) );
  NOR2_X1 U898 ( .A1(KEYINPUT33), .A2(n796), .ZN(n801) );
  NAND2_X1 U899 ( .A1(n797), .A2(KEYINPUT33), .ZN(n798) );
  NOR2_X1 U900 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U901 ( .A1(n801), .A2(n800), .ZN(n803) );
  XOR2_X1 U902 ( .A(G1981), .B(KEYINPUT100), .Z(n802) );
  XNOR2_X1 U903 ( .A(G305), .B(n802), .ZN(n915) );
  AND2_X1 U904 ( .A1(n803), .A2(n915), .ZN(n804) );
  NAND2_X1 U905 ( .A1(n805), .A2(n804), .ZN(n807) );
  NAND2_X1 U906 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n830) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n902), .ZN(n979) );
  INV_X1 U911 ( .A(n816), .ZN(n820) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n880), .ZN(n971) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n817) );
  NOR2_X1 U914 ( .A1(n971), .A2(n817), .ZN(n818) );
  XOR2_X1 U915 ( .A(KEYINPUT103), .B(n818), .Z(n819) );
  NOR2_X1 U916 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U917 ( .A1(n979), .A2(n821), .ZN(n822) );
  XNOR2_X1 U918 ( .A(n822), .B(KEYINPUT39), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n826) );
  NAND2_X1 U920 ( .A1(n905), .A2(n825), .ZN(n976) );
  NAND2_X1 U921 ( .A1(n826), .A2(n976), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n830), .A2(n829), .ZN(n832) );
  XNOR2_X1 U924 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n831) );
  XNOR2_X1 U925 ( .A(n832), .B(n831), .ZN(G329) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n833), .ZN(G217) );
  NAND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n835) );
  INV_X1 U928 ( .A(G661), .ZN(n834) );
  NOR2_X1 U929 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U930 ( .A(n836), .B(KEYINPUT107), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U932 ( .A1(n838), .A2(n837), .ZN(G188) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NOR2_X1 U937 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U939 ( .A(n930), .B(KEYINPUT113), .ZN(n842) );
  XNOR2_X1 U940 ( .A(G171), .B(n919), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n845) );
  XOR2_X1 U942 ( .A(G286), .B(n843), .Z(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n846) );
  NOR2_X1 U944 ( .A1(G37), .A2(n846), .ZN(G397) );
  XOR2_X1 U945 ( .A(G2100), .B(KEYINPUT109), .Z(n848) );
  XNOR2_X1 U946 ( .A(KEYINPUT108), .B(G2678), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U948 ( .A(KEYINPUT42), .B(G2090), .Z(n850) );
  XNOR2_X1 U949 ( .A(G2067), .B(G2072), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U951 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U952 ( .A(KEYINPUT43), .B(G2096), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(n856) );
  XOR2_X1 U954 ( .A(G2078), .B(G2084), .Z(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(G227) );
  XOR2_X1 U956 ( .A(G1971), .B(G1956), .Z(n858) );
  XNOR2_X1 U957 ( .A(G1966), .B(G1961), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U959 ( .A(n859), .B(G2474), .Z(n861) );
  XNOR2_X1 U960 ( .A(G1986), .B(G1976), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U962 ( .A(KEYINPUT41), .B(G1981), .Z(n863) );
  XNOR2_X1 U963 ( .A(G1996), .B(G1991), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n865), .B(n864), .ZN(G229) );
  NAND2_X1 U966 ( .A1(G124), .A2(n887), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n866), .B(KEYINPUT44), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n886), .A2(G112), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U970 ( .A1(n882), .A2(G136), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G100), .A2(n883), .ZN(n869) );
  NAND2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U973 ( .A1(n872), .A2(n871), .ZN(G162) );
  NAND2_X1 U974 ( .A1(G118), .A2(n886), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G130), .A2(n887), .ZN(n873) );
  NAND2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n879) );
  NAND2_X1 U977 ( .A1(n882), .A2(G142), .ZN(n876) );
  NAND2_X1 U978 ( .A1(G106), .A2(n883), .ZN(n875) );
  NAND2_X1 U979 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U980 ( .A(n877), .B(KEYINPUT45), .Z(n878) );
  NOR2_X1 U981 ( .A1(n879), .A2(n878), .ZN(n881) );
  XNOR2_X1 U982 ( .A(n881), .B(n880), .ZN(n901) );
  NAND2_X1 U983 ( .A1(n882), .A2(G139), .ZN(n885) );
  NAND2_X1 U984 ( .A1(G103), .A2(n883), .ZN(n884) );
  NAND2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n893) );
  NAND2_X1 U986 ( .A1(G115), .A2(n886), .ZN(n889) );
  NAND2_X1 U987 ( .A1(G127), .A2(n887), .ZN(n888) );
  NAND2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U989 ( .A(KEYINPUT110), .B(n890), .Z(n891) );
  XNOR2_X1 U990 ( .A(KEYINPUT47), .B(n891), .ZN(n892) );
  NOR2_X1 U991 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U992 ( .A(KEYINPUT111), .B(n894), .ZN(n981) );
  XOR2_X1 U993 ( .A(KEYINPUT48), .B(KEYINPUT112), .Z(n896) );
  XNOR2_X1 U994 ( .A(G162), .B(KEYINPUT46), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n981), .B(n897), .ZN(n899) );
  XNOR2_X1 U997 ( .A(G164), .B(G160), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(n902), .B(n970), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n907), .ZN(G395) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1006 ( .A1(G397), .A2(n909), .ZN(n914) );
  NOR2_X1 U1007 ( .A1(n910), .A2(G401), .ZN(n911) );
  XOR2_X1 U1008 ( .A(KEYINPUT114), .B(n911), .Z(n912) );
  NOR2_X1 U1009 ( .A1(G395), .A2(n912), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1013 ( .A(G1966), .B(G168), .ZN(n916) );
  NAND2_X1 U1014 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(n917), .B(KEYINPUT57), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(KEYINPUT121), .B(n918), .ZN(n940) );
  XNOR2_X1 U1017 ( .A(G1348), .B(n919), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(n920), .B(KEYINPUT122), .ZN(n935) );
  NAND2_X1 U1019 ( .A1(G1971), .A2(G303), .ZN(n921) );
  NAND2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n924) );
  XNOR2_X1 U1021 ( .A(G1956), .B(G299), .ZN(n923) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n928) );
  NOR2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1025 ( .A(n929), .B(KEYINPUT123), .ZN(n933) );
  XNOR2_X1 U1026 ( .A(G1341), .B(n930), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(KEYINPUT124), .B(n931), .ZN(n932) );
  NOR2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n937) );
  XOR2_X1 U1030 ( .A(G171), .B(G1961), .Z(n936) );
  NOR2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(KEYINPUT125), .B(n938), .ZN(n939) );
  NOR2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n942) );
  XOR2_X1 U1034 ( .A(G16), .B(KEYINPUT56), .Z(n941) );
  NOR2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n969) );
  XOR2_X1 U1036 ( .A(G16), .B(KEYINPUT126), .Z(n966) );
  XNOR2_X1 U1037 ( .A(G5), .B(n943), .ZN(n961) );
  XOR2_X1 U1038 ( .A(G1348), .B(KEYINPUT59), .Z(n944) );
  XNOR2_X1 U1039 ( .A(G4), .B(n944), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(G20), .B(G1956), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(G1341), .B(G19), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(G1981), .B(G6), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(n951), .B(KEYINPUT60), .ZN(n959) );
  XNOR2_X1 U1047 ( .A(G1986), .B(G24), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(G22), .B(G1971), .ZN(n952) );
  NOR2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(G1976), .B(KEYINPUT127), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(n954), .B(G23), .ZN(n955) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(KEYINPUT58), .B(n957), .ZN(n958) );
  NOR2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(G21), .B(G1966), .ZN(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(n964), .B(KEYINPUT61), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(G11), .A2(n967), .ZN(n968) );
  NOR2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n998) );
  XNOR2_X1 U1062 ( .A(G160), .B(G2084), .ZN(n973) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n977) );
  NAND2_X1 U1066 ( .A1(n977), .A2(n976), .ZN(n992) );
  XOR2_X1 U1067 ( .A(G2090), .B(G162), .Z(n978) );
  NOR2_X1 U1068 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(KEYINPUT51), .B(n980), .ZN(n988) );
  XNOR2_X1 U1070 ( .A(G164), .B(G2078), .ZN(n984) );
  XNOR2_X1 U1071 ( .A(G2072), .B(KEYINPUT115), .ZN(n982) );
  XNOR2_X1 U1072 ( .A(n982), .B(n981), .ZN(n983) );
  NAND2_X1 U1073 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(n985), .B(KEYINPUT116), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(KEYINPUT50), .B(n986), .ZN(n987) );
  NOR2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1077 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1078 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1079 ( .A(n993), .B(KEYINPUT52), .ZN(n994) );
  XNOR2_X1 U1080 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n1017) );
  NAND2_X1 U1081 ( .A1(n994), .A2(n1017), .ZN(n995) );
  XNOR2_X1 U1082 ( .A(KEYINPUT118), .B(n995), .ZN(n996) );
  NAND2_X1 U1083 ( .A1(n996), .A2(G29), .ZN(n997) );
  NAND2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n1021) );
  XNOR2_X1 U1085 ( .A(KEYINPUT119), .B(G2067), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(n999), .B(G26), .ZN(n1009) );
  XOR2_X1 U1087 ( .A(G2072), .B(G33), .Z(n1000) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(G28), .ZN(n1007) );
  XNOR2_X1 U1089 ( .A(G27), .B(n1001), .ZN(n1005) );
  XNOR2_X1 U1090 ( .A(G1996), .B(G32), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(G1991), .B(G25), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(n1010), .B(KEYINPUT120), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(n1011), .B(KEYINPUT53), .ZN(n1014) );
  XOR2_X1 U1098 ( .A(G2084), .B(G34), .Z(n1012) );
  XNOR2_X1 U1099 ( .A(KEYINPUT54), .B(n1012), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XNOR2_X1 U1101 ( .A(G35), .B(G2090), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XNOR2_X1 U1103 ( .A(n1018), .B(n1017), .ZN(n1019) );
  NOR2_X1 U1104 ( .A1(G29), .A2(n1019), .ZN(n1020) );
  NOR2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1106 ( .A(n1022), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

