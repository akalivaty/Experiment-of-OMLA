//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n785, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n207));
  INV_X1    g006(.A(G113gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(G120gat), .ZN(new_n209));
  INV_X1    g008(.A(G120gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(G113gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n207), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G134gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G127gat), .ZN(new_n214));
  INV_X1    g013(.A(G127gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G134gat), .ZN(new_n216));
  AND3_X1   g015(.A1(new_n214), .A2(new_n216), .A3(KEYINPUT68), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT68), .B1(new_n214), .B2(new_n216), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n212), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT69), .ZN(new_n220));
  XNOR2_X1  g019(.A(G127gat), .B(G134gat), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n221), .B(new_n207), .C1(new_n209), .C2(new_n211), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT69), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n223), .B(new_n212), .C1(new_n217), .C2(new_n218), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n220), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT74), .B1(G155gat), .B2(G162gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(G141gat), .B(G148gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n228), .B1(G155gat), .B2(G162gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n226), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G155gat), .B(G162gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G155gat), .A2(G162gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT2), .ZN(new_n235));
  INV_X1    g034(.A(G141gat), .ZN(new_n236));
  INV_X1    g035(.A(G148gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G141gat), .A2(G148gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n235), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(new_n231), .A3(new_n226), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n233), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n225), .B(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G225gat), .A2(G233gat), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT5), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n233), .A2(KEYINPUT77), .A3(new_n241), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT77), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n240), .A2(new_n231), .A3(new_n226), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n231), .B1(new_n240), .B2(new_n226), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n225), .B1(new_n246), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT78), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n224), .A2(new_n222), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n221), .A2(KEYINPUT68), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n215), .A2(G134gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n213), .A2(G127gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n223), .B1(new_n260), .B2(new_n212), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n250), .A2(new_n246), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n252), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT78), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n262), .A2(new_n252), .A3(new_n242), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n253), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n244), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT75), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT3), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n270), .B1(new_n242), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n248), .A2(new_n249), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n262), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT76), .B1(new_n273), .B2(KEYINPUT3), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT76), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n242), .A2(new_n277), .A3(new_n271), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n269), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n245), .B1(new_n268), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n262), .A2(new_n263), .A3(new_n252), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT4), .B1(new_n225), .B2(new_n273), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT5), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n280), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  OAI211_X1 g085(.A(KEYINPUT6), .B(new_n206), .C1(new_n281), .C2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT79), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n267), .B1(new_n264), .B2(new_n265), .ZN(new_n290));
  AOI211_X1 g089(.A(KEYINPUT78), .B(new_n252), .C1(new_n262), .C2(new_n263), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n280), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n245), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(new_n285), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n295), .A2(KEYINPUT79), .A3(KEYINPUT6), .A4(new_n206), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT6), .B1(new_n295), .B2(new_n206), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n292), .A2(new_n293), .B1(new_n280), .B2(new_n284), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n205), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n289), .A2(new_n296), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT91), .ZN(new_n301));
  INV_X1    g100(.A(G169gat), .ZN(new_n302));
  INV_X1    g101(.A(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT26), .ZN(new_n305));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(KEYINPUT66), .ZN(new_n307));
  NOR2_X1   g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT66), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n305), .B(new_n306), .C1(new_n311), .C2(KEYINPUT26), .ZN(new_n312));
  XOR2_X1   g111(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT27), .B(G183gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n313), .B1(new_n315), .B2(G190gat), .ZN(new_n316));
  INV_X1    g115(.A(G190gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n314), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G183gat), .A2(G190gat), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n312), .A2(new_n316), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(G183gat), .A2(G190gat), .ZN(new_n322));
  AND2_X1   g121(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n322), .B1(new_n323), .B2(G190gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT24), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n307), .A2(KEYINPUT23), .A3(new_n310), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT25), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n306), .A2(KEYINPUT23), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n329), .B1(new_n330), .B2(new_n304), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n327), .A2(new_n328), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT64), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n326), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n320), .A2(KEYINPUT64), .A3(new_n325), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n324), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT23), .ZN(new_n337));
  NOR3_X1   g136(.A1(new_n337), .A2(G169gat), .A3(G176gat), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(new_n304), .B2(new_n330), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT25), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT65), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n332), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AOI211_X1 g141(.A(KEYINPUT65), .B(KEYINPUT25), .C1(new_n336), .C2(new_n339), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n321), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n262), .ZN(new_n345));
  INV_X1    g144(.A(G227gat), .ZN(new_n346));
  INV_X1    g145(.A(G233gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n225), .B(new_n321), .C1(new_n342), .C2(new_n343), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n345), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT32), .ZN(new_n351));
  XNOR2_X1  g150(.A(G15gat), .B(G43gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT70), .ZN(new_n353));
  XNOR2_X1  g152(.A(G71gat), .B(G99gat), .ZN(new_n354));
  XOR2_X1   g153(.A(new_n353), .B(new_n354), .Z(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n351), .B1(KEYINPUT33), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n355), .B1(new_n350), .B2(KEYINPUT32), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT71), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT33), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n350), .A2(new_n361), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n360), .B1(new_n359), .B2(new_n362), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n358), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n330), .A2(new_n304), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n308), .A2(KEYINPUT23), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n369), .B1(G183gat), .B2(G190gat), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT64), .B1(new_n320), .B2(new_n325), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n368), .B1(new_n335), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT65), .B1(new_n373), .B2(KEYINPUT25), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n340), .A2(new_n341), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(new_n375), .A3(new_n332), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n225), .B1(new_n376), .B2(new_n321), .ZN(new_n377));
  INV_X1    g176(.A(new_n349), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT34), .B1(new_n379), .B2(new_n348), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT34), .ZN(new_n381));
  OAI221_X1 g180(.A(new_n381), .B1(new_n346), .B2(new_n347), .C1(new_n377), .C2(new_n378), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n365), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n351), .A2(new_n362), .A3(new_n356), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT71), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n383), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(new_n389), .A3(new_n358), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT81), .B(G22gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G78gat), .B(G106gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT31), .B(G50gat), .ZN(new_n394));
  XOR2_X1   g193(.A(new_n393), .B(new_n394), .Z(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n397));
  XNOR2_X1  g196(.A(G197gat), .B(G204gat), .ZN(new_n398));
  INV_X1    g197(.A(G211gat), .ZN(new_n399));
  INV_X1    g198(.A(G218gat), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n398), .B1(KEYINPUT22), .B2(new_n401), .ZN(new_n402));
  XOR2_X1   g201(.A(G211gat), .B(G218gat), .Z(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT29), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT3), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n406), .A2(new_n263), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n273), .A2(KEYINPUT76), .A3(KEYINPUT3), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n277), .B1(new_n242), .B2(new_n271), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n405), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n404), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n407), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G228gat), .A2(G233gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n397), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT29), .B1(new_n276), .B2(new_n278), .ZN(new_n416));
  OAI22_X1  g215(.A1(new_n416), .A2(new_n404), .B1(new_n263), .B2(new_n406), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n417), .A2(KEYINPUT80), .A3(new_n413), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n416), .A2(new_n404), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n414), .B1(new_n406), .B2(new_n242), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n396), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  AOI211_X1 g223(.A(new_n395), .B(new_n422), .C1(new_n415), .C2(new_n418), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n392), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n412), .A2(new_n397), .A3(new_n414), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT80), .B1(new_n417), .B2(new_n413), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n423), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n395), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n419), .A2(new_n396), .A3(new_n423), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n391), .A3(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n384), .A2(new_n390), .A3(new_n426), .A4(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(G8gat), .B(G36gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n435), .B(KEYINPUT72), .ZN(new_n436));
  XNOR2_X1  g235(.A(G64gat), .B(G92gat), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n436), .B(new_n437), .Z(new_n438));
  NAND2_X1  g237(.A1(G226gat), .A2(G233gat), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n321), .B(new_n439), .C1(new_n342), .C2(new_n343), .ZN(new_n440));
  AND4_X1   g239(.A1(new_n312), .A2(new_n316), .A3(new_n319), .A4(new_n320), .ZN(new_n441));
  INV_X1    g240(.A(new_n332), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n336), .A2(new_n339), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n329), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n444), .B2(KEYINPUT65), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n441), .B1(new_n445), .B2(new_n375), .ZN(new_n446));
  INV_X1    g245(.A(new_n439), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n447), .A2(KEYINPUT29), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n404), .B(new_n440), .C1(new_n446), .C2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n344), .B1(KEYINPUT29), .B2(new_n447), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n404), .B1(new_n451), .B2(new_n440), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n438), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n440), .B1(new_n446), .B2(new_n448), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n411), .ZN(new_n455));
  INV_X1    g254(.A(new_n438), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n455), .A2(KEYINPUT30), .A3(new_n449), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT73), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n453), .A2(new_n457), .A3(KEYINPUT73), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n455), .A2(new_n449), .A3(new_n456), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT30), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n460), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n289), .A2(new_n296), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n206), .B1(new_n281), .B2(new_n286), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n299), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n465), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n434), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n464), .A2(new_n453), .A3(new_n457), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n300), .A2(KEYINPUT35), .A3(new_n472), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n471), .A2(KEYINPUT35), .B1(new_n473), .B2(new_n434), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT40), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n275), .A2(new_n279), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n282), .A2(new_n283), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(KEYINPUT83), .B(KEYINPUT39), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n269), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n205), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n243), .A2(new_n244), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT39), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(new_n269), .B2(new_n478), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n475), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n478), .A2(new_n269), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n486), .A2(KEYINPUT39), .A3(new_n482), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n487), .A2(KEYINPUT40), .A3(new_n205), .A4(new_n480), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n472), .A2(new_n485), .A3(new_n488), .A4(new_n467), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n489), .A2(new_n432), .A3(new_n426), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n205), .B1(new_n294), .B2(new_n285), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT79), .B1(new_n491), .B2(KEYINPUT6), .ZN(new_n492));
  NOR4_X1   g291(.A1(new_n298), .A2(new_n288), .A3(new_n468), .A4(new_n205), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n469), .B(new_n462), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n450), .A2(new_n452), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT37), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n456), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n450), .A2(KEYINPUT84), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT84), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n449), .A2(new_n500), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n499), .A2(new_n452), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n498), .B1(new_n502), .B2(new_n497), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT38), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n496), .A2(new_n497), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n505), .A2(new_n504), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n503), .A2(new_n504), .B1(new_n498), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n490), .B1(new_n495), .B2(new_n508), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n384), .A2(new_n390), .A3(KEYINPUT36), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT36), .B1(new_n384), .B2(new_n390), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n426), .A2(new_n432), .ZN(new_n512));
  OAI22_X1  g311(.A1(new_n510), .A2(new_n511), .B1(new_n470), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n509), .B1(new_n513), .B2(KEYINPUT82), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT36), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n389), .B1(new_n388), .B2(new_n358), .ZN(new_n516));
  AOI211_X1 g315(.A(new_n383), .B(new_n357), .C1(new_n386), .C2(new_n387), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n384), .A2(new_n390), .A3(KEYINPUT36), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n426), .A2(new_n432), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(new_n300), .B2(new_n465), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT82), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n520), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n474), .B1(new_n514), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT90), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT18), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G29gat), .ZN(new_n529));
  INV_X1    g328(.A(G36gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT14), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT14), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(G29gat), .B2(G36gat), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n531), .B(new_n533), .C1(new_n529), .C2(new_n530), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT15), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G43gat), .B(G50gat), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n534), .A2(new_n535), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n539), .A3(new_n537), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(KEYINPUT87), .B(KEYINPUT17), .Z(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT88), .ZN(new_n544));
  XNOR2_X1  g343(.A(G15gat), .B(G22gat), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n545), .A2(G1gat), .ZN(new_n546));
  AOI21_X1  g345(.A(G8gat), .B1(new_n546), .B2(KEYINPUT89), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT16), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n545), .B1(new_n548), .B2(G1gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n547), .B(new_n550), .Z(new_n551));
  INV_X1    g350(.A(new_n541), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n551), .B1(KEYINPUT17), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n544), .A2(new_n553), .B1(new_n551), .B2(new_n541), .ZN(new_n554));
  NAND2_X1  g353(.A1(G229gat), .A2(G233gat), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n528), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n543), .A2(KEYINPUT88), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT88), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n558), .B1(new_n541), .B2(new_n542), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n553), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n551), .A2(new_n541), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n560), .A2(new_n555), .A3(new_n561), .A4(new_n528), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n547), .B(new_n550), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n552), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n555), .B(KEYINPUT13), .Z(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT86), .B1(new_n556), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G113gat), .B(G141gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G169gat), .B(G197gat), .Z(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT12), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(KEYINPUT86), .B(new_n575), .C1(new_n556), .C2(new_n568), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n301), .B1(new_n525), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n579), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n520), .A2(new_n523), .A3(new_n522), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n523), .B1(new_n520), .B2(new_n522), .ZN(new_n583));
  NOR3_X1   g382(.A1(new_n582), .A2(new_n583), .A3(new_n509), .ZN(new_n584));
  OAI211_X1 g383(.A(KEYINPUT91), .B(new_n581), .C1(new_n584), .C2(new_n474), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  AND2_X1   g385(.A1(G232gat), .A2(G233gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n587), .A2(KEYINPUT41), .ZN(new_n588));
  XNOR2_X1  g387(.A(G134gat), .B(G162gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT7), .ZN(new_n592));
  NAND2_X1  g391(.A1(G99gat), .A2(G106gat), .ZN(new_n593));
  INV_X1    g392(.A(G85gat), .ZN(new_n594));
  INV_X1    g393(.A(G92gat), .ZN(new_n595));
  AOI22_X1  g394(.A1(KEYINPUT8), .A2(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G99gat), .B(G106gat), .Z(new_n598));
  AOI21_X1  g397(.A(new_n597), .B1(KEYINPUT94), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n598), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT94), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n597), .A2(new_n601), .A3(new_n600), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n605), .B1(new_n552), .B2(KEYINPUT17), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n606), .B1(new_n557), .B2(new_n559), .ZN(new_n607));
  AOI22_X1  g406(.A1(new_n605), .A2(new_n541), .B1(KEYINPUT41), .B2(new_n587), .ZN(new_n608));
  XNOR2_X1  g407(.A(G190gat), .B(G218gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT95), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n610), .B1(new_n607), .B2(new_n608), .ZN(new_n613));
  OAI211_X1 g412(.A(KEYINPUT96), .B(new_n590), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n613), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n590), .A2(KEYINPUT96), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n590), .A2(KEYINPUT96), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .A4(new_n611), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G57gat), .B(G64gat), .Z(new_n620));
  INV_X1    g419(.A(KEYINPUT9), .ZN(new_n621));
  INV_X1    g420(.A(G71gat), .ZN(new_n622));
  INV_X1    g421(.A(G78gat), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G71gat), .B(G78gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(KEYINPUT21), .ZN(new_n628));
  XNOR2_X1  g427(.A(G127gat), .B(G155gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT21), .ZN(new_n631));
  INV_X1    g430(.A(new_n627), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n563), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n630), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G231gat), .A2(G233gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n635), .B(KEYINPUT93), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT92), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G183gat), .B(G211gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n634), .B(new_n641), .Z(new_n642));
  NAND2_X1  g441(.A1(new_n619), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(KEYINPUT97), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n619), .A2(new_n645), .A3(new_n642), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n603), .A3(new_n604), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT98), .B1(new_n592), .B2(new_n596), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n651), .A2(new_n598), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n627), .B1(new_n598), .B2(new_n651), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n649), .B(new_n650), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n605), .A2(KEYINPUT10), .A3(new_n627), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n648), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n653), .A2(new_n652), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n647), .B1(new_n657), .B2(new_n649), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G120gat), .B(G148gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(G176gat), .B(G204gat), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n660), .B(new_n661), .Z(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n656), .A2(new_n658), .A3(new_n663), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n664), .A2(KEYINPUT99), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT99), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n659), .A2(new_n668), .A3(new_n663), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n644), .A2(new_n646), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT100), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT100), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n644), .A2(new_n673), .A3(new_n646), .A4(new_n670), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT101), .B1(new_n586), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n678));
  AOI211_X1 g477(.A(new_n678), .B(new_n675), .C1(new_n580), .C2(new_n585), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n300), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g480(.A(KEYINPUT102), .B(KEYINPUT16), .ZN(new_n682));
  INV_X1    g481(.A(G8gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n472), .B(new_n684), .C1(new_n677), .C2(new_n679), .ZN(new_n685));
  INV_X1    g484(.A(new_n472), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n513), .A2(KEYINPUT82), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n512), .B(new_n489), .C1(new_n494), .C2(new_n507), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(new_n524), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n466), .A2(new_n469), .ZN(new_n690));
  INV_X1    g489(.A(new_n465), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT35), .B1(new_n692), .B2(new_n433), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n473), .A2(new_n434), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT91), .B1(new_n696), .B2(new_n581), .ZN(new_n697));
  AOI211_X1 g496(.A(new_n301), .B(new_n579), .C1(new_n689), .C2(new_n695), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n676), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(new_n678), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n586), .A2(KEYINPUT101), .A3(new_n676), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n686), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n685), .B1(new_n702), .B2(new_n683), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT42), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n685), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(G1325gat));
  NOR2_X1   g506(.A1(new_n677), .A2(new_n679), .ZN(new_n708));
  OAI21_X1  g507(.A(G15gat), .B1(new_n708), .B2(new_n520), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n516), .A2(new_n517), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n711), .A2(G15gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n709), .B1(new_n708), .B2(new_n712), .ZN(G1326gat));
  NOR2_X1   g512(.A1(new_n708), .A2(new_n512), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT43), .B(G22gat), .Z(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  INV_X1    g515(.A(new_n619), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n696), .A2(KEYINPUT44), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n688), .A2(new_n520), .A3(new_n522), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n619), .B1(new_n695), .B2(new_n719), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n720), .A2(KEYINPUT44), .ZN(new_n721));
  INV_X1    g520(.A(new_n670), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(new_n642), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n581), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n718), .A2(new_n721), .A3(new_n725), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n726), .A2(new_n690), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n723), .A2(new_n717), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(new_n580), .B2(new_n585), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n729), .A2(new_n529), .A3(new_n300), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n731));
  AOI22_X1  g530(.A1(G29gat), .A2(new_n727), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n731), .B2(new_n730), .ZN(G1328gat));
  INV_X1    g532(.A(new_n729), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n472), .A2(new_n530), .ZN(new_n735));
  OR3_X1    g534(.A1(new_n734), .A2(KEYINPUT46), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(G36gat), .B1(new_n726), .B2(new_n686), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT46), .B1(new_n734), .B2(new_n735), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(G1329gat));
  NOR2_X1   g538(.A1(new_n734), .A2(new_n711), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(G43gat), .ZN(new_n741));
  INV_X1    g540(.A(new_n520), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G43gat), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n726), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT47), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT47), .ZN(new_n746));
  OAI221_X1 g545(.A(new_n746), .B1(new_n726), .B2(new_n743), .C1(new_n740), .C2(G43gat), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1330gat));
  INV_X1    g547(.A(KEYINPUT104), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n718), .A2(new_n721), .A3(new_n521), .A4(new_n725), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G50gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT48), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT103), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n512), .A2(G50gat), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n753), .B1(new_n729), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n729), .A2(new_n753), .A3(new_n754), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n749), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n729), .A2(new_n754), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT103), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT48), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(new_n750), .B2(G50gat), .ZN(new_n762));
  AND4_X1   g561(.A1(new_n749), .A2(new_n760), .A3(new_n757), .A4(new_n762), .ZN(new_n763));
  AOI22_X1  g562(.A1(new_n729), .A2(new_n754), .B1(new_n750), .B2(G50gat), .ZN(new_n764));
  OAI22_X1  g563(.A1(new_n758), .A2(new_n763), .B1(KEYINPUT48), .B2(new_n764), .ZN(G1331gat));
  NAND2_X1  g564(.A1(new_n695), .A2(new_n719), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n644), .A2(new_n646), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n767), .A2(new_n579), .A3(new_n722), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n300), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g571(.A1(new_n769), .A2(new_n686), .ZN(new_n773));
  NOR2_X1   g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  AND2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n773), .B2(new_n774), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT105), .ZN(G1333gat));
  NAND3_X1  g577(.A1(new_n770), .A2(G71gat), .A3(new_n742), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n769), .A2(new_n711), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n780), .A2(KEYINPUT106), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n622), .B1(new_n780), .B2(KEYINPUT106), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n779), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n512), .ZN(new_n785));
  XNOR2_X1  g584(.A(KEYINPUT107), .B(G78gat), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1335gat));
  NAND2_X1  g586(.A1(new_n718), .A2(new_n721), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n581), .A2(new_n642), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n722), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(G85gat), .B1(new_n791), .B2(new_n690), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n720), .A2(new_n789), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n793), .A2(KEYINPUT51), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(KEYINPUT51), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(new_n722), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n300), .A2(new_n594), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n792), .B1(new_n796), .B2(new_n797), .ZN(G1336gat));
  OAI21_X1  g597(.A(G92gat), .B1(new_n791), .B2(new_n686), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n686), .A2(G92gat), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n794), .A2(new_n722), .A3(new_n795), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n801), .B2(KEYINPUT108), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n802), .B(new_n804), .ZN(G1337gat));
  NOR2_X1   g604(.A1(new_n796), .A2(new_n711), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n742), .A2(G99gat), .ZN(new_n807));
  OAI22_X1  g606(.A1(new_n806), .A2(G99gat), .B1(new_n791), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(KEYINPUT109), .ZN(G1338gat));
  NOR2_X1   g608(.A1(new_n791), .A2(new_n512), .ZN(new_n810));
  INV_X1    g609(.A(G106gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n521), .A2(new_n811), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n810), .A2(new_n811), .B1(new_n796), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT53), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815));
  OAI221_X1 g614(.A(new_n815), .B1(new_n796), .B2(new_n812), .C1(new_n810), .C2(new_n811), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(G1339gat));
  INV_X1    g616(.A(new_n642), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n656), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n654), .A2(new_n655), .A3(KEYINPUT110), .A4(new_n648), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT110), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n654), .A2(new_n655), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(new_n647), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n820), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826));
  AOI211_X1 g625(.A(new_n826), .B(new_n662), .C1(new_n656), .C2(new_n819), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n666), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n662), .B1(new_n656), .B2(new_n819), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT55), .B1(new_n825), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(new_n577), .A3(new_n578), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n560), .A2(new_n555), .A3(new_n561), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n526), .A3(new_n527), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n835), .A2(new_n567), .A3(new_n562), .A4(new_n575), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n554), .A2(new_n555), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n565), .A2(new_n566), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n574), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n836), .A2(new_n839), .A3(new_n669), .A4(new_n667), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n717), .B1(new_n833), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n832), .A2(new_n717), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n836), .A2(new_n839), .A3(KEYINPUT111), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT111), .B1(new_n836), .B2(new_n839), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n818), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n767), .A2(new_n579), .A3(new_n670), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n433), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(new_n300), .A3(new_n686), .ZN(new_n849));
  XOR2_X1   g648(.A(new_n849), .B(KEYINPUT112), .Z(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n208), .A3(new_n581), .ZN(new_n851));
  OAI21_X1  g650(.A(G113gat), .B1(new_n849), .B2(new_n579), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1340gat));
  NOR2_X1   g652(.A1(new_n670), .A2(G120gat), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT113), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(G120gat), .B1(new_n849), .B2(new_n670), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1341gat));
  NOR2_X1   g657(.A1(new_n849), .A2(new_n818), .ZN(new_n859));
  XNOR2_X1  g658(.A(KEYINPUT114), .B(G127gat), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n859), .B(new_n860), .ZN(G1342gat));
  NAND2_X1  g660(.A1(new_n717), .A2(new_n686), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n690), .B1(new_n862), .B2(KEYINPUT115), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(KEYINPUT115), .B2(new_n862), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(G134gat), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n848), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(KEYINPUT56), .Z(new_n867));
  OAI21_X1  g666(.A(G134gat), .B1(new_n849), .B2(new_n619), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1343gat));
  NAND2_X1  g668(.A1(new_n846), .A2(new_n847), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n871), .A3(new_n521), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n300), .A2(new_n686), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n742), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT116), .B1(new_n829), .B2(new_n831), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n665), .B1(new_n825), .B2(new_n827), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n825), .A2(new_n830), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n876), .B(new_n877), .C1(new_n878), .C2(KEYINPUT55), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n875), .A2(new_n879), .A3(new_n577), .A4(new_n578), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n717), .B1(new_n880), .B2(new_n840), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n818), .B1(new_n881), .B2(new_n845), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n512), .B1(new_n882), .B2(new_n847), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n872), .B(new_n874), .C1(new_n871), .C2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(G141gat), .B1(new_n884), .B2(new_n579), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n521), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n886), .A2(new_n742), .A3(new_n873), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n581), .A2(new_n236), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT117), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n890));
  AOI22_X1  g689(.A1(new_n887), .A2(new_n889), .B1(new_n890), .B2(KEYINPUT58), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n885), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n890), .A2(KEYINPUT58), .ZN(new_n893));
  XOR2_X1   g692(.A(new_n892), .B(new_n893), .Z(G1344gat));
  NAND3_X1  g693(.A1(new_n887), .A2(new_n237), .A3(new_n722), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n870), .A2(KEYINPUT57), .A3(new_n521), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT119), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT119), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n870), .A2(new_n899), .A3(KEYINPUT57), .A4(new_n521), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n672), .A2(new_n579), .A3(new_n674), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n882), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT120), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n512), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n882), .A2(new_n903), .A3(KEYINPUT120), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n871), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n902), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n722), .A3(new_n874), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n896), .B1(new_n911), .B2(G148gat), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n884), .A2(new_n670), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n913), .A2(KEYINPUT59), .A3(new_n237), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n895), .B1(new_n912), .B2(new_n914), .ZN(G1345gat));
  OAI21_X1  g714(.A(G155gat), .B1(new_n884), .B2(new_n818), .ZN(new_n916));
  INV_X1    g715(.A(G155gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n887), .A2(new_n917), .A3(new_n642), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1346gat));
  OR4_X1    g718(.A1(G162gat), .A2(new_n886), .A3(new_n742), .A4(new_n864), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT121), .B1(new_n884), .B2(new_n619), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G162gat), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n884), .A2(KEYINPUT121), .A3(new_n619), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(G1347gat));
  NAND4_X1  g723(.A1(new_n870), .A2(new_n690), .A3(new_n434), .A4(new_n472), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n925), .A2(new_n302), .A3(new_n579), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n925), .B(KEYINPUT122), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n581), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n926), .B1(new_n928), .B2(new_n302), .ZN(G1348gat));
  AOI21_X1  g728(.A(G176gat), .B1(new_n927), .B2(new_n722), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n930), .A2(KEYINPUT123), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n930), .A2(KEYINPUT123), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n925), .A2(new_n303), .A3(new_n670), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT124), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(G1349gat));
  NOR2_X1   g734(.A1(new_n925), .A2(new_n818), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n315), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n937), .B1(G183gat), .B2(new_n936), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n938), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g738(.A1(new_n927), .A2(new_n317), .A3(new_n717), .ZN(new_n940));
  OAI21_X1  g739(.A(G190gat), .B1(new_n925), .B2(new_n619), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT125), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n942), .A2(KEYINPUT61), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(KEYINPUT61), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(G1351gat));
  NAND2_X1  g744(.A1(new_n690), .A2(new_n472), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n742), .A2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n886), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(G197gat), .B1(new_n949), .B2(new_n581), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n948), .B1(new_n902), .B2(new_n909), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n581), .A2(G197gat), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(G1352gat));
  INV_X1    g752(.A(new_n951), .ZN(new_n954));
  OAI21_X1  g753(.A(G204gat), .B1(new_n954), .B2(new_n670), .ZN(new_n955));
  NOR4_X1   g754(.A1(new_n886), .A2(G204gat), .A3(new_n670), .A4(new_n948), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT62), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(G1353gat));
  AOI21_X1  g757(.A(KEYINPUT57), .B1(new_n906), .B2(new_n907), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n642), .B(new_n947), .C1(new_n959), .C2(new_n901), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n960), .A2(KEYINPUT127), .ZN(new_n961));
  OAI21_X1  g760(.A(G211gat), .B1(new_n960), .B2(KEYINPUT127), .ZN(new_n962));
  OAI21_X1  g761(.A(KEYINPUT63), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n951), .A2(new_n964), .A3(new_n642), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT63), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n960), .A2(KEYINPUT127), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n965), .A2(new_n966), .A3(G211gat), .A4(new_n967), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n949), .A2(new_n399), .A3(new_n642), .ZN(new_n969));
  XOR2_X1   g768(.A(new_n969), .B(KEYINPUT126), .Z(new_n970));
  NAND3_X1  g769(.A1(new_n963), .A2(new_n968), .A3(new_n970), .ZN(G1354gat));
  OAI21_X1  g770(.A(G218gat), .B1(new_n954), .B2(new_n619), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n949), .A2(new_n400), .A3(new_n717), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(G1355gat));
endmodule


