//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G57gat), .B(G85gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT5), .ZN(new_n208));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT2), .ZN(new_n210));
  INV_X1    g009(.A(G141gat), .ZN(new_n211));
  INV_X1    g010(.A(G148gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  AND3_X1   g014(.A1(KEYINPUT75), .A2(G155gat), .A3(G162gat), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT76), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(G155gat), .B2(G162gat), .ZN(new_n220));
  INV_X1    g019(.A(G155gat), .ZN(new_n221));
  INV_X1    g020(.A(G162gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT76), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n215), .A2(new_n218), .A3(new_n220), .A4(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT2), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n221), .B(new_n222), .C1(new_n225), .C2(KEYINPUT77), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(new_n209), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n213), .A2(new_n214), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n210), .A2(KEYINPUT77), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G134gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G127gat), .ZN(new_n233));
  INV_X1    g032(.A(G127gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G134gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G113gat), .B(G120gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n236), .B1(new_n237), .B2(KEYINPUT1), .ZN(new_n238));
  INV_X1    g037(.A(G120gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G113gat), .ZN(new_n240));
  INV_X1    g039(.A(G113gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G120gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G127gat), .B(G134gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT1), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n238), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT78), .B1(new_n231), .B2(new_n247), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n238), .A2(new_n246), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT78), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n249), .A2(new_n250), .A3(new_n230), .A4(new_n224), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n231), .A2(new_n247), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n248), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G225gat), .A2(G233gat), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n208), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n248), .A2(new_n251), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n231), .A2(KEYINPUT3), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT3), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n224), .A2(new_n230), .A3(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n247), .A3(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n231), .A2(new_n247), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT4), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n258), .A2(new_n254), .A3(new_n262), .A4(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n256), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT79), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT79), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n256), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n248), .A2(new_n251), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT4), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT81), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n263), .A2(KEYINPUT4), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n257), .B1(new_n248), .B2(new_n251), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT81), .B1(new_n277), .B2(new_n274), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n262), .A2(new_n208), .A3(new_n254), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n207), .B1(new_n270), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT6), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n256), .A2(new_n265), .A3(new_n268), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n268), .B1(new_n256), .B2(new_n265), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n280), .A2(new_n207), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n283), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT82), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n288), .A2(new_n281), .A3(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n280), .A2(new_n207), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT6), .B1(new_n291), .B2(new_n270), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n280), .B1(new_n284), .B2(new_n285), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(new_n206), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT82), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n282), .B1(new_n290), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT83), .ZN(new_n297));
  XOR2_X1   g096(.A(G197gat), .B(G204gat), .Z(new_n298));
  AND2_X1   g097(.A1(G211gat), .A2(G218gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(G211gat), .A2(G218gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n299), .A2(KEYINPUT22), .ZN(new_n302));
  OR3_X1    g101(.A1(new_n298), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(new_n298), .B2(new_n302), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G226gat), .A2(G233gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(KEYINPUT69), .ZN(new_n309));
  NAND2_X1  g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT26), .ZN(new_n312));
  NOR2_X1   g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n309), .A2(new_n314), .B1(G183gat), .B2(G190gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT27), .B(G183gat), .ZN(new_n316));
  INV_X1    g115(.A(G190gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT28), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n316), .A2(KEYINPUT28), .A3(new_n317), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n315), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G183gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n317), .ZN(new_n325));
  NAND3_X1  g124(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n327), .B1(KEYINPUT68), .B2(KEYINPUT24), .ZN(new_n328));
  AND2_X1   g127(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n325), .B(new_n326), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G169gat), .ZN(new_n331));
  INV_X1    g130(.A(G176gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT66), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT66), .B1(new_n313), .B2(KEYINPUT23), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n310), .A2(KEYINPUT25), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n339), .B1(KEYINPUT23), .B2(new_n313), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n330), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  XOR2_X1   g140(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n342));
  AOI21_X1  g141(.A(new_n334), .B1(new_n333), .B2(new_n335), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n313), .A2(KEYINPUT66), .A3(KEYINPUT23), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n310), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT24), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n327), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(new_n325), .A3(new_n326), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n313), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT65), .B1(new_n313), .B2(KEYINPUT23), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n342), .B1(new_n345), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT67), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n341), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI211_X1 g153(.A(KEYINPUT67), .B(new_n342), .C1(new_n345), .C2(new_n351), .ZN(new_n355));
  AOI211_X1 g154(.A(new_n307), .B(new_n323), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n307), .A2(KEYINPUT29), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n352), .A2(new_n353), .ZN(new_n358));
  INV_X1    g157(.A(new_n341), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(new_n355), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n323), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n305), .B1(new_n356), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n360), .A2(new_n361), .A3(new_n306), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n303), .A2(new_n304), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n323), .B1(new_n354), .B2(new_n355), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n364), .B(new_n365), .C1(new_n366), .C2(new_n357), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n363), .A2(KEYINPUT72), .A3(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n356), .A2(new_n362), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT72), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(new_n370), .A3(new_n365), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(G8gat), .B(G36gat), .Z(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(KEYINPUT73), .ZN(new_n374));
  XNOR2_X1  g173(.A(G64gat), .B(G92gat), .ZN(new_n375));
  XOR2_X1   g174(.A(new_n374), .B(new_n375), .Z(new_n376));
  NAND2_X1  g175(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT74), .B(KEYINPUT30), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n372), .A2(KEYINPUT30), .A3(new_n376), .ZN(new_n380));
  INV_X1    g179(.A(new_n376), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n368), .A2(new_n371), .A3(new_n381), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n296), .A2(new_n297), .A3(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n294), .A2(new_n283), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n289), .B1(new_n288), .B2(new_n281), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n292), .A2(KEYINPUT82), .A3(new_n294), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT83), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n305), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n304), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n299), .A2(new_n300), .A3(new_n392), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT29), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT3), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n224), .A2(new_n230), .ZN(new_n398));
  INV_X1    g197(.A(G228gat), .ZN(new_n399));
  INV_X1    g198(.A(G233gat), .ZN(new_n400));
  OAI22_X1  g199(.A1(new_n397), .A2(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT29), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n365), .B1(new_n402), .B2(new_n261), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT86), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n404), .A2(KEYINPUT86), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n401), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n260), .B1(new_n305), .B2(KEYINPUT29), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n231), .ZN(new_n410));
  AOI211_X1 g209(.A(new_n399), .B(new_n400), .C1(new_n410), .C2(new_n404), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n391), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n393), .A2(new_n396), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n260), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n414), .A2(new_n231), .B1(G228gat), .B2(G233gat), .ZN(new_n415));
  INV_X1    g214(.A(new_n407), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(new_n416), .A3(new_n405), .ZN(new_n417));
  INV_X1    g216(.A(new_n411), .ZN(new_n418));
  INV_X1    g217(.A(new_n391), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G78gat), .B(G106gat), .ZN(new_n421));
  INV_X1    g220(.A(G50gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(G22gat), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n412), .A2(new_n420), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n424), .B1(new_n412), .B2(new_n420), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(G227gat), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(new_n400), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n366), .A2(new_n249), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n366), .A2(new_n249), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT32), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT33), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(G71gat), .B(G99gat), .Z(new_n436));
  XNOR2_X1  g235(.A(G15gat), .B(G43gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n433), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT70), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n434), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n441), .B1(new_n440), .B2(new_n438), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n432), .A2(KEYINPUT32), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  OR2_X1    g243(.A1(new_n366), .A2(new_n249), .ZN(new_n445));
  INV_X1    g244(.A(new_n429), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n366), .A2(new_n249), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT34), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT34), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n445), .A2(new_n450), .A3(new_n446), .A4(new_n447), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT71), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n444), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n439), .A2(new_n452), .A3(KEYINPUT71), .A4(new_n443), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n427), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n384), .A2(new_n390), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT35), .ZN(new_n458));
  XNOR2_X1  g257(.A(KEYINPUT87), .B(KEYINPUT35), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n292), .A2(new_n294), .ZN(new_n460));
  AOI211_X1 g259(.A(new_n459), .B(new_n427), .C1(new_n282), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n452), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n449), .A2(new_n451), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(new_n439), .A3(new_n443), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n465), .A2(new_n389), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n458), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n384), .A2(new_n390), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n427), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT36), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n471), .B1(new_n454), .B2(new_n455), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT36), .B1(new_n462), .B2(new_n464), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n381), .A2(KEYINPUT37), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n382), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n363), .A2(new_n367), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT38), .B1(new_n477), .B2(KEYINPUT37), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n479), .A2(new_n282), .A3(new_n460), .A4(new_n377), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT38), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n368), .A2(KEYINPUT37), .A3(new_n371), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n482), .B1(new_n476), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n427), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n276), .A2(new_n278), .A3(new_n262), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(new_n255), .ZN(new_n488));
  OR2_X1    g287(.A1(new_n253), .A2(new_n255), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(KEYINPUT39), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT39), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n487), .A2(new_n491), .A3(new_n255), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n207), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT40), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n490), .A2(KEYINPUT40), .A3(new_n207), .A4(new_n492), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(new_n294), .A3(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n383), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n474), .B1(new_n486), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n470), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n468), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(G29gat), .A2(G36gat), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT14), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(G29gat), .A2(G36gat), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(G43gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(G50gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n422), .A2(G43gat), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT15), .ZN(new_n511));
  INV_X1    g310(.A(G29gat), .ZN(new_n512));
  INV_X1    g311(.A(G36gat), .ZN(new_n513));
  OR3_X1    g312(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT90), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT90), .B1(new_n512), .B2(new_n513), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n505), .A2(new_n511), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n422), .A2(G43gat), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT89), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n517), .B1(new_n518), .B2(new_n510), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n422), .A2(KEYINPUT89), .A3(G43gat), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT15), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI22_X1  g320(.A1(new_n507), .A2(new_n511), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n522), .B(KEYINPUT17), .Z(new_n523));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n524), .A2(G1gat), .ZN(new_n525));
  INV_X1    g324(.A(G8gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT16), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n524), .B1(new_n527), .B2(G1gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT92), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT91), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n525), .A2(new_n531), .A3(new_n528), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n532), .B(G8gat), .C1(new_n531), .C2(new_n528), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  OR3_X1    g333(.A1(new_n523), .A2(KEYINPUT93), .A3(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n523), .A2(new_n534), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n522), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT93), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n535), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT18), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n534), .B(new_n522), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n540), .B(KEYINPUT13), .Z(new_n544));
  AOI22_X1  g343(.A1(new_n541), .A2(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n536), .A2(new_n538), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n546), .A2(new_n535), .B1(G229gat), .B2(G233gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT18), .ZN(new_n548));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(G169gat), .B(G197gat), .Z(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT12), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n545), .A2(new_n548), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n554), .B1(new_n545), .B2(new_n548), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT94), .B1(new_n502), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n457), .A2(KEYINPUT35), .B1(new_n466), .B2(new_n461), .ZN(new_n560));
  INV_X1    g359(.A(new_n427), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n561), .B1(new_n384), .B2(new_n390), .ZN(new_n562));
  INV_X1    g361(.A(new_n455), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n439), .A2(new_n443), .B1(new_n452), .B2(KEYINPUT71), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT36), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n463), .A2(new_n439), .A3(new_n443), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n463), .B1(new_n443), .B2(new_n439), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n471), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n561), .B1(new_n480), .B2(new_n484), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n569), .B1(new_n570), .B2(new_n498), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n562), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g371(.A(KEYINPUT94), .B(new_n558), .C1(new_n560), .C2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n559), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(new_n296), .ZN(new_n576));
  NAND2_X1  g375(.A1(G85gat), .A2(G92gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT7), .ZN(new_n578));
  NAND2_X1  g377(.A1(G99gat), .A2(G106gat), .ZN(new_n579));
  INV_X1    g378(.A(G85gat), .ZN(new_n580));
  INV_X1    g379(.A(G92gat), .ZN(new_n581));
  AOI22_X1  g380(.A1(KEYINPUT8), .A2(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G99gat), .B(G106gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n523), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n522), .A2(new_n585), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT41), .ZN(new_n588));
  NAND2_X1  g387(.A1(G232gat), .A2(G233gat), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(G190gat), .B(G218gat), .Z(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n589), .A2(new_n588), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT95), .ZN(new_n595));
  XOR2_X1   g394(.A(G134gat), .B(G162gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n593), .A2(new_n597), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G57gat), .B(G64gat), .Z(new_n602));
  INV_X1    g401(.A(KEYINPUT9), .ZN(new_n603));
  INV_X1    g402(.A(G71gat), .ZN(new_n604));
  INV_X1    g403(.A(G78gat), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G71gat), .B(G78gat), .Z(new_n608));
  OR2_X1    g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT21), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G127gat), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n530), .B(new_n533), .C1(new_n612), .C2(new_n611), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(new_n221), .ZN(new_n622));
  XNOR2_X1  g421(.A(G183gat), .B(G211gat), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n622), .B(new_n623), .Z(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n618), .A2(new_n619), .A3(new_n624), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G120gat), .B(G148gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(G176gat), .B(G204gat), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n629), .B(new_n630), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n585), .B(new_n611), .ZN(new_n632));
  NAND2_X1  g431(.A1(G230gat), .A2(G233gat), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT96), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n631), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n637), .B1(new_n636), .B2(new_n635), .ZN(new_n638));
  INV_X1    g437(.A(new_n633), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT10), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n632), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n585), .A2(KEYINPUT10), .A3(new_n610), .A4(new_n609), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n638), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n631), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n643), .B2(new_n634), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n601), .A2(new_n628), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n576), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(G1gat), .ZN(G1324gat));
  NOR3_X1   g452(.A1(new_n575), .A2(new_n650), .A3(new_n383), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT16), .B(G8gat), .Z(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(new_n526), .B2(new_n654), .ZN(new_n657));
  MUX2_X1   g456(.A(new_n656), .B(new_n657), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g457(.A(KEYINPUT94), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n560), .A2(new_n572), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n659), .B1(new_n660), .B2(new_n557), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n573), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n651), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n465), .ZN(new_n665));
  AOI21_X1  g464(.A(G15gat), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n474), .A2(G15gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n667), .B(KEYINPUT97), .Z(new_n668));
  AOI21_X1  g467(.A(new_n666), .B1(new_n664), .B2(new_n668), .ZN(G1326gat));
  NOR2_X1   g468(.A1(new_n663), .A2(new_n561), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT43), .B(G22gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1327gat));
  NOR3_X1   g471(.A1(new_n601), .A2(new_n628), .A3(new_n648), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n576), .A2(new_n512), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT45), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n648), .B(KEYINPUT98), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n678), .A2(new_n557), .A3(new_n628), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(KEYINPUT99), .A2(KEYINPUT44), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(KEYINPUT99), .A2(KEYINPUT44), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(new_n660), .B2(new_n601), .ZN(new_n686));
  INV_X1    g485(.A(new_n601), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n687), .B(new_n681), .C1(new_n560), .C2(new_n572), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n680), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(G29gat), .B1(new_n690), .B2(new_n296), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n675), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n676), .A2(new_n691), .A3(new_n692), .ZN(G1328gat));
  OAI21_X1  g492(.A(G36gat), .B1(new_n690), .B2(new_n383), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n575), .A2(new_n383), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n695), .A2(new_n513), .A3(new_n673), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT100), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT100), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n695), .A2(new_n699), .A3(new_n513), .A4(new_n673), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n698), .B1(new_n697), .B2(new_n700), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n694), .B1(new_n701), .B2(new_n702), .ZN(G1329gat));
  OAI21_X1  g502(.A(G43gat), .B1(new_n690), .B2(new_n569), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n673), .A2(new_n508), .A3(new_n665), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n575), .B2(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g506(.A(new_n422), .B1(new_n689), .B2(new_n427), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n427), .A2(new_n422), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n673), .B1(KEYINPUT102), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n710), .B1(KEYINPUT102), .B2(new_n709), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(new_n559), .B2(new_n574), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT48), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT103), .B1(new_n708), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n684), .B1(new_n502), .B2(new_n687), .ZN(new_n715));
  INV_X1    g514(.A(new_n688), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n427), .B(new_n679), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G50gat), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n718), .A2(new_n719), .A3(KEYINPUT48), .A4(new_n712), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n714), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n712), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n722), .B1(new_n718), .B2(KEYINPUT101), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT101), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT48), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT104), .B1(new_n721), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT48), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n712), .B1(new_n708), .B2(new_n724), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n718), .A2(KEYINPUT101), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n714), .A2(new_n720), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n727), .A2(new_n734), .ZN(G1331gat));
  INV_X1    g534(.A(new_n628), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n687), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n502), .A2(new_n737), .A3(new_n557), .A4(new_n678), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n388), .ZN(new_n740));
  XNOR2_X1  g539(.A(KEYINPUT105), .B(G57gat), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1332gat));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n389), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n744));
  XOR2_X1   g543(.A(KEYINPUT49), .B(G64gat), .Z(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n743), .B2(new_n745), .ZN(G1333gat));
  OAI21_X1  g545(.A(G71gat), .B1(new_n738), .B2(new_n569), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n665), .A2(new_n604), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n738), .B2(new_n748), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g549(.A1(new_n739), .A2(new_n427), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT107), .ZN(new_n752));
  XOR2_X1   g551(.A(KEYINPUT106), .B(G78gat), .Z(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1335gat));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n660), .A2(new_n601), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n756), .A2(KEYINPUT108), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n558), .A2(new_n628), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(KEYINPUT108), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n757), .A2(KEYINPUT51), .A3(new_n758), .A4(new_n759), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n755), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n762), .A2(KEYINPUT109), .A3(new_n764), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n296), .A2(G85gat), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n766), .A2(new_n648), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n686), .A2(new_n688), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n558), .A2(new_n628), .A3(new_n649), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(G85gat), .B1(new_n772), .B2(new_n296), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n769), .A2(new_n773), .ZN(G1336gat));
  NOR3_X1   g573(.A1(new_n677), .A2(G92gat), .A3(new_n383), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(new_n763), .B2(new_n765), .ZN(new_n776));
  INV_X1    g575(.A(new_n772), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n581), .B1(new_n777), .B2(new_n389), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(KEYINPUT52), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n775), .B(KEYINPUT110), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n762), .B2(new_n764), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT52), .B1(new_n782), .B2(new_n778), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n783), .ZN(G1337gat));
  NOR2_X1   g583(.A1(new_n465), .A2(G99gat), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n766), .A2(new_n648), .A3(new_n767), .A4(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G99gat), .B1(new_n772), .B2(new_n569), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(G1338gat));
  INV_X1    g587(.A(G106gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n678), .A2(new_n789), .A3(new_n427), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n762), .B2(new_n764), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n789), .B1(new_n777), .B2(new_n427), .ZN(new_n792));
  OR3_X1    g591(.A1(new_n791), .A2(KEYINPUT53), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(KEYINPUT53), .B1(new_n791), .B2(new_n792), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(G1339gat));
  NOR3_X1   g594(.A1(new_n650), .A2(new_n556), .A3(new_n555), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n543), .A2(new_n544), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n797), .A2(KEYINPUT112), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(KEYINPUT112), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n798), .B(new_n799), .C1(new_n540), .C2(new_n539), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n553), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n545), .A2(new_n548), .A3(new_n554), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n802), .A3(new_n648), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n641), .A2(new_n639), .A3(new_n642), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(KEYINPUT111), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n805), .A2(KEYINPUT54), .A3(new_n644), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n631), .B1(new_n643), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  AOI22_X1  g609(.A1(new_n809), .A2(new_n810), .B1(new_n644), .B2(new_n638), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n806), .A2(KEYINPUT55), .A3(new_n808), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n601), .B(new_n803), .C1(new_n557), .C2(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n811), .A2(new_n802), .A3(new_n812), .A4(new_n801), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n628), .B1(new_n815), .B2(new_n687), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n796), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n817), .A2(new_n296), .A3(new_n427), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n466), .ZN(new_n819));
  OAI21_X1  g618(.A(G113gat), .B1(new_n819), .B2(new_n557), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n818), .B(new_n383), .C1(new_n564), .C2(new_n563), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n557), .A2(G113gat), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT113), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n820), .B1(new_n821), .B2(new_n823), .ZN(G1340gat));
  NOR3_X1   g623(.A1(new_n819), .A2(new_n239), .A3(new_n677), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n821), .A2(new_n649), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n825), .B1(new_n826), .B2(new_n239), .ZN(G1341gat));
  NOR3_X1   g626(.A1(new_n819), .A2(new_n234), .A3(new_n736), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n821), .A2(new_n736), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n829), .A2(KEYINPUT114), .ZN(new_n830));
  AOI21_X1  g629(.A(G127gat), .B1(new_n829), .B2(KEYINPUT114), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(G1342gat));
  NOR3_X1   g631(.A1(new_n821), .A2(G134gat), .A3(new_n601), .ZN(new_n833));
  XOR2_X1   g632(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n834));
  OR2_X1    g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(G134gat), .B1(new_n819), .B2(new_n601), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n833), .A2(new_n834), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(G1343gat));
  NOR3_X1   g637(.A1(new_n474), .A2(new_n296), .A3(new_n389), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n814), .A2(new_n816), .ZN(new_n840));
  INV_X1    g639(.A(new_n796), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT57), .B1(new_n842), .B2(new_n427), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n817), .A2(new_n844), .A3(new_n561), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n839), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(G141gat), .B1(new_n846), .B2(new_n557), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n842), .A2(new_n427), .A3(new_n839), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(new_n211), .A3(new_n558), .ZN(new_n849));
  XNOR2_X1  g648(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n849), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n846), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g653(.A(KEYINPUT116), .B(new_n839), .C1(new_n843), .C2(new_n845), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(new_n558), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n852), .B1(new_n856), .B2(G141gat), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT58), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n851), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g660(.A(KEYINPUT118), .B(new_n851), .C1(new_n857), .C2(new_n858), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1344gat));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n212), .A3(new_n648), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865));
  OR3_X1    g664(.A1(new_n843), .A2(new_n845), .A3(KEYINPUT119), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n843), .A2(KEYINPUT119), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n648), .A3(new_n839), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n865), .B1(new_n869), .B2(G148gat), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n871));
  AOI211_X1 g670(.A(KEYINPUT59), .B(new_n212), .C1(new_n871), .C2(new_n648), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n864), .B1(new_n870), .B2(new_n872), .ZN(G1345gat));
  NAND3_X1  g672(.A1(new_n848), .A2(new_n221), .A3(new_n628), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n871), .A2(new_n628), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n875), .B2(new_n221), .ZN(G1346gat));
  NAND3_X1  g675(.A1(new_n848), .A2(new_n222), .A3(new_n687), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n871), .A2(new_n687), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n222), .ZN(G1347gat));
  NOR2_X1   g678(.A1(new_n817), .A2(new_n427), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n296), .A2(new_n389), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(new_n465), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n331), .B1(new_n883), .B2(new_n558), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(KEYINPUT121), .ZN(new_n885));
  INV_X1    g684(.A(new_n456), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n817), .A2(new_n886), .A3(new_n881), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT120), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n331), .A3(new_n558), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n885), .A2(new_n889), .ZN(G1348gat));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n332), .A3(new_n648), .ZN(new_n891));
  INV_X1    g690(.A(new_n883), .ZN(new_n892));
  OAI21_X1  g691(.A(G176gat), .B1(new_n892), .B2(new_n677), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(G1349gat));
  AOI21_X1  g693(.A(new_n324), .B1(new_n883), .B2(new_n628), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n887), .A2(new_n628), .A3(new_n316), .ZN(new_n896));
  OAI22_X1  g695(.A1(new_n895), .A2(new_n896), .B1(KEYINPUT122), .B2(KEYINPUT60), .ZN(new_n897));
  NAND2_X1  g696(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT123), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n897), .B(new_n899), .ZN(G1350gat));
  NAND3_X1  g699(.A1(new_n888), .A2(new_n317), .A3(new_n687), .ZN(new_n901));
  OAI21_X1  g700(.A(G190gat), .B1(new_n892), .B2(new_n601), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n902), .A2(KEYINPUT124), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(KEYINPUT124), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n904), .B1(new_n903), .B2(new_n905), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n901), .B1(new_n906), .B2(new_n907), .ZN(G1351gat));
  NOR2_X1   g707(.A1(new_n474), .A2(new_n881), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n868), .A2(G197gat), .A3(new_n558), .A4(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(G197gat), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n842), .A2(new_n427), .A3(new_n909), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n912), .B2(new_n557), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n910), .A2(new_n913), .ZN(G1352gat));
  NOR3_X1   g713(.A1(new_n912), .A2(G204gat), .A3(new_n649), .ZN(new_n915));
  NAND2_X1  g714(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n916));
  OR2_X1    g715(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n918), .B1(new_n916), .B2(new_n915), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n866), .A2(new_n867), .A3(new_n678), .A4(new_n909), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(G204gat), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT126), .ZN(G1353gat));
  OR3_X1    g722(.A1(new_n912), .A2(G211gat), .A3(new_n736), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n868), .A2(new_n628), .A3(new_n909), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n925), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT63), .B1(new_n925), .B2(G211gat), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(G1354gat));
  NOR3_X1   g727(.A1(new_n912), .A2(G218gat), .A3(new_n601), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n866), .A2(new_n867), .A3(new_n687), .A4(new_n909), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n930), .B2(G218gat), .ZN(new_n931));
  XOR2_X1   g730(.A(new_n931), .B(KEYINPUT127), .Z(G1355gat));
endmodule


