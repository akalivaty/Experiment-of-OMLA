//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1301, new_n1302, new_n1303,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT64), .Z(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT65), .B(G244), .ZN(new_n218));
  AND2_X1   g0018(.A1(new_n218), .A2(G77), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  XOR2_X1   g0043(.A(KEYINPUT8), .B(G58), .Z(new_n244));
  NAND2_X1  g0044(.A1(new_n206), .A2(G20), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n215), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G13), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(G1), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G20), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  OAI22_X1  g0053(.A1(new_n246), .A2(new_n253), .B1(new_n252), .B2(new_n244), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT67), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(new_n207), .A3(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(KEYINPUT67), .B1(G20), .B2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G159), .ZN(new_n260));
  INV_X1    g0060(.A(G58), .ZN(new_n261));
  INV_X1    g0061(.A(G68), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(G20), .B1(new_n263), .B2(new_n201), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(new_n268), .A3(KEYINPUT74), .ZN(new_n269));
  OR3_X1    g0069(.A1(new_n256), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(new_n270), .A3(new_n207), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n262), .B1(new_n271), .B2(KEYINPUT7), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n269), .A2(new_n270), .A3(new_n207), .A4(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n265), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n249), .B1(new_n275), .B2(KEYINPUT16), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT16), .ZN(new_n277));
  INV_X1    g0077(.A(new_n265), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n273), .B1(new_n279), .B2(G20), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n267), .A2(new_n268), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n262), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT76), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n278), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI211_X1 g0085(.A(KEYINPUT76), .B(new_n262), .C1(new_n280), .C2(new_n282), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n277), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n254), .B1(new_n276), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G169), .ZN(new_n289));
  AND2_X1   g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(new_n215), .ZN(new_n291));
  INV_X1    g0091(.A(G226), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G1698), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(G223), .B2(G1698), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(new_n270), .B2(new_n269), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G87), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n291), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT66), .ZN(new_n299));
  OAI21_X1  g0099(.A(G274), .B1(new_n290), .B2(new_n215), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G274), .ZN(new_n303));
  AND2_X1   g0103(.A1(G1), .A2(G13), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G41), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G41), .ZN(new_n307));
  INV_X1    g0107(.A(G45), .ZN(new_n308));
  AOI21_X1  g0108(.A(G1), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(KEYINPUT66), .A3(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n291), .A2(new_n309), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n302), .A2(new_n310), .B1(new_n311), .B2(G232), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n289), .B1(new_n298), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n304), .A2(new_n305), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n269), .A2(new_n270), .ZN(new_n315));
  INV_X1    g0115(.A(new_n294), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n314), .B1(new_n317), .B2(new_n296), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n311), .A2(G232), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n300), .A2(new_n299), .A3(new_n301), .ZN(new_n320));
  AOI21_X1  g0120(.A(KEYINPUT66), .B1(new_n306), .B2(new_n309), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n313), .B1(new_n323), .B2(G179), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT18), .B1(new_n288), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n254), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT7), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT75), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT75), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT7), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n207), .B2(new_n281), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n279), .A2(new_n327), .A3(G20), .ZN(new_n333));
  OAI21_X1  g0133(.A(G68), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n265), .B1(new_n334), .B2(KEYINPUT76), .ZN(new_n335));
  INV_X1    g0135(.A(new_n286), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT16), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n271), .A2(KEYINPUT7), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n338), .A2(G68), .A3(new_n274), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n339), .A2(KEYINPUT16), .A3(new_n278), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n248), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n326), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT18), .ZN(new_n343));
  INV_X1    g0143(.A(new_n324), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G200), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n318), .B2(new_n322), .ZN(new_n347));
  INV_X1    g0147(.A(G190), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n298), .A2(new_n312), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n350), .B(new_n326), .C1(new_n337), .C2(new_n341), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT77), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n354), .A2(KEYINPUT17), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n355), .B1(new_n288), .B2(new_n350), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n325), .B(new_n345), .C1(new_n353), .C2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G97), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n229), .A2(G1698), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(G226), .B2(G1698), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n359), .B1(new_n361), .B2(new_n281), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n362), .A2(new_n291), .B1(new_n311), .B2(G238), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT13), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n302), .A2(new_n310), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n364), .B1(new_n363), .B2(new_n365), .ZN(new_n368));
  OAI21_X1  g0168(.A(G169), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT14), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n366), .A2(KEYINPUT71), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n366), .A2(KEYINPUT71), .ZN(new_n372));
  INV_X1    g0172(.A(new_n368), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n371), .A2(G179), .A3(new_n372), .A4(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT14), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n375), .B(G169), .C1(new_n367), .C2(new_n368), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n370), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n250), .A2(new_n207), .A3(G1), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(new_n248), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n379), .A2(G68), .A3(new_n245), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT73), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n262), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n382), .B(KEYINPUT12), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n259), .A2(KEYINPUT72), .A3(G50), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT72), .B1(new_n259), .B2(G50), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n256), .A2(G20), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G77), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n389), .A2(new_n390), .B1(new_n207), .B2(G68), .ZN(new_n391));
  OAI211_X1 g0191(.A(KEYINPUT11), .B(new_n248), .C1(new_n387), .C2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT11), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n387), .A2(new_n391), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n393), .B1(new_n394), .B2(new_n249), .ZN(new_n395));
  AND3_X1   g0195(.A1(new_n384), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n377), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n371), .A2(G190), .A3(new_n372), .A4(new_n373), .ZN(new_n399));
  OAI21_X1  g0199(.A(G200), .B1(new_n367), .B2(new_n368), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n396), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n379), .A2(G77), .A3(new_n245), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(G77), .B2(new_n252), .ZN(new_n404));
  XOR2_X1   g0204(.A(KEYINPUT15), .B(G87), .Z(new_n405));
  AOI22_X1  g0205(.A1(new_n405), .A2(new_n388), .B1(G20), .B2(G77), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n244), .A2(new_n259), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n249), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n311), .A2(new_n218), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n365), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT70), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT70), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n365), .A2(new_n413), .A3(new_n410), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n279), .A2(G238), .A3(G1698), .ZN(new_n415));
  INV_X1    g0215(.A(G1698), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n279), .A2(G232), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G107), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n415), .B(new_n417), .C1(new_n418), .C2(new_n279), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n291), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n412), .A2(new_n414), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n409), .B1(new_n421), .B2(new_n289), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n411), .A2(KEYINPUT70), .B1(new_n291), .B2(new_n419), .ZN(new_n423));
  INV_X1    g0223(.A(G179), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(new_n414), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n245), .A2(KEYINPUT68), .A3(G50), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT68), .B1(new_n245), .B2(G50), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n430), .A2(new_n379), .B1(new_n202), .B2(new_n378), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n203), .A2(G20), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT8), .B(G58), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n432), .B1(new_n433), .B2(new_n389), .ZN(new_n434));
  INV_X1    g0234(.A(G150), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(new_n257), .B2(new_n258), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n248), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n431), .A2(KEYINPUT9), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n314), .B1(new_n281), .B2(new_n390), .ZN(new_n439));
  MUX2_X1   g0239(.A(G222), .B(G223), .S(G1698), .Z(new_n440));
  OAI21_X1  g0240(.A(new_n439), .B1(new_n281), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n311), .A2(G226), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n441), .A2(new_n365), .A3(G190), .A4(new_n442), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n431), .A2(new_n437), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT9), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n441), .A2(new_n365), .A3(new_n442), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n445), .A2(new_n446), .B1(new_n447), .B2(G200), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT10), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n444), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n447), .A2(G200), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n244), .A2(new_n388), .B1(G20), .B2(new_n203), .ZN(new_n452));
  INV_X1    g0252(.A(new_n436), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n249), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n378), .A2(new_n202), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n245), .A2(G50), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT68), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n427), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n455), .B1(new_n459), .B2(new_n253), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n446), .B1(new_n454), .B2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n451), .A2(new_n461), .A3(new_n438), .A4(new_n443), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT10), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n450), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n421), .A2(G200), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n412), .A2(G190), .A3(new_n414), .A4(new_n420), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(new_n409), .A3(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n441), .A2(new_n365), .A3(new_n424), .A4(new_n442), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT69), .ZN(new_n469));
  XNOR2_X1  g0269(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n454), .A2(new_n460), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n471), .B1(new_n289), .B2(new_n447), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  AND4_X1   g0273(.A1(new_n426), .A2(new_n464), .A3(new_n467), .A4(new_n473), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n358), .A2(new_n402), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT83), .ZN(new_n477));
  XNOR2_X1  g0277(.A(G97), .B(G107), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT6), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G97), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n479), .A2(new_n481), .A3(G107), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n484), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n485));
  OAI21_X1  g0285(.A(G107), .B1(new_n332), .B2(new_n333), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n249), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OR3_X1    g0287(.A1(new_n252), .A2(KEYINPUT78), .A3(G97), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT78), .B1(new_n252), .B2(G97), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n256), .A2(G1), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n378), .A2(new_n248), .A3(new_n490), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n488), .A2(new_n489), .B1(G97), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n477), .B1(new_n487), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n259), .A2(G77), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n482), .B1(new_n479), .B2(new_n478), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(new_n207), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n418), .B1(new_n280), .B2(new_n282), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n248), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n499), .A2(KEYINPUT83), .A3(new_n492), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT80), .ZN(new_n502));
  INV_X1    g0302(.A(G244), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(G1698), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT4), .B1(new_n315), .B2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n267), .A2(new_n268), .A3(G250), .A4(G1698), .ZN(new_n506));
  AND2_X1   g0306(.A1(KEYINPUT4), .A2(G244), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n267), .A2(new_n268), .A3(new_n507), .A4(new_n416), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G283), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT79), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(KEYINPUT79), .A2(G33), .A3(G283), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n506), .A2(new_n508), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n502), .B1(new_n505), .B2(new_n514), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n506), .A2(new_n508), .A3(new_n513), .ZN(new_n516));
  INV_X1    g0316(.A(new_n504), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n517), .B1(new_n269), .B2(new_n270), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n516), .B(KEYINPUT80), .C1(KEYINPUT4), .C2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n515), .A2(new_n519), .A3(new_n291), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT81), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n307), .A2(KEYINPUT5), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n206), .A2(G45), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n308), .A2(G1), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT5), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G41), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(KEYINPUT81), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n307), .A2(KEYINPUT5), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n524), .A2(new_n528), .A3(new_n306), .A4(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n524), .A2(new_n528), .A3(new_n529), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n314), .ZN(new_n532));
  INV_X1    g0332(.A(G257), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n520), .A2(G179), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n289), .B1(new_n520), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n501), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n405), .A2(new_n252), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n491), .A2(new_n405), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT19), .B1(new_n388), .B2(G97), .ZN(new_n542));
  INV_X1    g0342(.A(G87), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(new_n481), .A3(new_n418), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT86), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT86), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n546), .A2(new_n543), .A3(new_n481), .A4(new_n418), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT19), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n359), .B2(new_n207), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n542), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n315), .A2(new_n207), .A3(G68), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n540), .B(new_n541), .C1(new_n553), .C2(new_n249), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT84), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n300), .B2(new_n523), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n306), .A2(KEYINPUT84), .A3(new_n525), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n314), .A2(G250), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n206), .A2(KEYINPUT85), .A3(G45), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT85), .B1(new_n206), .B2(G45), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n556), .A2(new_n557), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(G238), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n416), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n503), .A2(G1698), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n566), .B1(new_n269), .B2(new_n270), .ZN(new_n567));
  INV_X1    g0367(.A(G116), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n256), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n291), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n562), .A2(new_n570), .A3(new_n424), .ZN(new_n571));
  AOI21_X1  g0371(.A(G169), .B1(new_n562), .B2(new_n570), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n562), .A2(new_n570), .A3(G190), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n346), .B1(new_n562), .B2(new_n570), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n249), .B1(new_n551), .B2(new_n552), .ZN(new_n577));
  INV_X1    g0377(.A(new_n491), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n578), .A2(new_n543), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n577), .A2(new_n539), .A3(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n554), .A2(new_n573), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n487), .A2(new_n493), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n520), .A2(G190), .A3(new_n535), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n346), .B1(new_n520), .B2(new_n535), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n582), .B(new_n583), .C1(new_n584), .C2(KEYINPUT82), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n584), .A2(KEYINPUT82), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n538), .B(new_n581), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT23), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n588), .A2(new_n418), .A3(G20), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT88), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n589), .A2(new_n590), .B1(new_n591), .B2(G20), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT22), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n207), .A2(G87), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n594), .B1(new_n281), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n589), .A2(new_n590), .B1(KEYINPUT23), .B2(G107), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n593), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(KEYINPUT22), .A2(G87), .ZN(new_n599));
  AOI211_X1 g0399(.A(G20), .B(new_n599), .C1(new_n269), .C2(new_n270), .ZN(new_n600));
  OAI21_X1  g0400(.A(KEYINPUT24), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n315), .A2(KEYINPUT22), .A3(new_n207), .A4(G87), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT24), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n604));
  OAI22_X1  g0404(.A1(new_n604), .A2(KEYINPUT88), .B1(new_n588), .B2(new_n418), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n605), .A2(new_n592), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n602), .A2(new_n603), .A3(new_n596), .A4(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n249), .B1(new_n601), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT25), .B1(new_n378), .B2(new_n418), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n378), .A2(KEYINPUT25), .A3(new_n418), .ZN(new_n610));
  OAI22_X1  g0410(.A1(new_n578), .A2(new_n418), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n533), .A2(G1698), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(G250), .B2(G1698), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n270), .B2(new_n269), .ZN(new_n615));
  INV_X1    g0415(.A(G294), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n256), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n291), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n531), .A2(G264), .A3(new_n314), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(new_n530), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n346), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(G190), .B2(new_n620), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n612), .A2(new_n622), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n620), .A2(G179), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n620), .A2(new_n289), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n624), .B(new_n625), .C1(new_n608), .C2(new_n611), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n533), .A2(new_n416), .ZN(new_n628));
  INV_X1    g0428(.A(G264), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(G1698), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n269), .B2(new_n270), .ZN(new_n632));
  OR2_X1    g0432(.A1(KEYINPUT87), .A2(G303), .ZN(new_n633));
  NAND2_X1  g0433(.A1(KEYINPUT87), .A2(G303), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n279), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n291), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n531), .A2(G270), .A3(new_n314), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(new_n637), .A3(new_n530), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G200), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n378), .A2(new_n568), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n491), .A2(G116), .ZN(new_n641));
  AOI21_X1  g0441(.A(G20), .B1(new_n256), .B2(G97), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n513), .A2(new_n642), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n247), .A2(new_n215), .B1(G20), .B2(new_n568), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n643), .A2(new_n644), .A3(KEYINPUT20), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT20), .B1(new_n643), .B2(new_n644), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n640), .B(new_n641), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n639), .B(new_n648), .C1(new_n348), .C2(new_n638), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n647), .A2(new_n638), .A3(G169), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT21), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n647), .A2(new_n638), .A3(KEYINPUT21), .A4(G169), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n636), .A2(new_n637), .A3(G179), .A4(new_n530), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n647), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n649), .A2(new_n652), .A3(new_n653), .A4(new_n656), .ZN(new_n657));
  NOR4_X1   g0457(.A1(new_n476), .A2(new_n587), .A3(new_n627), .A4(new_n657), .ZN(G372));
  NAND2_X1  g0458(.A1(new_n325), .A2(new_n345), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n396), .A2(new_n399), .A3(new_n400), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n398), .B1(new_n660), .B2(new_n426), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n351), .B1(new_n354), .B2(KEYINPUT17), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n351), .B2(new_n352), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n659), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n464), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n473), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n626), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n652), .A2(new_n653), .A3(new_n656), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n623), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n587), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n576), .A2(new_n580), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n573), .A2(new_n554), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT26), .B1(new_n538), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n520), .A2(G179), .A3(new_n535), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n508), .A2(new_n513), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n677), .B(new_n506), .C1(new_n518), .C2(KEYINPUT4), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n314), .B1(new_n678), .B2(new_n502), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n534), .B1(new_n679), .B2(new_n519), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n676), .B1(new_n680), .B2(new_n289), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT26), .ZN(new_n682));
  INV_X1    g0482(.A(new_n582), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n581), .A2(new_n681), .A3(new_n682), .A4(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n675), .A2(new_n673), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n475), .B1(new_n671), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n667), .A2(new_n686), .ZN(G369));
  NAND2_X1  g0487(.A1(new_n251), .A2(new_n207), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(new_n690), .A3(G213), .ZN(new_n691));
  INV_X1    g0491(.A(G343), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n612), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT89), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n696), .A2(new_n626), .A3(new_n623), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n695), .A2(KEYINPUT89), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n669), .A2(new_n694), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n699), .A2(new_n701), .B1(new_n668), .B2(new_n694), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n648), .A2(new_n694), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n669), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n657), .B2(new_n703), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G330), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n697), .A2(new_n698), .B1(new_n626), .B2(new_n694), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n702), .A2(new_n709), .ZN(G399));
  NOR2_X1   g0510(.A1(new_n548), .A2(G116), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n210), .A2(new_n307), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G1), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n214), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n694), .B1(new_n671), .B2(new_n685), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT90), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT29), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT90), .B(new_n694), .C1(new_n671), .C2(new_n685), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT91), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n719), .A2(KEYINPUT91), .A3(new_n720), .A4(new_n721), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n520), .A2(new_n535), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G169), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n582), .B1(new_n727), .B2(new_n676), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n728), .A2(KEYINPUT92), .A3(KEYINPUT26), .A4(new_n581), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n581), .A2(new_n681), .A3(KEYINPUT26), .A4(new_n683), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT92), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n727), .A2(new_n676), .B1(new_n494), .B2(new_n500), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT26), .B1(new_n733), .B2(new_n581), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n673), .B(new_n729), .C1(new_n732), .C2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT93), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n671), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n729), .A2(new_n673), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n738), .B(KEYINPUT93), .C1(new_n734), .C2(new_n732), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n693), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n724), .A2(new_n725), .B1(KEYINPUT29), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT30), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n618), .A2(new_n619), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n562), .A2(new_n570), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n655), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n742), .B1(new_n746), .B2(new_n726), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n654), .A2(new_n743), .A3(new_n744), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n680), .A2(new_n748), .A3(KEYINPUT30), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n620), .A2(new_n424), .A3(new_n744), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n726), .A2(new_n750), .A3(new_n638), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n747), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n693), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT31), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n752), .A2(KEYINPUT31), .A3(new_n693), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n657), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n758), .A2(new_n626), .A3(new_n623), .A4(new_n694), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n587), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n741), .B1(G330), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n716), .B1(new_n763), .B2(G1), .ZN(G364));
  INV_X1    g0564(.A(new_n712), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n250), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n206), .B1(new_n766), .B2(G45), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n707), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(G330), .B2(new_n705), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n210), .A2(new_n279), .ZN(new_n772));
  INV_X1    g0572(.A(G355), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n772), .A2(new_n773), .B1(G116), .B2(new_n210), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n239), .A2(new_n308), .ZN(new_n775));
  INV_X1    g0575(.A(new_n315), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n210), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(new_n308), .B2(new_n214), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n774), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n304), .B1(new_n207), .B2(G169), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n780), .A2(KEYINPUT94), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(KEYINPUT94), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G13), .A2(G33), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n769), .B1(new_n779), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n346), .A2(G179), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n207), .A2(G190), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G179), .A2(G200), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G283), .A2(new_n793), .B1(new_n796), .B2(G329), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT97), .Z(new_n798));
  NAND3_X1  g0598(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(G190), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(KEYINPUT33), .B(G317), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT98), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n803), .B2(new_n802), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n799), .A2(new_n348), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(KEYINPUT96), .B(G326), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n207), .B1(new_n794), .B2(G190), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n809), .B1(G294), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n424), .A2(G200), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n791), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n279), .B1(new_n815), .B2(G311), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n207), .A2(new_n348), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n790), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n817), .A2(new_n813), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G303), .A2(new_n819), .B1(new_n821), .B2(G322), .ZN(new_n822));
  AND3_X1   g0622(.A1(new_n812), .A2(new_n816), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n798), .A2(new_n805), .A3(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G58), .A2(new_n821), .B1(new_n815), .B2(G77), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n202), .B2(new_n807), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT95), .Z(new_n827));
  INV_X1    g0627(.A(G159), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n795), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT32), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n279), .B1(new_n818), .B2(new_n543), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(G107), .B2(new_n793), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n810), .A2(new_n481), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(new_n800), .B2(G68), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n830), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n824), .B1(new_n827), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n789), .B1(new_n836), .B2(new_n783), .ZN(new_n837));
  INV_X1    g0637(.A(new_n786), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n837), .B1(new_n705), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n771), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G396));
  OAI21_X1  g0641(.A(new_n693), .B1(new_n408), .B2(new_n404), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n467), .A2(new_n842), .B1(new_n425), .B2(new_n422), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n422), .A2(new_n425), .A3(new_n694), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(KEYINPUT99), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n466), .A2(new_n409), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n346), .B1(new_n423), .B2(new_n414), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n842), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n426), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT99), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n850), .A2(new_n851), .A3(new_n844), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n846), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n853), .B(new_n694), .C1(new_n671), .C2(new_n685), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n719), .A2(new_n721), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n854), .B1(new_n855), .B2(new_n853), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n762), .A2(G330), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n769), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n857), .B2(new_n856), .ZN(new_n859));
  INV_X1    g0659(.A(new_n783), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n785), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n769), .B1(new_n861), .B2(G77), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n279), .B(new_n833), .C1(G294), .C2(new_n821), .ZN(new_n863));
  AOI22_X1  g0663(.A1(G116), .A2(new_n815), .B1(new_n796), .B2(G311), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n792), .A2(new_n543), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(G107), .B2(new_n819), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G283), .A2(new_n800), .B1(new_n806), .B2(G303), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n863), .A2(new_n864), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(G132), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n795), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n792), .A2(new_n262), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n870), .B(new_n871), .C1(G50), .C2(new_n819), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n776), .B1(G58), .B2(new_n811), .ZN(new_n873));
  AOI22_X1  g0673(.A1(G143), .A2(new_n821), .B1(new_n815), .B2(G159), .ZN(new_n874));
  INV_X1    g0674(.A(G137), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n874), .B1(new_n801), .B2(new_n435), .C1(new_n875), .C2(new_n807), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT34), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n872), .B(new_n873), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n868), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n862), .B1(new_n880), .B2(new_n783), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n853), .B2(new_n785), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n859), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(G384));
  OAI211_X1 g0684(.A(new_n214), .B(G77), .C1(new_n261), .C2(new_n262), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n202), .A2(G68), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n206), .B(G13), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT101), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n484), .A2(KEYINPUT35), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n484), .A2(KEYINPUT35), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n889), .A2(G116), .A3(new_n216), .A4(new_n890), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n891), .B(KEYINPUT36), .Z(new_n892));
  INV_X1    g0692(.A(KEYINPUT100), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n888), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n893), .B2(new_n892), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n666), .B1(new_n741), .B2(new_n475), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n288), .A2(new_n691), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n357), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n351), .B1(new_n288), .B2(new_n324), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT37), .B1(new_n899), .B2(new_n897), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n342), .A2(new_n344), .ZN(new_n901));
  INV_X1    g0701(.A(new_n691), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n342), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT37), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n901), .A2(new_n903), .A3(new_n904), .A4(new_n351), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT38), .B1(new_n898), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT102), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n339), .A2(new_n278), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n277), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n254), .B1(new_n276), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n913), .A2(new_n691), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n357), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n351), .B1(new_n691), .B2(new_n913), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n913), .A2(new_n324), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT37), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n905), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n915), .A2(new_n919), .A3(KEYINPUT38), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n908), .A2(new_n909), .A3(new_n910), .A4(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n398), .A2(new_n693), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n357), .A2(new_n897), .B1(new_n900), .B2(new_n905), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n920), .B(new_n910), .C1(KEYINPUT38), .C2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT102), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n915), .A2(new_n919), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT38), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n910), .B1(new_n928), .B2(new_n920), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n921), .B(new_n922), .C1(new_n925), .C2(new_n929), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n398), .B(new_n401), .C1(new_n396), .C2(new_n694), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n397), .B(new_n693), .C1(new_n660), .C2(new_n377), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(new_n854), .B2(new_n844), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n928), .A2(new_n920), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n935), .A2(new_n936), .B1(new_n659), .B2(new_n691), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n930), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n896), .B(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT103), .B1(new_n757), .B2(new_n760), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n931), .A2(new_n932), .B1(new_n852), .B2(new_n846), .ZN(new_n942));
  INV_X1    g0742(.A(new_n587), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n627), .A2(new_n657), .A3(new_n693), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT103), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n945), .A2(new_n946), .A3(new_n755), .A4(new_n756), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n941), .A2(new_n942), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT40), .B1(new_n928), .B2(new_n920), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n941), .A2(new_n942), .A3(new_n947), .ZN(new_n951));
  AND3_X1   g0751(.A1(new_n915), .A2(new_n919), .A3(KEYINPUT38), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n952), .A2(new_n907), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT40), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n955), .A2(new_n475), .A3(new_n941), .A4(new_n947), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n920), .B1(new_n923), .B2(KEYINPUT38), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n957), .A2(new_n941), .A3(new_n947), .A4(new_n942), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n958), .A2(KEYINPUT40), .B1(new_n948), .B2(new_n949), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n941), .A2(new_n947), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n959), .B1(new_n476), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n956), .A2(new_n961), .A3(G330), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n940), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n206), .B2(new_n766), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n940), .A2(new_n962), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n895), .B1(new_n964), .B2(new_n965), .ZN(G367));
  OAI221_X1 g0766(.A(new_n538), .B1(new_n582), .B2(new_n694), .C1(new_n585), .C2(new_n586), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n728), .A2(new_n693), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n699), .A2(new_n701), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT42), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n538), .B1(new_n970), .B2(new_n626), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n694), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n976), .A2(KEYINPUT104), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(KEYINPUT104), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n580), .A2(new_n694), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n980), .A2(new_n554), .A3(new_n573), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n674), .B2(new_n980), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n709), .A2(new_n970), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n982), .B(KEYINPUT43), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n979), .A2(new_n988), .ZN(new_n989));
  AND3_X1   g0789(.A1(new_n985), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n987), .B1(new_n985), .B2(new_n989), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n724), .A2(new_n725), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n740), .A2(KEYINPUT29), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n857), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n709), .A2(KEYINPUT106), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n702), .A2(KEYINPUT45), .A3(new_n969), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT45), .ZN(new_n999));
  INV_X1    g0799(.A(new_n702), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n999), .B1(new_n1000), .B2(new_n970), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n997), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n702), .A2(new_n969), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT44), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n709), .A2(KEYINPUT106), .ZN(new_n1005));
  AND3_X1   g0805(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1005), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n971), .B1(new_n708), .B2(new_n701), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(new_n706), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n763), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1008), .B1(new_n1012), .B2(KEYINPUT105), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n996), .A2(new_n1010), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT105), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n996), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n712), .B(KEYINPUT41), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n767), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n992), .A2(new_n1019), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n982), .A2(new_n838), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n405), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n787), .B1(new_n210), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n777), .A2(new_n235), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n769), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n818), .A2(new_n568), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n1026), .A2(KEYINPUT46), .B1(new_n616), .B2(new_n801), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(KEYINPUT107), .B(G311), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n807), .A2(new_n1028), .B1(new_n418), .B2(new_n810), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G283), .A2(new_n815), .B1(new_n796), .B2(G317), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n633), .A2(new_n634), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1032), .A2(new_n821), .B1(new_n793), .B2(G97), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n315), .B1(new_n1026), .B2(KEYINPUT46), .ZN(new_n1034));
  AND4_X1   g0834(.A1(new_n1030), .A2(new_n1031), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n793), .A2(G77), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n435), .B2(new_n820), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n279), .B1(new_n818), .B2(new_n261), .C1(new_n828), .C2(new_n801), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n811), .A2(G68), .ZN(new_n1039));
  INV_X1    g0839(.A(G143), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1039), .B1(new_n807), .B2(new_n1040), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n814), .A2(new_n202), .B1(new_n795), .B2(new_n875), .ZN(new_n1042));
  NOR4_X1   g0842(.A1(new_n1037), .A2(new_n1038), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1035), .A2(new_n1043), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1044), .A2(KEYINPUT47), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n860), .B1(new_n1044), .B2(KEYINPUT47), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1025), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1021), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1020), .A2(new_n1048), .ZN(G387));
  NAND2_X1  g0849(.A1(new_n996), .A2(new_n1010), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1012), .A2(new_n765), .A3(new_n1050), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n708), .A2(new_n838), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n711), .A2(new_n772), .B1(G107), .B2(new_n210), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n711), .ZN(new_n1054));
  AOI211_X1 g0854(.A(G45), .B(new_n1054), .C1(G68), .C2(G77), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n433), .A2(G50), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT50), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n777), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1058), .A2(KEYINPUT108), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n232), .A2(new_n308), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n1058), .B2(KEYINPUT108), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1053), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n769), .B1(new_n1062), .B2(new_n788), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n806), .A2(G159), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT109), .Z(new_n1065));
  NAND2_X1  g0865(.A1(new_n819), .A2(G77), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n202), .B2(new_n820), .C1(new_n435), .C2(new_n795), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n315), .B1(new_n262), .B2(new_n814), .C1(new_n481), .C2(new_n792), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n811), .A2(new_n405), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n801), .B2(new_n433), .ZN(new_n1070));
  OR4_X1    g0870(.A1(new_n1065), .A2(new_n1067), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n819), .A2(G294), .B1(new_n811), .B2(G283), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G317), .A2(new_n821), .B1(new_n815), .B2(new_n1032), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n806), .A2(G322), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1073), .B(new_n1074), .C1(new_n801), .C2(new_n1028), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT48), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1072), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT110), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1078), .A2(KEYINPUT49), .A3(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n795), .A2(new_n808), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G116), .B2(new_n793), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(new_n776), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(KEYINPUT49), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1071), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1063), .B1(new_n1085), .B2(new_n783), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1011), .A2(new_n768), .B1(new_n1052), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1051), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(KEYINPUT111), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT111), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1051), .A2(new_n1090), .A3(new_n1087), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1091), .ZN(G393));
  INV_X1    g0892(.A(new_n1008), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n768), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n787), .B1(new_n481), .B2(new_n210), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n777), .A2(new_n242), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n769), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n810), .A2(new_n390), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1098), .B(new_n776), .C1(G50), .C2(new_n800), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n814), .A2(new_n433), .B1(new_n795), .B2(new_n1040), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n865), .B(new_n1100), .C1(G68), .C2(new_n819), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n807), .A2(new_n435), .B1(new_n820), .B2(new_n828), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1102), .B(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1099), .A2(new_n1101), .A3(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G283), .A2(new_n819), .B1(new_n796), .B2(G322), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1106), .B(new_n281), .C1(new_n418), .C2(new_n792), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT113), .Z(new_n1108));
  AOI22_X1  g0908(.A1(new_n821), .A2(G311), .B1(G317), .B2(new_n806), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT52), .Z(new_n1110));
  NAND2_X1  g0910(.A1(new_n1032), .A2(new_n800), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(G294), .A2(new_n815), .B1(new_n811), .B2(G116), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1105), .B1(new_n1108), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1097), .B1(new_n1114), .B2(new_n783), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n969), .B2(new_n838), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1012), .A2(KEYINPUT105), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1117), .A2(new_n1016), .A3(new_n1093), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n765), .B1(new_n1093), .B2(new_n1014), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1094), .B(new_n1116), .C1(new_n1118), .C2(new_n1119), .ZN(G390));
  OAI21_X1  g0920(.A(new_n921), .B1(new_n925), .B2(new_n929), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n854), .A2(new_n844), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n933), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n922), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1123), .A2(KEYINPUT114), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT114), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n935), .B2(new_n922), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1121), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n953), .A2(new_n922), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n845), .B1(new_n740), .B2(new_n853), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1129), .B1(new_n1130), .B2(new_n934), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(G330), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n846), .B2(new_n852), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n941), .A2(new_n947), .A3(new_n933), .A4(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n993), .A2(new_n475), .A3(new_n994), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n941), .A2(new_n947), .A3(new_n475), .A4(G330), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT115), .Z(new_n1140));
  AND3_X1   g0940(.A1(new_n1138), .A2(new_n1140), .A3(new_n667), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n762), .A2(new_n933), .A3(new_n1134), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1128), .A2(new_n1131), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1134), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n934), .B1(new_n960), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1130), .A2(new_n1142), .A3(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n934), .B1(new_n761), .B2(new_n1144), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1135), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1148), .A2(KEYINPUT116), .A3(new_n1122), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT116), .B1(new_n1148), .B2(new_n1122), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1146), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1137), .A2(new_n1141), .A3(new_n1143), .A4(new_n1152), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1128), .A2(new_n1131), .A3(new_n1142), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1135), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1151), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1145), .A2(new_n1142), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1156), .A2(new_n1149), .B1(new_n1130), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1138), .A2(new_n1140), .A3(new_n667), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n1154), .A2(new_n1155), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1153), .A2(new_n1160), .A3(new_n765), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT119), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n820), .A2(new_n568), .B1(new_n814), .B2(new_n481), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n871), .B(new_n1163), .C1(G294), .C2(new_n796), .ZN(new_n1164));
  INV_X1    g0964(.A(G283), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n807), .A2(new_n1165), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1098), .B(new_n1166), .C1(G107), .C2(new_n800), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n281), .B1(new_n818), .B2(new_n543), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT117), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1164), .A2(new_n1167), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n818), .A2(new_n435), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT53), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n820), .A2(new_n869), .B1(new_n792), .B2(new_n202), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G125), .B2(new_n796), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT54), .B(G143), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n279), .B1(new_n814), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G137), .B2(new_n800), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n811), .A2(G159), .B1(G128), .B2(new_n806), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1174), .A2(new_n1176), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1172), .A2(KEYINPUT118), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n783), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT118), .B1(new_n1172), .B2(new_n1181), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n769), .B1(new_n244), .B2(new_n861), .C1(new_n1183), .C2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n1121), .B2(new_n784), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1186), .B1(new_n1187), .B2(new_n768), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1161), .A2(new_n1162), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1162), .B1(new_n1161), .B2(new_n1188), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(G378));
  XNOR2_X1  g0992(.A(KEYINPUT123), .B(KEYINPUT55), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT121), .ZN(new_n1197));
  AOI221_X4 g0997(.A(new_n1197), .B1(new_n470), .B2(new_n472), .C1(new_n450), .C2(new_n463), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT121), .B1(new_n464), .B2(new_n473), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1196), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n449), .B1(new_n444), .B2(new_n448), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n462), .A2(KEYINPUT10), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n473), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n1197), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n464), .A2(KEYINPUT121), .A3(new_n473), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(new_n1205), .A3(new_n1195), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n471), .A2(new_n691), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AND3_X1   g1008(.A1(new_n1200), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1208), .B1(new_n1200), .B2(new_n1206), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1194), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1198), .A2(new_n1199), .A3(new_n1196), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1195), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1207), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1200), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1214), .A2(new_n1193), .A3(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1211), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n955), .B2(G330), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1133), .B(new_n1217), .C1(new_n950), .C2(new_n954), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n938), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1217), .B1(new_n959), .B2(new_n1133), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n955), .A2(G330), .A3(new_n1218), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n939), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1221), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n768), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n769), .B1(new_n861), .B2(G50), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT120), .Z(new_n1228));
  OAI22_X1  g1028(.A1(new_n801), .A2(new_n869), .B1(new_n810), .B2(new_n435), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1177), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(G128), .A2(new_n821), .B1(new_n819), .B2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n875), .B2(new_n814), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1229), .B(new_n1232), .C1(G125), .C2(new_n806), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n256), .B(new_n307), .C1(new_n792), .C2(new_n828), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G124), .B2(new_n796), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1235), .A2(new_n1236), .A3(new_n1238), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(G107), .A2(new_n821), .B1(new_n796), .B2(G283), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1022), .B2(new_n814), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n793), .A2(G58), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(G97), .A2(new_n800), .B1(new_n806), .B2(G116), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1066), .A2(new_n1242), .A3(new_n1243), .A4(new_n1039), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n776), .A2(new_n307), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1241), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1246), .A2(KEYINPUT58), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(KEYINPUT58), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1245), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1249));
  AND4_X1   g1049(.A1(new_n1239), .A2(new_n1247), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n1228), .B1(new_n860), .B2(new_n1250), .C1(new_n1218), .C2(new_n785), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1226), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1153), .A2(new_n1141), .B1(new_n1221), .B2(new_n1224), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n765), .B1(new_n1254), .B2(KEYINPUT57), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT124), .B1(new_n1256), .B2(new_n938), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1225), .B2(KEYINPUT124), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1159), .B1(new_n1187), .B2(new_n1152), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT57), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1253), .B1(new_n1255), .B2(new_n1261), .ZN(G375));
  INV_X1    g1062(.A(KEYINPUT125), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(new_n1158), .A2(new_n1263), .A3(new_n767), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT125), .B1(new_n1152), .B2(new_n768), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n769), .B1(new_n861), .B2(G68), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n933), .A2(new_n785), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(G97), .A2(new_n819), .B1(new_n796), .B2(G303), .ZN(new_n1268));
  OAI221_X1 g1068(.A(new_n1268), .B1(new_n418), .B2(new_n814), .C1(new_n1165), .C2(new_n820), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(G116), .A2(new_n800), .B1(new_n806), .B2(G294), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1036), .A2(new_n1270), .A3(new_n1069), .A4(new_n281), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(G137), .A2(new_n821), .B1(new_n819), .B2(G159), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(G58), .A2(new_n793), .B1(new_n796), .B2(G128), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n815), .A2(G150), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1272), .A2(new_n1273), .A3(new_n315), .A4(new_n1274), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(G50), .A2(new_n811), .B1(new_n1230), .B2(new_n800), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n869), .B2(new_n807), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n1269), .A2(new_n1271), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1266), .B(new_n1267), .C1(new_n783), .C2(new_n1278), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1264), .A2(new_n1265), .A3(new_n1279), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1141), .A2(new_n1152), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1152), .A2(new_n896), .A3(new_n1140), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1018), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1280), .B1(new_n1281), .B2(new_n1284), .ZN(G381));
  NAND3_X1  g1085(.A1(new_n1089), .A2(new_n840), .A3(new_n1091), .ZN(new_n1286));
  NOR4_X1   g1086(.A1(G390), .A2(new_n1286), .A3(G381), .A4(G384), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n992), .A2(new_n1019), .B1(new_n1021), .B2(new_n1047), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1137), .A2(new_n1143), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1141), .B1(new_n1289), .B2(new_n1282), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1225), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n712), .B1(new_n1291), .B2(new_n1260), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT124), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1293), .B1(new_n1221), .B2(new_n1224), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1290), .B(KEYINPUT57), .C1(new_n1257), .C2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1252), .B1(new_n1292), .B2(new_n1295), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1161), .A2(KEYINPUT126), .A3(new_n1188), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT126), .B1(new_n1161), .B2(new_n1188), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1287), .A2(new_n1288), .A3(new_n1296), .A4(new_n1299), .ZN(G407));
  NAND2_X1  g1100(.A1(new_n692), .A2(G213), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1296), .A2(new_n1299), .A3(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(G407), .A2(G213), .A3(new_n1303), .ZN(G409));
  NAND3_X1  g1104(.A1(new_n1290), .A2(new_n1283), .A3(new_n1225), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n768), .B1(new_n1294), .B2(new_n1257), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1305), .A2(new_n1251), .A3(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1161), .A2(new_n1188), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT126), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1161), .A2(KEYINPUT126), .A3(new_n1188), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1307), .A2(new_n1310), .A3(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1308), .A2(KEYINPUT119), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1189), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1312), .B1(G375), .B2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1281), .B1(KEYINPUT60), .B2(new_n1282), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1158), .A2(new_n1159), .A3(KEYINPUT60), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n765), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1280), .B1(new_n1316), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n883), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1280), .B(G384), .C1(new_n1316), .C2(new_n1318), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1315), .A2(new_n1301), .A3(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(KEYINPUT62), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1302), .A2(G2897), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1302), .A2(KEYINPUT127), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1320), .A2(new_n1321), .A3(new_n1326), .A4(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1320), .A2(new_n1321), .A3(new_n1327), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1329), .A2(G2897), .A3(new_n1302), .ZN(new_n1330));
  AOI22_X1  g1130(.A1(new_n1296), .A2(G378), .B1(new_n1299), .B2(new_n1307), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1328), .B(new_n1330), .C1(new_n1331), .C2(new_n1302), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT61), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT62), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1315), .A2(new_n1334), .A3(new_n1301), .A4(new_n1323), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1325), .A2(new_n1332), .A3(new_n1333), .A4(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1091), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1090), .B1(new_n1051), .B2(new_n1087), .ZN(new_n1338));
  OAI21_X1  g1138(.A(G396), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  AND3_X1   g1139(.A1(new_n1339), .A2(G390), .A3(new_n1286), .ZN(new_n1340));
  AOI21_X1  g1140(.A(G390), .B1(new_n1339), .B2(new_n1286), .ZN(new_n1341));
  OAI21_X1  g1141(.A(G387), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1339), .A2(new_n1286), .ZN(new_n1343));
  INV_X1    g1143(.A(G390), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1339), .A2(G390), .A3(new_n1286), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1345), .A2(new_n1288), .A3(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1342), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1336), .A2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT63), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1348), .B1(new_n1350), .B2(new_n1324), .ZN(new_n1351));
  OR2_X1    g1151(.A1(new_n1324), .A2(new_n1350), .ZN(new_n1352));
  XNOR2_X1  g1152(.A(new_n1329), .B(new_n1326), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1315), .A2(new_n1301), .ZN(new_n1354));
  AOI21_X1  g1154(.A(KEYINPUT61), .B1(new_n1353), .B2(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1351), .A2(new_n1352), .A3(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1349), .A2(new_n1356), .ZN(G405));
  NAND2_X1  g1157(.A1(new_n1296), .A2(G378), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(G375), .A2(new_n1299), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1358), .A2(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1360), .A2(new_n1323), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1358), .A2(new_n1359), .A3(new_n1322), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  XNOR2_X1  g1163(.A(new_n1363), .B(new_n1348), .ZN(G402));
endmodule


