//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n595,
    new_n598, new_n600, new_n601, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  AND3_X1   g043(.A1(new_n468), .A2(G101), .A3(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n469), .B1(new_n470), .B2(G137), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(G160));
  OAI21_X1  g047(.A(G2104), .B1(new_n468), .B2(G112), .ZN(new_n473));
  OR3_X1    g048(.A1(KEYINPUT67), .A2(G100), .A3(G2105), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT67), .B1(G100), .B2(G2105), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n468), .B1(new_n463), .B2(new_n464), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  AOI211_X1 g054(.A(new_n476), .B(new_n479), .C1(G136), .C2(new_n470), .ZN(G162));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  INV_X1    g056(.A(G138), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n484));
  NOR2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  AND2_X1   g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n483), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  XNOR2_X1  g063(.A(KEYINPUT3), .B(G2104), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n484), .B1(new_n489), .B2(new_n483), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n486), .C2(new_n485), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n481), .B1(new_n491), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n483), .B1(new_n486), .B2(new_n485), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(new_n487), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n492), .A2(new_n495), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT68), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  OR2_X1    g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n510), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  INV_X1    g095(.A(G89), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n522));
  INV_X1    g097(.A(G51), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n514), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n525));
  OAI221_X1 g100(.A(new_n520), .B1(new_n521), .B2(new_n512), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n526), .A2(new_n528), .ZN(G168));
  AOI22_X1  g104(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n509), .ZN(new_n531));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n512), .A2(new_n532), .B1(new_n514), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(G171));
  INV_X1    g110(.A(G81), .ZN(new_n536));
  INV_X1    g111(.A(G43), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n512), .A2(new_n536), .B1(new_n514), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT70), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n509), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  INV_X1    g123(.A(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(KEYINPUT6), .A2(G651), .ZN(new_n550));
  NAND2_X1  g125(.A1(KEYINPUT6), .A2(G651), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G53), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT9), .ZN(new_n554));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(new_n507), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n512), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n558), .A2(G651), .B1(new_n559), .B2(G91), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n554), .A2(new_n560), .ZN(G299));
  INV_X1    g136(.A(G171), .ZN(G301));
  INV_X1    g137(.A(G168), .ZN(G286));
  OAI21_X1  g138(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n564));
  INV_X1    g139(.A(G49), .ZN(new_n565));
  INV_X1    g140(.A(G87), .ZN(new_n566));
  OAI221_X1 g141(.A(new_n564), .B1(new_n514), .B2(new_n565), .C1(new_n566), .C2(new_n512), .ZN(G288));
  NAND2_X1  g142(.A1(new_n552), .A2(G48), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n507), .A2(new_n511), .A3(G86), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(G61), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(new_n505), .B2(new_n506), .ZN(new_n572));
  AND2_X1   g147(.A1(G73), .A2(G543), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(G305));
  AOI22_X1  g150(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(new_n509), .ZN(new_n577));
  INV_X1    g152(.A(G85), .ZN(new_n578));
  INV_X1    g153(.A(G47), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n512), .A2(new_n578), .B1(new_n514), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G290));
  NAND2_X1  g157(.A1(G301), .A2(G868), .ZN(new_n583));
  AND3_X1   g158(.A1(new_n507), .A2(new_n511), .A3(G92), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT10), .ZN(new_n585));
  NAND2_X1  g160(.A1(G79), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G66), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n556), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(G54), .B2(new_n552), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n583), .B1(new_n591), .B2(G868), .ZN(G321));
  XNOR2_X1  g167(.A(G321), .B(KEYINPUT71), .ZN(G284));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  NAND2_X1  g169(.A1(G299), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(G168), .B2(new_n594), .ZN(G297));
  OAI21_X1  g171(.A(new_n595), .B1(G168), .B2(new_n594), .ZN(G280));
  INV_X1    g172(.A(G559), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n591), .B1(new_n598), .B2(G860), .ZN(G148));
  NAND2_X1  g174(.A1(new_n542), .A2(new_n594), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n590), .A2(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(new_n594), .ZN(G323));
  XNOR2_X1  g177(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g178(.A(G2104), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(G2105), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n489), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g181(.A(KEYINPUT72), .B(KEYINPUT12), .Z(new_n607));
  XNOR2_X1  g182(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT13), .ZN(new_n609));
  XOR2_X1   g184(.A(KEYINPUT73), .B(G2100), .Z(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(KEYINPUT74), .Z(new_n612));
  NAND2_X1  g187(.A1(new_n470), .A2(G135), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n477), .A2(G123), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n468), .A2(G111), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(G2096), .Z(new_n618));
  OAI211_X1 g193(.A(new_n612), .B(new_n618), .C1(new_n610), .C2(new_n609), .ZN(G156));
  XNOR2_X1  g194(.A(G2427), .B(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT15), .B(G2435), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n623), .A2(KEYINPUT14), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2443), .B(G2446), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G1341), .B(G1348), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(G2451), .B(G2454), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT75), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n629), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(G14), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT76), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(G401));
  INV_X1    g212(.A(KEYINPUT18), .ZN(new_n638));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT17), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n639), .A2(new_n640), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n638), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2100), .ZN(new_n645));
  XOR2_X1   g220(.A(G2072), .B(G2078), .Z(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(new_n641), .B2(KEYINPUT18), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2096), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n645), .B(new_n648), .ZN(G227));
  XOR2_X1   g224(.A(G1971), .B(G1976), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT19), .ZN(new_n651));
  XOR2_X1   g226(.A(G1956), .B(G2474), .Z(new_n652));
  XOR2_X1   g227(.A(G1961), .B(G1966), .Z(new_n653));
  AND2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT20), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n652), .A2(new_n653), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  MUX2_X1   g234(.A(new_n659), .B(new_n658), .S(new_n651), .Z(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT77), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n661), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G1991), .B(G1996), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT78), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1981), .B(G1986), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G229));
  INV_X1    g244(.A(G29), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n670), .A2(G32), .ZN(new_n671));
  NAND3_X1  g246(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT26), .Z(new_n673));
  NAND2_X1  g248(.A1(new_n470), .A2(G141), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n477), .A2(G129), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n605), .A2(G105), .ZN(new_n676));
  NAND4_X1  g251(.A1(new_n673), .A2(new_n674), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n671), .B1(new_n677), .B2(G29), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT86), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT27), .B(G1996), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT87), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n670), .A2(G33), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT25), .ZN(new_n685));
  AOI22_X1  g260(.A1(new_n489), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n686), .A2(new_n468), .ZN(new_n687));
  AOI211_X1 g262(.A(new_n685), .B(new_n687), .C1(G139), .C2(new_n470), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n683), .B1(new_n688), .B2(new_n670), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(G2072), .Z(new_n690));
  INV_X1    g265(.A(G34), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n691), .A2(KEYINPUT24), .ZN(new_n692));
  AOI21_X1  g267(.A(G29), .B1(new_n691), .B2(KEYINPUT24), .ZN(new_n693));
  AOI22_X1  g268(.A1(G160), .A2(G29), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G2084), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT85), .Z(new_n696));
  NAND3_X1  g271(.A1(new_n682), .A2(new_n690), .A3(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT88), .Z(new_n698));
  NAND2_X1  g273(.A1(new_n670), .A2(G35), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G162), .B2(new_n670), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT29), .Z(new_n701));
  INV_X1    g276(.A(G2090), .ZN(new_n702));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G21), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G168), .B2(new_n703), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n701), .A2(new_n702), .B1(G1966), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(G5), .A2(G16), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT89), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G301), .B2(new_n703), .ZN(new_n709));
  INV_X1    g284(.A(G1961), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G2084), .B2(new_n694), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n679), .A2(new_n680), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n709), .A2(new_n710), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT31), .B(G11), .ZN(new_n715));
  INV_X1    g290(.A(G28), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(KEYINPUT30), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT30), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n670), .B1(new_n718), .B2(G28), .ZN(new_n719));
  OAI221_X1 g294(.A(new_n715), .B1(new_n717), .B2(new_n719), .C1(new_n617), .C2(new_n670), .ZN(new_n720));
  NOR4_X1   g295(.A1(new_n712), .A2(new_n713), .A3(new_n714), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n706), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n670), .A2(G27), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G164), .B2(new_n670), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G2078), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n670), .A2(G26), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT84), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT28), .ZN(new_n728));
  AOI22_X1  g303(.A1(G128), .A2(new_n477), .B1(new_n470), .B2(G140), .ZN(new_n729));
  INV_X1    g304(.A(G104), .ZN(new_n730));
  AND3_X1   g305(.A1(new_n730), .A2(new_n468), .A3(KEYINPUT83), .ZN(new_n731));
  AOI21_X1  g306(.A(KEYINPUT83), .B1(new_n730), .B2(new_n468), .ZN(new_n732));
  OAI221_X1 g307(.A(G2104), .B1(G116), .B2(new_n468), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n728), .B1(new_n735), .B2(new_n670), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G2067), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n703), .A2(G20), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT23), .Z(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G299), .B2(G16), .ZN(new_n740));
  INV_X1    g315(.A(G1956), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NOR4_X1   g317(.A1(new_n722), .A2(new_n725), .A3(new_n737), .A4(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G16), .A2(G19), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n543), .B2(G16), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT82), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(G1341), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n703), .A2(G4), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n591), .B2(new_n703), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT81), .B(G1348), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  OAI221_X1 g326(.A(new_n751), .B1(G1966), .B2(new_n705), .C1(new_n701), .C2(new_n702), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n746), .B2(G1341), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n698), .A2(new_n743), .A3(new_n747), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n703), .A2(G22), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G166), .B2(new_n703), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1971), .ZN(new_n757));
  NOR2_X1   g332(.A1(G6), .A2(G16), .ZN(new_n758));
  INV_X1    g333(.A(G305), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(G16), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT32), .B(G1981), .Z(new_n761));
  XOR2_X1   g336(.A(new_n760), .B(new_n761), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n703), .A2(G23), .ZN(new_n763));
  INV_X1    g338(.A(G288), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n703), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT33), .B(G1976), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n765), .B(new_n766), .Z(new_n767));
  NOR3_X1   g342(.A1(new_n757), .A2(new_n762), .A3(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT34), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n470), .A2(G131), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n477), .A2(G119), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n468), .A2(G107), .ZN(new_n773));
  OAI21_X1  g348(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n771), .B(new_n772), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  MUX2_X1   g350(.A(G25), .B(new_n775), .S(G29), .Z(new_n776));
  XOR2_X1   g351(.A(KEYINPUT35), .B(G1991), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n778), .A2(KEYINPUT79), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n778), .A2(KEYINPUT79), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n703), .A2(G24), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n581), .B2(new_n703), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1986), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n779), .A2(new_n780), .A3(new_n783), .ZN(new_n784));
  AND3_X1   g359(.A1(new_n770), .A2(KEYINPUT80), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(KEYINPUT80), .B1(new_n770), .B2(new_n784), .ZN(new_n786));
  OAI22_X1  g361(.A1(new_n785), .A2(new_n786), .B1(new_n769), .B2(new_n768), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT36), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(KEYINPUT36), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n754), .B1(new_n788), .B2(new_n789), .ZN(G311));
  XOR2_X1   g365(.A(G311), .B(KEYINPUT90), .Z(G150));
  NAND2_X1  g366(.A1(new_n542), .A2(KEYINPUT92), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(new_n509), .ZN(new_n794));
  INV_X1    g369(.A(G93), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT91), .B(G55), .Z(new_n796));
  OAI22_X1  g371(.A1(new_n512), .A2(new_n795), .B1(new_n514), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT92), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n539), .A2(new_n799), .A3(new_n541), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n792), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n542), .B(KEYINPUT92), .C1(new_n794), .C2(new_n797), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT38), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n591), .A2(G559), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(KEYINPUT39), .ZN(new_n807));
  INV_X1    g382(.A(G860), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(KEYINPUT39), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n798), .A2(new_n808), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT37), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n812), .ZN(G145));
  AOI21_X1  g388(.A(new_n496), .B1(new_n499), .B2(new_n487), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n734), .B(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n677), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(new_n688), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n608), .B(new_n775), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n477), .A2(G130), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n468), .A2(G118), .ZN(new_n821));
  OAI21_X1  g396(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(G142), .B2(new_n470), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n819), .B(new_n824), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n818), .A2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT93), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n818), .B2(new_n825), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n826), .A2(new_n828), .ZN(new_n830));
  XNOR2_X1  g405(.A(G160), .B(new_n617), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G162), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n832), .B1(new_n818), .B2(new_n825), .ZN(new_n834));
  AOI21_X1  g409(.A(G37), .B1(new_n826), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g412(.A(KEYINPUT97), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n798), .A2(G868), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT94), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n590), .A2(G299), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n590), .A2(G299), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n841), .B1(new_n844), .B2(KEYINPUT41), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT41), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n844), .B(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n846), .B1(new_n848), .B2(KEYINPUT94), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n803), .B(new_n601), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n844), .B2(new_n850), .ZN(new_n852));
  NAND2_X1  g427(.A1(KEYINPUT96), .A2(KEYINPUT42), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n581), .B(G288), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(KEYINPUT95), .ZN(new_n856));
  XNOR2_X1  g431(.A(G303), .B(G305), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n855), .A2(KEYINPUT95), .ZN(new_n859));
  MUX2_X1   g434(.A(new_n858), .B(new_n857), .S(new_n859), .Z(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(KEYINPUT96), .B2(KEYINPUT42), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n854), .A2(new_n862), .ZN(new_n863));
  AND3_X1   g438(.A1(new_n852), .A2(KEYINPUT96), .A3(KEYINPUT42), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n852), .B1(KEYINPUT96), .B2(KEYINPUT42), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n838), .B(new_n840), .C1(new_n867), .C2(new_n594), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n594), .B1(new_n863), .B2(new_n866), .ZN(new_n869));
  OAI21_X1  g444(.A(KEYINPUT97), .B1(new_n869), .B2(new_n839), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(G295));
  OAI21_X1  g446(.A(new_n840), .B1(new_n867), .B2(new_n594), .ZN(G331));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n873));
  INV_X1    g448(.A(new_n844), .ZN(new_n874));
  OAI21_X1  g449(.A(G301), .B1(new_n526), .B2(new_n528), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n524), .A2(new_n525), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n520), .B1(new_n512), .B2(new_n521), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(new_n527), .A3(G171), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n801), .A2(new_n802), .A3(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n882), .A2(KEYINPUT100), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n803), .A2(new_n880), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(KEYINPUT100), .ZN(new_n885));
  AND4_X1   g460(.A1(new_n874), .A2(new_n883), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n882), .A2(KEYINPUT98), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT98), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n801), .A2(new_n888), .A3(new_n802), .A4(new_n881), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n884), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(KEYINPUT99), .A3(new_n849), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT99), .ZN(new_n893));
  AOI22_X1  g468(.A1(new_n887), .A2(new_n889), .B1(new_n803), .B2(new_n880), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n844), .B(KEYINPUT41), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n845), .B1(new_n895), .B2(new_n841), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n893), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n886), .B1(new_n892), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n860), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n895), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n890), .A2(new_n874), .A3(new_n884), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n860), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n903), .A2(G37), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n899), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n899), .ZN(new_n907));
  INV_X1    g482(.A(G37), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(new_n898), .B2(new_n860), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT101), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT101), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n911), .B(new_n908), .C1(new_n898), .C2(new_n860), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n907), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n873), .B(new_n906), .C1(new_n913), .C2(new_n905), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n899), .A2(new_n905), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n915), .B1(new_n910), .B2(new_n912), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n905), .B1(new_n899), .B2(new_n904), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT44), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n914), .A2(new_n918), .ZN(G397));
  NAND3_X1  g494(.A1(new_n467), .A2(new_n471), .A3(G40), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n467), .A2(new_n471), .A3(KEYINPUT103), .A4(G40), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n500), .A2(new_n501), .ZN(new_n925));
  XOR2_X1   g500(.A(KEYINPUT102), .B(G1384), .Z(new_n926));
  AOI21_X1  g501(.A(KEYINPUT45), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n734), .B(G2067), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT104), .ZN(new_n930));
  INV_X1    g505(.A(G1996), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n677), .B(new_n931), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n775), .B(new_n777), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n581), .B(G1986), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n928), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(KEYINPUT107), .B(G8), .Z(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(G286), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  OR2_X1    g517(.A1(new_n942), .A2(KEYINPUT51), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n944));
  INV_X1    g519(.A(G1384), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n925), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n944), .B1(new_n946), .B2(KEYINPUT50), .ZN(new_n947));
  AOI21_X1  g522(.A(G1384), .B1(new_n497), .B2(new_n502), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT50), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n500), .A2(KEYINPUT68), .A3(new_n501), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT68), .B1(new_n500), .B2(new_n501), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n945), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n953), .A2(new_n944), .A3(KEYINPUT50), .ZN(new_n954));
  XOR2_X1   g529(.A(KEYINPUT113), .B(G2084), .Z(new_n955));
  NAND4_X1  g530(.A1(new_n950), .A2(new_n954), .A3(new_n924), .A4(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G1966), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(G1384), .B1(new_n500), .B2(new_n501), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n922), .B(new_n923), .C1(KEYINPUT45), .C2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n957), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n956), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n940), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT122), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n943), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n963), .A2(KEYINPUT122), .A3(new_n940), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(KEYINPUT120), .B(KEYINPUT51), .ZN(new_n969));
  INV_X1    g544(.A(G8), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n970), .B1(new_n956), .B2(new_n962), .ZN(new_n971));
  OAI211_X1 g546(.A(KEYINPUT121), .B(new_n969), .C1(new_n971), .C2(new_n942), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n969), .B1(new_n971), .B2(new_n942), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT121), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n968), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n963), .A2(new_n942), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT45), .B1(new_n503), .B2(new_n945), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n925), .A2(new_n926), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n922), .B(new_n923), .C1(new_n980), .C2(new_n958), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G2078), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n950), .A2(new_n924), .A3(new_n954), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n984), .A2(new_n985), .B1(new_n986), .B2(new_n710), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n988));
  OR4_X1    g563(.A1(new_n988), .A2(new_n959), .A3(new_n961), .A4(G2078), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  XOR2_X1   g565(.A(G171), .B(KEYINPUT54), .Z(new_n991));
  AND2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n922), .A2(new_n923), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n960), .A2(new_n949), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT111), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n503), .A2(new_n949), .A3(new_n945), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT50), .B1(new_n814), .B2(G1384), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n997), .A2(new_n998), .A3(new_n922), .A4(new_n923), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n995), .A2(new_n702), .A3(new_n996), .A4(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1971), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n979), .B2(new_n981), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n940), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(G166), .B2(new_n970), .ZN(new_n1006));
  NAND3_X1  g581(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1004), .A2(KEYINPUT112), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n939), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1011), .B1(new_n1012), .B2(new_n1008), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n950), .A2(new_n954), .A3(new_n702), .A4(new_n924), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n970), .B1(new_n1014), .B2(new_n1002), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1006), .A2(KEYINPUT106), .A3(new_n1007), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT106), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n922), .A2(new_n960), .A3(new_n923), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n764), .A2(G1976), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1020), .A2(new_n1021), .A3(new_n940), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT52), .ZN(new_n1023));
  INV_X1    g598(.A(G1981), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n570), .A2(KEYINPUT109), .A3(new_n1024), .A4(new_n574), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n574), .A2(new_n1024), .A3(new_n569), .A4(new_n568), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT109), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n1025), .A2(new_n1028), .B1(G305), .B2(G1981), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT49), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1020), .B(new_n940), .C1(new_n1029), .C2(KEYINPUT49), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1023), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G1976), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT52), .B1(G288), .B2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1020), .A2(new_n1021), .A3(new_n940), .A4(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT108), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1033), .A2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1010), .A2(new_n1013), .A3(new_n1019), .A4(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n920), .A2(KEYINPUT124), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n920), .A2(KEYINPUT124), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1041), .A2(new_n927), .A3(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n980), .A2(new_n958), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n1044), .A2(new_n988), .A3(G2078), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n991), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n987), .A2(new_n1046), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n992), .A2(new_n1040), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n978), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n981), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n953), .A2(new_n958), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(new_n1052), .A3(new_n931), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n1054));
  XOR2_X1   g629(.A(KEYINPUT58), .B(G1341), .Z(new_n1055));
  NAND2_X1  g630(.A1(new_n1020), .A2(new_n1055), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1053), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1054), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n543), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1059), .B(new_n1062), .ZN(new_n1063));
  XOR2_X1   g638(.A(G299), .B(KEYINPUT57), .Z(new_n1064));
  INV_X1    g639(.A(new_n995), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n996), .A2(new_n999), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n741), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT56), .B(G2072), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n982), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1064), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1067), .A2(new_n1064), .A3(new_n1069), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(KEYINPUT61), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1067), .A2(new_n1069), .A3(KEYINPUT115), .A4(new_n1064), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1070), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1063), .B(new_n1073), .C1(KEYINPUT61), .C2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT60), .ZN(new_n1079));
  INV_X1    g654(.A(new_n750), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n953), .A2(KEYINPUT50), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n993), .B1(new_n1081), .B2(new_n947), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1080), .B1(new_n1082), .B2(new_n954), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1020), .A2(G2067), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT116), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n986), .B2(new_n750), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1079), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1089), .A2(new_n1090), .A3(new_n591), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1093));
  AOI211_X1 g668(.A(KEYINPUT116), .B(new_n1084), .C1(new_n986), .C2(new_n750), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT60), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n590), .B1(new_n1095), .B2(KEYINPUT119), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1091), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1085), .A2(new_n1088), .A3(new_n1079), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1078), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1093), .A2(new_n1094), .A3(new_n590), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(new_n1070), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1101), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1050), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1015), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n1009), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT63), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1107), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n963), .A2(G168), .A3(new_n940), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1106), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT110), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n1033), .B2(new_n1038), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1036), .B(KEYINPUT108), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1020), .A2(new_n940), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1029), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT49), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n1030), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1114), .A2(new_n1119), .A3(KEYINPUT110), .A4(new_n1023), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1113), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1104), .B1(new_n1111), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1107), .B1(new_n1040), .B2(new_n1109), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1109), .B1(new_n1009), .B2(new_n1105), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1113), .A2(new_n1120), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(KEYINPUT114), .A3(new_n1125), .A4(new_n1108), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1122), .A2(new_n1123), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1119), .A2(new_n1034), .A3(new_n764), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1115), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1019), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1130), .B1(new_n1125), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1127), .A2(new_n1132), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n966), .A2(new_n967), .B1(new_n973), .B2(new_n974), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1134), .A2(new_n972), .B1(new_n942), .B2(new_n963), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n990), .A2(G171), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1040), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n978), .B2(KEYINPUT62), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1133), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n938), .B1(new_n1103), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n928), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1144), .A2(KEYINPUT46), .A3(new_n931), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT46), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n928), .B2(G1996), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n930), .A2(new_n816), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1145), .B(new_n1147), .C1(new_n1148), .C2(new_n928), .ZN(new_n1149));
  XOR2_X1   g724(.A(new_n1149), .B(KEYINPUT47), .Z(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n777), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n775), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n933), .A2(new_n1153), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n734), .A2(G2067), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n928), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n935), .A2(new_n1144), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n928), .A2(G1986), .A3(G290), .ZN(new_n1158));
  XNOR2_X1  g733(.A(KEYINPUT125), .B(KEYINPUT48), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1158), .B(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1156), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1151), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT126), .B1(new_n1143), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n938), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n1077), .A2(KEYINPUT61), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1063), .A2(new_n1073), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n591), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1095), .A2(KEYINPUT119), .A3(new_n590), .ZN(new_n1168));
  AOI22_X1  g743(.A1(new_n1167), .A2(new_n1168), .B1(new_n1090), .B2(new_n1089), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1098), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1165), .B(new_n1166), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1102), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1049), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1139), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n1175));
  OAI211_X1 g750(.A(new_n1127), .B(new_n1132), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1164), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1162), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1163), .A2(new_n1180), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g756(.A(new_n906), .B1(new_n913), .B2(new_n905), .ZN(new_n1183));
  NOR3_X1   g757(.A1(G229), .A2(new_n460), .A3(G227), .ZN(new_n1184));
  NAND2_X1  g758(.A1(new_n1184), .A2(new_n636), .ZN(new_n1185));
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n1186));
  XNOR2_X1  g760(.A(new_n1185), .B(new_n1186), .ZN(new_n1187));
  AND3_X1   g761(.A1(new_n1183), .A2(new_n836), .A3(new_n1187), .ZN(G308));
  NAND3_X1  g762(.A1(new_n1183), .A2(new_n836), .A3(new_n1187), .ZN(G225));
endmodule


