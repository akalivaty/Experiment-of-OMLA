

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594;

  XNOR2_X1 U327 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U328 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U329 ( .A(n398), .B(n397), .ZN(n401) );
  XNOR2_X1 U330 ( .A(n414), .B(n413), .ZN(n415) );
  INV_X1 U331 ( .A(KEYINPUT36), .ZN(n425) );
  XNOR2_X1 U332 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n455) );
  XNOR2_X1 U333 ( .A(n550), .B(n425), .ZN(n591) );
  XNOR2_X1 U334 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U335 ( .A(n311), .B(n310), .Z(n539) );
  XNOR2_X1 U336 ( .A(n330), .B(n329), .ZN(n557) );
  XNOR2_X1 U337 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n460) );
  XNOR2_X1 U338 ( .A(n461), .B(n460), .ZN(G1351GAT) );
  XOR2_X1 U339 ( .A(G169GAT), .B(G113GAT), .Z(n367) );
  XOR2_X1 U340 ( .A(G190GAT), .B(G134GAT), .Z(n408) );
  XNOR2_X1 U341 ( .A(n367), .B(n408), .ZN(n297) );
  XOR2_X1 U342 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n296) );
  XNOR2_X1 U343 ( .A(KEYINPUT88), .B(KEYINPUT18), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n335) );
  XNOR2_X1 U345 ( .A(n297), .B(n335), .ZN(n303) );
  XOR2_X1 U346 ( .A(G120GAT), .B(G127GAT), .Z(n299) );
  XNOR2_X1 U347 ( .A(KEYINPUT85), .B(KEYINPUT0), .ZN(n298) );
  XNOR2_X1 U348 ( .A(n299), .B(n298), .ZN(n328) );
  XOR2_X1 U349 ( .A(G15GAT), .B(n328), .Z(n301) );
  NAND2_X1 U350 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U352 ( .A(n303), .B(n302), .Z(n311) );
  XOR2_X1 U353 ( .A(KEYINPUT86), .B(G71GAT), .Z(n305) );
  XNOR2_X1 U354 ( .A(G43GAT), .B(G99GAT), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U356 ( .A(G176GAT), .B(G183GAT), .Z(n307) );
  XNOR2_X1 U357 ( .A(KEYINPUT20), .B(KEYINPUT87), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U359 ( .A(n309), .B(n308), .ZN(n310) );
  INV_X1 U360 ( .A(n539), .ZN(n467) );
  XOR2_X1 U361 ( .A(KEYINPUT78), .B(G85GAT), .Z(n313) );
  XNOR2_X1 U362 ( .A(G29GAT), .B(G134GAT), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U364 ( .A(G155GAT), .B(G148GAT), .Z(n315) );
  XNOR2_X1 U365 ( .A(G113GAT), .B(G162GAT), .ZN(n314) );
  XNOR2_X1 U366 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U367 ( .A(n317), .B(n316), .Z(n322) );
  XOR2_X1 U368 ( .A(KEYINPUT1), .B(G57GAT), .Z(n319) );
  NAND2_X1 U369 ( .A1(G225GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U370 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U371 ( .A(KEYINPUT6), .B(n320), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U373 ( .A(KEYINPUT4), .B(KEYINPUT92), .Z(n324) );
  XNOR2_X1 U374 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U376 ( .A(n326), .B(n325), .Z(n330) );
  XNOR2_X1 U377 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n327), .B(KEYINPUT2), .ZN(n450) );
  XNOR2_X1 U379 ( .A(n328), .B(n450), .ZN(n329) );
  INV_X1 U380 ( .A(KEYINPUT54), .ZN(n433) );
  XOR2_X1 U381 ( .A(G92GAT), .B(G218GAT), .Z(n332) );
  XNOR2_X1 U382 ( .A(G36GAT), .B(G190GAT), .ZN(n331) );
  XNOR2_X1 U383 ( .A(n332), .B(n331), .ZN(n346) );
  XOR2_X1 U384 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n334) );
  XNOR2_X1 U385 ( .A(G169GAT), .B(KEYINPUT93), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n334), .B(n333), .ZN(n339) );
  XOR2_X1 U387 ( .A(G64GAT), .B(n335), .Z(n337) );
  NAND2_X1 U388 ( .A1(G226GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U389 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U390 ( .A(n339), .B(n338), .ZN(n344) );
  XOR2_X1 U391 ( .A(G197GAT), .B(KEYINPUT21), .Z(n437) );
  XOR2_X1 U392 ( .A(KEYINPUT80), .B(G211GAT), .Z(n341) );
  XNOR2_X1 U393 ( .A(G8GAT), .B(G183GAT), .ZN(n340) );
  XNOR2_X1 U394 ( .A(n341), .B(n340), .ZN(n360) );
  XNOR2_X1 U395 ( .A(n437), .B(n360), .ZN(n342) );
  XOR2_X1 U396 ( .A(G176GAT), .B(G204GAT), .Z(n394) );
  XNOR2_X1 U397 ( .A(n342), .B(n394), .ZN(n343) );
  XNOR2_X1 U398 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U399 ( .A(n346), .B(n345), .Z(n525) );
  INV_X1 U400 ( .A(n525), .ZN(n466) );
  XOR2_X1 U401 ( .A(KEYINPUT13), .B(KEYINPUT71), .Z(n348) );
  XNOR2_X1 U402 ( .A(G71GAT), .B(G57GAT), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U404 ( .A(G64GAT), .B(n349), .ZN(n403) );
  XOR2_X1 U405 ( .A(G22GAT), .B(G155GAT), .Z(n438) );
  XOR2_X1 U406 ( .A(KEYINPUT12), .B(KEYINPUT81), .Z(n351) );
  XNOR2_X1 U407 ( .A(G127GAT), .B(G78GAT), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U409 ( .A(n438), .B(n352), .Z(n354) );
  NAND2_X1 U410 ( .A1(G231GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U412 ( .A(KEYINPUT82), .B(KEYINPUT14), .Z(n356) );
  XNOR2_X1 U413 ( .A(KEYINPUT83), .B(KEYINPUT15), .ZN(n355) );
  XNOR2_X1 U414 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U415 ( .A(n358), .B(n357), .Z(n362) );
  XNOR2_X1 U416 ( .A(G15GAT), .B(G1GAT), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n359), .B(KEYINPUT68), .ZN(n370) );
  XNOR2_X1 U418 ( .A(n370), .B(n360), .ZN(n361) );
  XNOR2_X1 U419 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U420 ( .A(n403), .B(n363), .Z(n463) );
  INV_X1 U421 ( .A(n463), .ZN(n588) );
  XOR2_X1 U422 ( .A(KEYINPUT114), .B(n588), .Z(n546) );
  XOR2_X1 U423 ( .A(KEYINPUT64), .B(KEYINPUT65), .Z(n365) );
  XNOR2_X1 U424 ( .A(G197GAT), .B(G8GAT), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U426 ( .A(n366), .B(G22GAT), .Z(n369) );
  XNOR2_X1 U427 ( .A(n367), .B(G141GAT), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n374) );
  XOR2_X1 U429 ( .A(KEYINPUT69), .B(n370), .Z(n372) );
  NAND2_X1 U430 ( .A1(G229GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U432 ( .A(n374), .B(n373), .Z(n383) );
  XNOR2_X1 U433 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n375), .B(G29GAT), .ZN(n376) );
  XOR2_X1 U435 ( .A(n376), .B(KEYINPUT8), .Z(n378) );
  XNOR2_X1 U436 ( .A(G43GAT), .B(G50GAT), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n378), .B(n377), .ZN(n418) );
  XOR2_X1 U438 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n380) );
  XNOR2_X1 U439 ( .A(KEYINPUT29), .B(KEYINPUT66), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n418), .B(n381), .ZN(n382) );
  XNOR2_X1 U442 ( .A(n383), .B(n382), .ZN(n579) );
  INV_X1 U443 ( .A(KEYINPUT41), .ZN(n405) );
  XOR2_X1 U444 ( .A(KEYINPUT73), .B(G92GAT), .Z(n385) );
  XNOR2_X1 U445 ( .A(G99GAT), .B(G85GAT), .ZN(n384) );
  XNOR2_X1 U446 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U447 ( .A(G106GAT), .B(n386), .ZN(n419) );
  XNOR2_X1 U448 ( .A(G120GAT), .B(KEYINPUT32), .ZN(n392) );
  INV_X1 U449 ( .A(KEYINPUT74), .ZN(n387) );
  NAND2_X1 U450 ( .A1(KEYINPUT31), .A2(n387), .ZN(n390) );
  INV_X1 U451 ( .A(KEYINPUT31), .ZN(n388) );
  NAND2_X1 U452 ( .A1(n388), .A2(KEYINPUT74), .ZN(n389) );
  NAND2_X1 U453 ( .A1(n390), .A2(n389), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U455 ( .A(n394), .B(n393), .ZN(n398) );
  AND2_X1 U456 ( .A1(G230GAT), .A2(G233GAT), .ZN(n396) );
  INV_X1 U457 ( .A(KEYINPUT75), .ZN(n395) );
  XNOR2_X1 U458 ( .A(G78GAT), .B(KEYINPUT72), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n399), .B(G148GAT), .ZN(n443) );
  XNOR2_X1 U460 ( .A(n443), .B(KEYINPUT33), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U462 ( .A(n419), .B(n402), .Z(n404) );
  XOR2_X1 U463 ( .A(n404), .B(n403), .Z(n584) );
  XNOR2_X1 U464 ( .A(n405), .B(n584), .ZN(n510) );
  NOR2_X1 U465 ( .A1(n579), .A2(n510), .ZN(n406) );
  XNOR2_X1 U466 ( .A(n406), .B(KEYINPUT46), .ZN(n407) );
  NOR2_X1 U467 ( .A1(n546), .A2(n407), .ZN(n422) );
  XOR2_X1 U468 ( .A(KEYINPUT9), .B(KEYINPUT78), .Z(n410) );
  XOR2_X1 U469 ( .A(G218GAT), .B(G162GAT), .Z(n442) );
  XNOR2_X1 U470 ( .A(n408), .B(n442), .ZN(n409) );
  XNOR2_X1 U471 ( .A(n410), .B(n409), .ZN(n416) );
  XOR2_X1 U472 ( .A(KEYINPUT77), .B(KEYINPUT11), .Z(n412) );
  XNOR2_X1 U473 ( .A(KEYINPUT76), .B(KEYINPUT10), .ZN(n411) );
  XNOR2_X1 U474 ( .A(n412), .B(n411), .ZN(n414) );
  AND2_X1 U475 ( .A1(G232GAT), .A2(G233GAT), .ZN(n413) );
  XOR2_X1 U476 ( .A(n418), .B(n417), .Z(n421) );
  INV_X1 U477 ( .A(n419), .ZN(n420) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n566) );
  NAND2_X1 U479 ( .A1(n422), .A2(n566), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n423), .B(KEYINPUT47), .ZN(n430) );
  INV_X1 U481 ( .A(KEYINPUT79), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n424), .B(n566), .ZN(n462) );
  INV_X1 U483 ( .A(n462), .ZN(n550) );
  NOR2_X1 U484 ( .A1(n591), .A2(n588), .ZN(n426) );
  XNOR2_X1 U485 ( .A(KEYINPUT45), .B(n426), .ZN(n427) );
  NAND2_X1 U486 ( .A1(n427), .A2(n584), .ZN(n428) );
  XOR2_X1 U487 ( .A(n579), .B(KEYINPUT70), .Z(n568) );
  NOR2_X1 U488 ( .A1(n428), .A2(n568), .ZN(n429) );
  NOR2_X1 U489 ( .A1(n430), .A2(n429), .ZN(n431) );
  XNOR2_X1 U490 ( .A(n431), .B(KEYINPUT48), .ZN(n555) );
  NOR2_X1 U491 ( .A1(n466), .A2(n555), .ZN(n432) );
  XNOR2_X1 U492 ( .A(n433), .B(n432), .ZN(n434) );
  NOR2_X1 U493 ( .A1(n557), .A2(n434), .ZN(n578) );
  XOR2_X1 U494 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n436) );
  XNOR2_X1 U495 ( .A(KEYINPUT24), .B(KEYINPUT91), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n454) );
  XOR2_X1 U497 ( .A(G211GAT), .B(G204GAT), .Z(n440) );
  XNOR2_X1 U498 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U499 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U500 ( .A(n441), .B(G106GAT), .Z(n448) );
  XOR2_X1 U501 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U502 ( .A1(G228GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U503 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U504 ( .A(G50GAT), .B(n446), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U506 ( .A(n449), .B(KEYINPUT90), .Z(n452) );
  XNOR2_X1 U507 ( .A(n450), .B(KEYINPUT89), .ZN(n451) );
  XNOR2_X1 U508 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U509 ( .A(n454), .B(n453), .Z(n477) );
  NAND2_X1 U510 ( .A1(n578), .A2(n477), .ZN(n456) );
  NOR2_X1 U511 ( .A1(n467), .A2(n457), .ZN(n574) );
  NAND2_X1 U512 ( .A1(n574), .A2(n546), .ZN(n459) );
  XNOR2_X1 U513 ( .A(G183GAT), .B(KEYINPUT124), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n459), .B(n458), .ZN(G1350GAT) );
  NAND2_X1 U515 ( .A1(n574), .A2(n550), .ZN(n461) );
  XNOR2_X1 U516 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n485) );
  NAND2_X1 U517 ( .A1(n568), .A2(n584), .ZN(n498) );
  XOR2_X1 U518 ( .A(KEYINPUT84), .B(KEYINPUT16), .Z(n465) );
  NAND2_X1 U519 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U520 ( .A(n465), .B(n464), .ZN(n483) );
  NOR2_X1 U521 ( .A1(n467), .A2(n466), .ZN(n468) );
  XOR2_X1 U522 ( .A(KEYINPUT98), .B(n468), .Z(n469) );
  NAND2_X1 U523 ( .A1(n477), .A2(n469), .ZN(n470) );
  XNOR2_X1 U524 ( .A(KEYINPUT25), .B(n470), .ZN(n475) );
  NOR2_X1 U525 ( .A1(n477), .A2(n539), .ZN(n472) );
  XNOR2_X1 U526 ( .A(KEYINPUT26), .B(KEYINPUT96), .ZN(n471) );
  XNOR2_X1 U527 ( .A(n472), .B(n471), .ZN(n577) );
  XOR2_X1 U528 ( .A(KEYINPUT27), .B(n525), .Z(n478) );
  INV_X1 U529 ( .A(n478), .ZN(n473) );
  NAND2_X1 U530 ( .A1(n577), .A2(n473), .ZN(n554) );
  XNOR2_X1 U531 ( .A(KEYINPUT97), .B(n554), .ZN(n474) );
  NOR2_X1 U532 ( .A1(n475), .A2(n474), .ZN(n476) );
  NOR2_X1 U533 ( .A1(n557), .A2(n476), .ZN(n481) );
  XOR2_X1 U534 ( .A(n477), .B(KEYINPUT28), .Z(n532) );
  NOR2_X1 U535 ( .A1(n478), .A2(n532), .ZN(n479) );
  NAND2_X1 U536 ( .A1(n557), .A2(n479), .ZN(n537) );
  NOR2_X1 U537 ( .A1(n539), .A2(n537), .ZN(n480) );
  NOR2_X1 U538 ( .A1(n481), .A2(n480), .ZN(n495) );
  INV_X1 U539 ( .A(n495), .ZN(n482) );
  NAND2_X1 U540 ( .A1(n483), .A2(n482), .ZN(n512) );
  NOR2_X1 U541 ( .A1(n498), .A2(n512), .ZN(n492) );
  NAND2_X1 U542 ( .A1(n557), .A2(n492), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(G1324GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n487) );
  NAND2_X1 U545 ( .A1(n492), .A2(n525), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U547 ( .A(G8GAT), .B(n488), .ZN(G1325GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U549 ( .A1(n492), .A2(n539), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U551 ( .A(G15GAT), .B(n491), .Z(G1326GAT) );
  NAND2_X1 U552 ( .A1(n492), .A2(n532), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n493), .B(KEYINPUT102), .ZN(n494) );
  XNOR2_X1 U554 ( .A(G22GAT), .B(n494), .ZN(G1327GAT) );
  NOR2_X1 U555 ( .A1(n591), .A2(n495), .ZN(n496) );
  NAND2_X1 U556 ( .A1(n588), .A2(n496), .ZN(n497) );
  XOR2_X1 U557 ( .A(KEYINPUT37), .B(n497), .Z(n522) );
  NOR2_X1 U558 ( .A1(n522), .A2(n498), .ZN(n501) );
  XOR2_X1 U559 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n499) );
  XNOR2_X1 U560 ( .A(KEYINPUT38), .B(n499), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(n508) );
  NAND2_X1 U562 ( .A1(n508), .A2(n557), .ZN(n504) );
  XNOR2_X1 U563 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n502), .B(KEYINPUT39), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n504), .B(n503), .ZN(G1328GAT) );
  NAND2_X1 U566 ( .A1(n525), .A2(n508), .ZN(n505) );
  XNOR2_X1 U567 ( .A(G36GAT), .B(n505), .ZN(G1329GAT) );
  NAND2_X1 U568 ( .A1(n539), .A2(n508), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n506), .B(KEYINPUT40), .ZN(n507) );
  XNOR2_X1 U570 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  NAND2_X1 U571 ( .A1(n508), .A2(n532), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n509), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n514) );
  INV_X1 U574 ( .A(n510), .ZN(n573) );
  NAND2_X1 U575 ( .A1(n573), .A2(n579), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n511), .B(KEYINPUT106), .ZN(n521) );
  NOR2_X1 U577 ( .A1(n521), .A2(n512), .ZN(n518) );
  NAND2_X1 U578 ( .A1(n557), .A2(n518), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(G1332GAT) );
  XOR2_X1 U580 ( .A(G64GAT), .B(KEYINPUT107), .Z(n516) );
  NAND2_X1 U581 ( .A1(n518), .A2(n525), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(G1333GAT) );
  NAND2_X1 U583 ( .A1(n539), .A2(n518), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n517), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U585 ( .A(G78GAT), .B(KEYINPUT43), .Z(n520) );
  NAND2_X1 U586 ( .A1(n518), .A2(n532), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  NOR2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n523), .B(KEYINPUT108), .ZN(n531) );
  NAND2_X1 U590 ( .A1(n531), .A2(n557), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n524), .B(G85GAT), .ZN(G1336GAT) );
  XOR2_X1 U592 ( .A(G92GAT), .B(KEYINPUT109), .Z(n527) );
  NAND2_X1 U593 ( .A1(n525), .A2(n531), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n527), .B(n526), .ZN(G1337GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n529) );
  NAND2_X1 U596 ( .A1(n531), .A2(n539), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U598 ( .A(G99GAT), .B(n530), .ZN(G1338GAT) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n536) );
  XOR2_X1 U600 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n534) );
  NAND2_X1 U601 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U602 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(G1339GAT) );
  NOR2_X1 U604 ( .A1(n555), .A2(n537), .ZN(n538) );
  NAND2_X1 U605 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n540), .B(KEYINPUT115), .ZN(n551) );
  NAND2_X1 U607 ( .A1(n551), .A2(n568), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n541), .B(KEYINPUT116), .ZN(n542) );
  XNOR2_X1 U609 ( .A(G113GAT), .B(n542), .ZN(G1340GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n544) );
  NAND2_X1 U611 ( .A1(n551), .A2(n573), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U613 ( .A(G120GAT), .B(n545), .Z(G1341GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n548) );
  NAND2_X1 U615 ( .A1(n551), .A2(n546), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U617 ( .A(G127GAT), .B(n549), .Z(G1342GAT) );
  XOR2_X1 U618 ( .A(G134GAT), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U619 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  NOR2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n565) );
  NOR2_X1 U623 ( .A1(n579), .A2(n565), .ZN(n558) );
  XOR2_X1 U624 ( .A(G141GAT), .B(n558), .Z(G1344GAT) );
  NOR2_X1 U625 ( .A1(n510), .A2(n565), .ZN(n563) );
  XOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n560) );
  XNOR2_X1 U627 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(KEYINPUT119), .B(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  NOR2_X1 U631 ( .A1(n588), .A2(n565), .ZN(n564) );
  XOR2_X1 U632 ( .A(G155GAT), .B(n564), .Z(G1346GAT) );
  NOR2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U634 ( .A(G162GAT), .B(n567), .Z(G1347GAT) );
  NAND2_X1 U635 ( .A1(n574), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n571) );
  XNOR2_X1 U638 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n570) );
  XNOR2_X1 U639 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U640 ( .A(KEYINPUT56), .B(n572), .Z(n576) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(G1349GAT) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n590) );
  NOR2_X1 U644 ( .A1(n590), .A2(n579), .ZN(n583) );
  XOR2_X1 U645 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n581) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n590), .ZN(n586) );
  XNOR2_X1 U650 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(G204GAT), .B(n587), .ZN(G1353GAT) );
  NOR2_X1 U653 ( .A1(n588), .A2(n590), .ZN(n589) );
  XOR2_X1 U654 ( .A(G211GAT), .B(n589), .Z(G1354GAT) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n593) );
  XNOR2_X1 U656 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

