

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738;

  XNOR2_X1 U378 ( .A(n410), .B(n446), .ZN(n611) );
  INV_X1 U379 ( .A(G953), .ZN(n715) );
  NOR2_X2 U380 ( .A1(n551), .A2(n664), .ZN(n412) );
  NOR2_X1 U381 ( .A1(n611), .A2(n723), .ZN(n655) );
  OR2_X2 U382 ( .A1(n669), .A2(n539), .ZN(n377) );
  XNOR2_X2 U383 ( .A(n534), .B(n465), .ZN(n487) );
  XNOR2_X2 U384 ( .A(n466), .B(G143), .ZN(n534) );
  NOR2_X1 U385 ( .A1(n667), .A2(n447), .ZN(n460) );
  XNOR2_X1 U386 ( .A(n433), .B(n432), .ZN(n667) );
  NOR2_X2 U387 ( .A1(n672), .A2(n673), .ZN(n434) );
  INV_X1 U388 ( .A(n559), .ZN(n596) );
  XOR2_X1 U389 ( .A(G119), .B(KEYINPUT3), .Z(n488) );
  AND2_X1 U390 ( .A1(n558), .A2(n628), .ZN(n442) );
  NAND2_X1 U391 ( .A1(n738), .A2(n635), .ZN(n554) );
  NAND2_X1 U392 ( .A1(n386), .A2(n384), .ZN(n648) );
  XNOR2_X1 U393 ( .A(n541), .B(n394), .ZN(n393) );
  NOR2_X1 U394 ( .A1(n567), .A2(n566), .ZN(n571) );
  NAND2_X1 U395 ( .A1(n588), .A2(n374), .ZN(n597) );
  NOR2_X1 U396 ( .A1(n663), .A2(n662), .ZN(n603) );
  XNOR2_X1 U397 ( .A(n378), .B(n508), .ZN(n669) );
  XNOR2_X1 U398 ( .A(n488), .B(G146), .ZN(n489) );
  XNOR2_X1 U399 ( .A(G902), .B(KEYINPUT15), .ZN(n493) );
  NOR2_X1 U400 ( .A1(n735), .A2(n734), .ZN(n370) );
  NOR2_X1 U401 ( .A1(n654), .A2(n444), .ZN(n443) );
  INV_X1 U402 ( .A(n737), .ZN(n444) );
  XNOR2_X1 U403 ( .A(n424), .B(n422), .ZN(n697) );
  XNOR2_X1 U404 ( .A(n423), .B(n517), .ZN(n422) );
  XNOR2_X1 U405 ( .A(n524), .B(n521), .ZN(n424) );
  XNOR2_X1 U406 ( .A(n523), .B(n518), .ZN(n423) );
  XNOR2_X1 U407 ( .A(n486), .B(G137), .ZN(n464) );
  XNOR2_X1 U408 ( .A(G134), .B(G131), .ZN(n486) );
  NAND2_X1 U409 ( .A1(n356), .A2(n419), .ZN(n368) );
  XNOR2_X1 U410 ( .A(n390), .B(KEYINPUT97), .ZN(n551) );
  NAND2_X1 U411 ( .A1(n648), .A2(n631), .ZN(n390) );
  XNOR2_X1 U412 ( .A(n379), .B(G125), .ZN(n497) );
  INV_X1 U413 ( .A(G146), .ZN(n379) );
  INV_X1 U414 ( .A(G128), .ZN(n466) );
  XNOR2_X1 U415 ( .A(n420), .B(G107), .ZN(n533) );
  XNOR2_X1 U416 ( .A(G116), .B(G122), .ZN(n420) );
  XOR2_X1 U417 ( .A(G113), .B(G104), .Z(n517) );
  NAND2_X1 U418 ( .A1(G234), .A2(G237), .ZN(n477) );
  XOR2_X1 U419 ( .A(KEYINPUT92), .B(KEYINPUT14), .Z(n478) );
  NAND2_X1 U420 ( .A1(n660), .A2(n659), .ZN(n663) );
  XNOR2_X1 U421 ( .A(n575), .B(KEYINPUT1), .ZN(n673) );
  XNOR2_X1 U422 ( .A(n471), .B(KEYINPUT90), .ZN(n472) );
  XNOR2_X1 U423 ( .A(n371), .B(n721), .ZN(n622) );
  XNOR2_X1 U424 ( .A(n372), .B(n358), .ZN(n371) );
  XNOR2_X1 U425 ( .A(n489), .B(n373), .ZN(n372) );
  XNOR2_X1 U426 ( .A(n498), .B(n382), .ZN(n381) );
  XNOR2_X1 U427 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n382) );
  XNOR2_X1 U428 ( .A(n499), .B(KEYINPUT70), .ZN(n439) );
  XNOR2_X1 U429 ( .A(G128), .B(G119), .ZN(n499) );
  XNOR2_X1 U430 ( .A(n497), .B(n437), .ZN(n722) );
  XNOR2_X1 U431 ( .A(n438), .B(G140), .ZN(n437) );
  INV_X1 U432 ( .A(KEYINPUT10), .ZN(n438) );
  XNOR2_X1 U433 ( .A(n414), .B(n501), .ZN(n527) );
  XNOR2_X1 U434 ( .A(n500), .B(n415), .ZN(n414) );
  INV_X1 U435 ( .A(KEYINPUT68), .ZN(n415) );
  XNOR2_X1 U436 ( .A(G134), .B(KEYINPUT9), .ZN(n528) );
  XOR2_X1 U437 ( .A(KEYINPUT100), .B(KEYINPUT7), .Z(n529) );
  AND2_X2 U438 ( .A1(n435), .A2(n440), .ZN(n699) );
  NOR2_X1 U439 ( .A1(n615), .A2(n493), .ZN(n435) );
  INV_X1 U440 ( .A(KEYINPUT33), .ZN(n432) );
  AND2_X1 U441 ( .A1(n571), .A2(n568), .ZN(n428) );
  NOR2_X1 U442 ( .A1(n597), .A2(n602), .ZN(n598) );
  INV_X1 U443 ( .A(KEYINPUT22), .ZN(n394) );
  NAND2_X1 U444 ( .A1(n601), .A2(n403), .ZN(n402) );
  XNOR2_X1 U445 ( .A(n525), .B(n430), .ZN(n547) );
  XNOR2_X1 U446 ( .A(n526), .B(n431), .ZN(n430) );
  INV_X1 U447 ( .A(G475), .ZN(n431) );
  XNOR2_X1 U448 ( .A(n507), .B(n506), .ZN(n508) );
  NOR2_X1 U449 ( .A1(n705), .A2(G902), .ZN(n378) );
  INV_X1 U450 ( .A(KEYINPUT94), .ZN(n506) );
  AND2_X1 U451 ( .A1(n393), .A2(n406), .ZN(n557) );
  XNOR2_X1 U452 ( .A(n512), .B(n407), .ZN(n515) );
  XNOR2_X1 U453 ( .A(n511), .B(n408), .ZN(n407) );
  NAND2_X1 U454 ( .A1(n699), .A2(G469), .ZN(n463) );
  NOR2_X1 U455 ( .A1(G953), .A2(G237), .ZN(n522) );
  OR2_X1 U456 ( .A1(G237), .A2(G902), .ZN(n474) );
  XNOR2_X1 U457 ( .A(n467), .B(G116), .ZN(n373) );
  XNOR2_X1 U458 ( .A(KEYINPUT5), .B(G113), .ZN(n467) );
  XNOR2_X1 U459 ( .A(G143), .B(G131), .ZN(n518) );
  XNOR2_X1 U460 ( .A(G122), .B(KEYINPUT12), .ZN(n519) );
  XOR2_X1 U461 ( .A(KEYINPUT98), .B(KEYINPUT11), .Z(n520) );
  XNOR2_X1 U462 ( .A(n413), .B(G101), .ZN(n490) );
  INV_X1 U463 ( .A(KEYINPUT65), .ZN(n413) );
  XNOR2_X1 U464 ( .A(n723), .B(n612), .ZN(n613) );
  INV_X1 U465 ( .A(KEYINPUT75), .ZN(n612) );
  INV_X1 U466 ( .A(KEYINPUT4), .ZN(n465) );
  XNOR2_X1 U467 ( .A(KEYINPUT78), .B(KEYINPUT17), .ZN(n454) );
  XNOR2_X1 U468 ( .A(KEYINPUT18), .B(KEYINPUT79), .ZN(n455) );
  XNOR2_X1 U469 ( .A(n497), .B(n468), .ZN(n396) );
  XNOR2_X1 U470 ( .A(n434), .B(KEYINPUT74), .ZN(n549) );
  INV_X1 U471 ( .A(n547), .ZN(n421) );
  XNOR2_X1 U472 ( .A(n596), .B(n595), .ZN(n660) );
  NOR2_X1 U473 ( .A1(n565), .A2(n564), .ZN(n576) );
  INV_X1 U474 ( .A(n539), .ZN(n403) );
  AND2_X1 U475 ( .A1(n676), .A2(n576), .ZN(n577) );
  INV_X1 U476 ( .A(KEYINPUT45), .ZN(n446) );
  AND2_X1 U477 ( .A1(n442), .A2(n552), .ZN(n441) );
  XNOR2_X1 U478 ( .A(n470), .B(n399), .ZN(n713) );
  XNOR2_X1 U479 ( .A(n533), .B(n469), .ZN(n399) );
  INV_X1 U480 ( .A(KEYINPUT16), .ZN(n469) );
  INV_X1 U481 ( .A(G107), .ZN(n509) );
  INV_X1 U482 ( .A(G104), .ZN(n408) );
  XNOR2_X1 U483 ( .A(G146), .B(G140), .ZN(n513) );
  XNOR2_X1 U484 ( .A(n490), .B(n397), .ZN(n512) );
  XNOR2_X1 U485 ( .A(G110), .B(KEYINPUT71), .ZN(n397) );
  XNOR2_X1 U486 ( .A(n365), .B(n713), .ZN(n616) );
  XNOR2_X1 U487 ( .A(n395), .B(n398), .ZN(n365) );
  XNOR2_X1 U488 ( .A(n512), .B(n396), .ZN(n395) );
  XNOR2_X1 U489 ( .A(n487), .B(n359), .ZN(n398) );
  XNOR2_X1 U490 ( .A(n405), .B(n404), .ZN(n689) );
  INV_X1 U491 ( .A(KEYINPUT93), .ZN(n404) );
  INV_X1 U492 ( .A(KEYINPUT31), .ZN(n389) );
  NAND2_X1 U493 ( .A1(n447), .A2(n389), .ZN(n387) );
  AND2_X1 U494 ( .A1(n376), .A2(n375), .ZN(n374) );
  XNOR2_X1 U495 ( .A(n585), .B(n586), .ZN(n376) );
  XNOR2_X1 U496 ( .A(KEYINPUT19), .B(KEYINPUT64), .ZN(n476) );
  XNOR2_X1 U497 ( .A(n623), .B(KEYINPUT62), .ZN(n624) );
  XNOR2_X1 U498 ( .A(n502), .B(n436), .ZN(n705) );
  XNOR2_X1 U499 ( .A(n380), .B(n722), .ZN(n436) );
  XNOR2_X1 U500 ( .A(n439), .B(n381), .ZN(n380) );
  BUF_X1 U501 ( .A(n699), .Z(n700) );
  XNOR2_X1 U502 ( .A(n532), .B(n417), .ZN(n698) );
  XNOR2_X1 U503 ( .A(n535), .B(n418), .ZN(n417) );
  INV_X1 U504 ( .A(KEYINPUT101), .ZN(n418) );
  AND2_X1 U505 ( .A1(n426), .A2(n425), .ZN(n654) );
  XNOR2_X1 U506 ( .A(n428), .B(n427), .ZN(n426) );
  XNOR2_X1 U507 ( .A(KEYINPUT105), .B(KEYINPUT43), .ZN(n427) );
  OR2_X1 U508 ( .A1(n604), .A2(n683), .ZN(n605) );
  NOR2_X1 U509 ( .A1(n406), .A2(n574), .ZN(n651) );
  INV_X1 U510 ( .A(KEYINPUT35), .ZN(n456) );
  AND2_X1 U511 ( .A1(n542), .A2(n409), .ZN(n392) );
  NAND2_X1 U512 ( .A1(n385), .A2(n383), .ZN(n384) );
  AND2_X1 U513 ( .A1(n388), .A2(n387), .ZN(n386) );
  NOR2_X1 U514 ( .A1(n447), .A2(n389), .ZN(n385) );
  XNOR2_X1 U515 ( .A(n599), .B(n429), .ZN(n642) );
  INV_X1 U516 ( .A(KEYINPUT104), .ZN(n429) );
  NAND2_X1 U517 ( .A1(n557), .A2(n543), .ZN(n635) );
  INV_X1 U518 ( .A(KEYINPUT60), .ZN(n449) );
  NAND2_X1 U519 ( .A1(n452), .A2(n451), .ZN(n450) );
  NAND2_X1 U520 ( .A1(n462), .A2(n451), .ZN(n461) );
  XNOR2_X1 U521 ( .A(n463), .B(n361), .ZN(n462) );
  NOR2_X1 U522 ( .A1(n692), .A2(G953), .ZN(n693) );
  AND2_X1 U523 ( .A1(n691), .A2(n360), .ZN(n400) );
  INV_X1 U524 ( .A(n406), .ZN(n409) );
  OR2_X1 U525 ( .A1(KEYINPUT47), .A2(n593), .ZN(n356) );
  XOR2_X1 U526 ( .A(n658), .B(KEYINPUT83), .Z(n357) );
  XOR2_X1 U527 ( .A(n490), .B(n491), .Z(n358) );
  XOR2_X1 U528 ( .A(n455), .B(n454), .Z(n359) );
  BUF_X1 U529 ( .A(n673), .Z(n406) );
  OR2_X1 U530 ( .A1(n667), .A2(n683), .ZN(n360) );
  XOR2_X1 U531 ( .A(n695), .B(n694), .Z(n361) );
  XOR2_X1 U532 ( .A(n697), .B(n696), .Z(n362) );
  XOR2_X1 U533 ( .A(n618), .B(n617), .Z(n363) );
  XNOR2_X1 U534 ( .A(n607), .B(KEYINPUT48), .ZN(n364) );
  NOR2_X1 U535 ( .A1(G952), .A2(n715), .ZN(n707) );
  INV_X1 U536 ( .A(n707), .ZN(n451) );
  NAND2_X1 U537 ( .A1(n553), .A2(n441), .ZN(n410) );
  XNOR2_X1 U538 ( .A(n366), .B(n364), .ZN(n445) );
  NAND2_X1 U539 ( .A1(n369), .A2(n367), .ZN(n366) );
  NOR2_X1 U540 ( .A1(n594), .A2(n368), .ZN(n367) );
  XNOR2_X1 U541 ( .A(n370), .B(KEYINPUT46), .ZN(n369) );
  XNOR2_X2 U542 ( .A(n487), .B(n464), .ZN(n721) );
  INV_X1 U543 ( .A(n587), .ZN(n375) );
  XNOR2_X2 U544 ( .A(n377), .B(KEYINPUT66), .ZN(n672) );
  INV_X1 U545 ( .A(n681), .ZN(n383) );
  NAND2_X1 U546 ( .A1(n681), .A2(n389), .ZN(n388) );
  XNOR2_X2 U547 ( .A(n391), .B(KEYINPUT32), .ZN(n738) );
  NAND2_X1 U548 ( .A1(n393), .A2(n392), .ZN(n391) );
  XNOR2_X1 U549 ( .A(n625), .B(n624), .ZN(n626) );
  NAND2_X1 U550 ( .A1(n699), .A2(G472), .ZN(n625) );
  NOR2_X2 U551 ( .A1(n620), .A2(n707), .ZN(n411) );
  NAND2_X1 U552 ( .A1(n357), .A2(n400), .ZN(n692) );
  NOR2_X2 U553 ( .A1(n626), .A2(n707), .ZN(n416) );
  OR2_X2 U554 ( .A1(n447), .A2(n402), .ZN(n541) );
  XNOR2_X1 U555 ( .A(n554), .B(n544), .ZN(n448) );
  NAND2_X1 U556 ( .A1(n554), .A2(KEYINPUT44), .ZN(n558) );
  NAND2_X1 U557 ( .A1(n401), .A2(n545), .ZN(n553) );
  NAND2_X1 U558 ( .A1(n448), .A2(n733), .ZN(n401) );
  XNOR2_X1 U559 ( .A(n453), .B(n362), .ZN(n452) );
  NOR2_X1 U560 ( .A1(n604), .A2(n581), .ZN(n641) );
  NAND2_X1 U561 ( .A1(n480), .A2(G952), .ZN(n405) );
  XNOR2_X2 U562 ( .A(n485), .B(n484), .ZN(n447) );
  XNOR2_X1 U563 ( .A(n411), .B(n621), .ZN(G51) );
  XNOR2_X1 U564 ( .A(n412), .B(KEYINPUT103), .ZN(n552) );
  XNOR2_X1 U565 ( .A(n416), .B(n627), .ZN(G57) );
  INV_X1 U566 ( .A(n651), .ZN(n419) );
  INV_X1 U567 ( .A(n548), .ZN(n540) );
  INV_X1 U568 ( .A(n662), .ZN(n601) );
  INV_X1 U569 ( .A(n660), .ZN(n602) );
  NAND2_X1 U570 ( .A1(n548), .A2(n421), .ZN(n662) );
  INV_X1 U571 ( .A(n596), .ZN(n425) );
  NAND2_X1 U572 ( .A1(n548), .A2(n547), .ZN(n599) );
  NAND2_X1 U573 ( .A1(n549), .A2(n555), .ZN(n433) );
  XNOR2_X2 U574 ( .A(n610), .B(KEYINPUT76), .ZN(n440) );
  NAND2_X1 U575 ( .A1(n657), .A2(n440), .ZN(n658) );
  NAND2_X1 U576 ( .A1(n445), .A2(n443), .ZN(n723) );
  NOR2_X1 U577 ( .A1(n447), .A2(n676), .ZN(n550) );
  XNOR2_X1 U578 ( .A(n450), .B(n449), .ZN(G60) );
  NAND2_X1 U579 ( .A1(n699), .A2(G475), .ZN(n453) );
  XNOR2_X2 U580 ( .A(n457), .B(n456), .ZN(n733) );
  NAND2_X1 U581 ( .A1(n459), .A2(n458), .ZN(n457) );
  INV_X1 U582 ( .A(n589), .ZN(n458) );
  XNOR2_X1 U583 ( .A(n460), .B(KEYINPUT34), .ZN(n459) );
  XNOR2_X1 U584 ( .A(n461), .B(KEYINPUT119), .ZN(G54) );
  XNOR2_X1 U585 ( .A(n619), .B(n363), .ZN(n620) );
  NOR2_X2 U586 ( .A1(n559), .A2(n584), .ZN(n570) );
  INV_X1 U587 ( .A(KEYINPUT85), .ZN(n544) );
  INV_X1 U588 ( .A(KEYINPUT84), .ZN(n607) );
  XNOR2_X1 U589 ( .A(n510), .B(n509), .ZN(n511) );
  NOR2_X1 U590 ( .A1(n655), .A2(KEYINPUT2), .ZN(n656) );
  INV_X1 U591 ( .A(KEYINPUT0), .ZN(n484) );
  INV_X1 U592 ( .A(n575), .ZN(n580) );
  XNOR2_X1 U593 ( .A(KEYINPUT87), .B(KEYINPUT63), .ZN(n627) );
  NAND2_X1 U594 ( .A1(G224), .A2(n715), .ZN(n468) );
  XNOR2_X1 U595 ( .A(n488), .B(n517), .ZN(n470) );
  NAND2_X1 U596 ( .A1(n616), .A2(n493), .ZN(n473) );
  NAND2_X1 U597 ( .A1(n474), .A2(G210), .ZN(n471) );
  XNOR2_X2 U598 ( .A(n473), .B(n472), .ZN(n559) );
  NAND2_X1 U599 ( .A1(G214), .A2(n474), .ZN(n475) );
  XNOR2_X1 U600 ( .A(KEYINPUT91), .B(n475), .ZN(n584) );
  XNOR2_X1 U601 ( .A(n570), .B(n476), .ZN(n581) );
  XNOR2_X1 U602 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U603 ( .A(KEYINPUT72), .B(n479), .Z(n480) );
  NOR2_X1 U604 ( .A1(G953), .A2(n689), .ZN(n562) );
  AND2_X1 U605 ( .A1(G953), .A2(n480), .ZN(n481) );
  NAND2_X1 U606 ( .A1(G902), .A2(n481), .ZN(n560) );
  NOR2_X1 U607 ( .A1(n560), .A2(G898), .ZN(n482) );
  NOR2_X1 U608 ( .A1(n562), .A2(n482), .ZN(n483) );
  NOR2_X1 U609 ( .A1(n581), .A2(n483), .ZN(n485) );
  NAND2_X1 U610 ( .A1(n522), .A2(G210), .ZN(n491) );
  NOR2_X1 U611 ( .A1(n622), .A2(G902), .ZN(n492) );
  XNOR2_X1 U612 ( .A(G472), .B(n492), .ZN(n583) );
  INV_X1 U613 ( .A(n583), .ZN(n676) );
  XNOR2_X1 U614 ( .A(n676), .B(KEYINPUT6), .ZN(n567) );
  INV_X1 U615 ( .A(n567), .ZN(n555) );
  XOR2_X1 U616 ( .A(KEYINPUT95), .B(KEYINPUT21), .Z(n496) );
  NAND2_X1 U617 ( .A1(G234), .A2(n493), .ZN(n494) );
  XNOR2_X1 U618 ( .A(KEYINPUT20), .B(n494), .ZN(n503) );
  NAND2_X1 U619 ( .A1(n503), .A2(G221), .ZN(n495) );
  XNOR2_X1 U620 ( .A(n496), .B(n495), .ZN(n670) );
  XNOR2_X1 U621 ( .A(KEYINPUT96), .B(n670), .ZN(n539) );
  XNOR2_X1 U622 ( .A(G137), .B(G110), .ZN(n498) );
  XOR2_X1 U623 ( .A(KEYINPUT8), .B(KEYINPUT67), .Z(n501) );
  NAND2_X1 U624 ( .A1(G234), .A2(n715), .ZN(n500) );
  NAND2_X1 U625 ( .A1(G221), .A2(n527), .ZN(n502) );
  XOR2_X1 U626 ( .A(KEYINPUT77), .B(KEYINPUT25), .Z(n505) );
  NAND2_X1 U627 ( .A1(n503), .A2(G217), .ZN(n504) );
  XNOR2_X1 U628 ( .A(n505), .B(n504), .ZN(n507) );
  NAND2_X1 U629 ( .A1(G227), .A2(n715), .ZN(n510) );
  XNOR2_X1 U630 ( .A(n721), .B(n513), .ZN(n514) );
  XNOR2_X1 U631 ( .A(n515), .B(n514), .ZN(n695) );
  NOR2_X1 U632 ( .A1(n695), .A2(G902), .ZN(n516) );
  XNOR2_X2 U633 ( .A(n516), .B(G469), .ZN(n575) );
  XNOR2_X1 U634 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n526) );
  XNOR2_X1 U635 ( .A(n520), .B(n519), .ZN(n521) );
  NAND2_X1 U636 ( .A1(G214), .A2(n522), .ZN(n523) );
  INV_X1 U637 ( .A(n722), .ZN(n524) );
  NOR2_X1 U638 ( .A1(G902), .A2(n697), .ZN(n525) );
  NAND2_X1 U639 ( .A1(G217), .A2(n527), .ZN(n531) );
  XNOR2_X1 U640 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U641 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U642 ( .A(n533), .B(n534), .ZN(n535) );
  NOR2_X1 U643 ( .A1(G902), .A2(n698), .ZN(n536) );
  XNOR2_X1 U644 ( .A(G478), .B(n536), .ZN(n548) );
  NAND2_X1 U645 ( .A1(n547), .A2(n540), .ZN(n589) );
  INV_X1 U646 ( .A(KEYINPUT44), .ZN(n537) );
  XNOR2_X1 U647 ( .A(n733), .B(n537), .ZN(n545) );
  INV_X1 U648 ( .A(n669), .ZN(n565) );
  XOR2_X1 U649 ( .A(KEYINPUT80), .B(n567), .Z(n538) );
  NOR2_X1 U650 ( .A1(n565), .A2(n538), .ZN(n542) );
  NOR2_X1 U651 ( .A1(n565), .A2(n676), .ZN(n543) );
  OR2_X1 U652 ( .A1(n547), .A2(n548), .ZN(n546) );
  XOR2_X1 U653 ( .A(n546), .B(KEYINPUT102), .Z(n636) );
  INV_X1 U654 ( .A(n636), .ZN(n649) );
  NAND2_X1 U655 ( .A1(n649), .A2(n599), .ZN(n582) );
  INV_X1 U656 ( .A(n582), .ZN(n664) );
  NAND2_X1 U657 ( .A1(n676), .A2(n549), .ZN(n681) );
  NOR2_X1 U658 ( .A1(n672), .A2(n575), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n588), .A2(n550), .ZN(n631) );
  NOR2_X1 U660 ( .A1(n555), .A2(n669), .ZN(n556) );
  NAND2_X1 U661 ( .A1(n557), .A2(n556), .ZN(n628) );
  NOR2_X1 U662 ( .A1(G900), .A2(n560), .ZN(n561) );
  NOR2_X1 U663 ( .A1(n562), .A2(n561), .ZN(n587) );
  NOR2_X1 U664 ( .A1(n670), .A2(n587), .ZN(n563) );
  XNOR2_X1 U665 ( .A(n563), .B(KEYINPUT69), .ZN(n564) );
  NAND2_X1 U666 ( .A1(n576), .A2(n642), .ZN(n566) );
  NOR2_X1 U667 ( .A1(n409), .A2(n584), .ZN(n568) );
  XNOR2_X1 U668 ( .A(KEYINPUT36), .B(KEYINPUT86), .ZN(n569) );
  XNOR2_X1 U669 ( .A(n569), .B(KEYINPUT109), .ZN(n573) );
  NAND2_X1 U670 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U671 ( .A(n573), .B(n572), .Z(n574) );
  XNOR2_X1 U672 ( .A(KEYINPUT28), .B(KEYINPUT107), .ZN(n578) );
  XOR2_X1 U673 ( .A(n578), .B(n577), .Z(n579) );
  NAND2_X1 U674 ( .A1(n580), .A2(n579), .ZN(n604) );
  NAND2_X1 U675 ( .A1(n641), .A2(n582), .ZN(n593) );
  NAND2_X1 U676 ( .A1(n593), .A2(KEYINPUT47), .ZN(n591) );
  XOR2_X1 U677 ( .A(KEYINPUT30), .B(KEYINPUT106), .Z(n586) );
  INV_X1 U678 ( .A(n584), .ZN(n659) );
  NAND2_X1 U679 ( .A1(n676), .A2(n659), .ZN(n585) );
  NOR2_X1 U680 ( .A1(n597), .A2(n589), .ZN(n590) );
  NAND2_X1 U681 ( .A1(n590), .A2(n596), .ZN(n639) );
  NAND2_X1 U682 ( .A1(n591), .A2(n639), .ZN(n592) );
  XNOR2_X1 U683 ( .A(n592), .B(KEYINPUT82), .ZN(n594) );
  XNOR2_X1 U684 ( .A(KEYINPUT38), .B(KEYINPUT73), .ZN(n595) );
  XNOR2_X1 U685 ( .A(KEYINPUT39), .B(n598), .ZN(n608) );
  NOR2_X1 U686 ( .A1(n599), .A2(n608), .ZN(n600) );
  XNOR2_X1 U687 ( .A(n600), .B(KEYINPUT40), .ZN(n735) );
  XOR2_X1 U688 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n606) );
  XNOR2_X1 U689 ( .A(KEYINPUT41), .B(n603), .ZN(n683) );
  XNOR2_X1 U690 ( .A(n606), .B(n605), .ZN(n734) );
  NOR2_X1 U691 ( .A1(n608), .A2(n649), .ZN(n609) );
  XOR2_X1 U692 ( .A(KEYINPUT110), .B(n609), .Z(n737) );
  NAND2_X1 U693 ( .A1(n655), .A2(KEYINPUT2), .ZN(n610) );
  NOR2_X1 U694 ( .A1(n611), .A2(n613), .ZN(n614) );
  NOR2_X1 U695 ( .A1(KEYINPUT2), .A2(n614), .ZN(n615) );
  NAND2_X1 U696 ( .A1(n699), .A2(G210), .ZN(n619) );
  XOR2_X1 U697 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n618) );
  XNOR2_X1 U698 ( .A(n616), .B(KEYINPUT88), .ZN(n617) );
  XNOR2_X1 U699 ( .A(KEYINPUT56), .B(KEYINPUT118), .ZN(n621) );
  XOR2_X1 U700 ( .A(n622), .B(KEYINPUT89), .Z(n623) );
  XNOR2_X1 U701 ( .A(G101), .B(n628), .ZN(G3) );
  INV_X1 U702 ( .A(n642), .ZN(n644) );
  NOR2_X1 U703 ( .A1(n644), .A2(n631), .ZN(n630) );
  XNOR2_X1 U704 ( .A(G104), .B(KEYINPUT111), .ZN(n629) );
  XNOR2_X1 U705 ( .A(n630), .B(n629), .ZN(G6) );
  NOR2_X1 U706 ( .A1(n649), .A2(n631), .ZN(n633) );
  XNOR2_X1 U707 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n632) );
  XNOR2_X1 U708 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U709 ( .A(G107), .B(n634), .ZN(G9) );
  XNOR2_X1 U710 ( .A(G110), .B(n635), .ZN(G12) );
  XOR2_X1 U711 ( .A(G128), .B(KEYINPUT29), .Z(n638) );
  NAND2_X1 U712 ( .A1(n641), .A2(n636), .ZN(n637) );
  XNOR2_X1 U713 ( .A(n638), .B(n637), .ZN(G30) );
  XNOR2_X1 U714 ( .A(G143), .B(KEYINPUT112), .ZN(n640) );
  XNOR2_X1 U715 ( .A(n640), .B(n639), .ZN(G45) );
  NAND2_X1 U716 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U717 ( .A(n643), .B(G146), .ZN(G48) );
  NOR2_X1 U718 ( .A1(n644), .A2(n648), .ZN(n646) );
  XNOR2_X1 U719 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n645) );
  XNOR2_X1 U720 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U721 ( .A(G113), .B(n647), .ZN(G15) );
  NOR2_X1 U722 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U723 ( .A(G116), .B(n650), .Z(G18) );
  XOR2_X1 U724 ( .A(KEYINPUT115), .B(KEYINPUT37), .Z(n653) );
  XNOR2_X1 U725 ( .A(G125), .B(n651), .ZN(n652) );
  XNOR2_X1 U726 ( .A(n653), .B(n652), .ZN(G27) );
  XOR2_X1 U727 ( .A(G140), .B(n654), .Z(G42) );
  XNOR2_X1 U728 ( .A(KEYINPUT81), .B(n656), .ZN(n657) );
  NOR2_X1 U729 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U730 ( .A1(n662), .A2(n661), .ZN(n666) );
  NOR2_X1 U731 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U732 ( .A1(n666), .A2(n665), .ZN(n668) );
  NOR2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n686) );
  NAND2_X1 U734 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U735 ( .A(KEYINPUT49), .B(n671), .Z(n679) );
  XOR2_X1 U736 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n675) );
  NAND2_X1 U737 ( .A1(n406), .A2(n672), .ZN(n674) );
  XNOR2_X1 U738 ( .A(n675), .B(n674), .ZN(n677) );
  NOR2_X1 U739 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U740 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U741 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U742 ( .A(KEYINPUT51), .B(n682), .ZN(n684) );
  NOR2_X1 U743 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U744 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U745 ( .A(KEYINPUT52), .B(n687), .ZN(n688) );
  NOR2_X1 U746 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U747 ( .A(n690), .B(KEYINPUT117), .ZN(n691) );
  XNOR2_X1 U748 ( .A(n693), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U749 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n694) );
  XOR2_X1 U750 ( .A(KEYINPUT59), .B(KEYINPUT120), .Z(n696) );
  XOR2_X1 U751 ( .A(n698), .B(KEYINPUT121), .Z(n702) );
  NAND2_X1 U752 ( .A1(n700), .A2(G478), .ZN(n701) );
  XNOR2_X1 U753 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U754 ( .A1(n707), .A2(n703), .ZN(G63) );
  NAND2_X1 U755 ( .A1(G217), .A2(n700), .ZN(n704) );
  XNOR2_X1 U756 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U757 ( .A1(n707), .A2(n706), .ZN(G66) );
  OR2_X1 U758 ( .A1(G953), .A2(n611), .ZN(n712) );
  NAND2_X1 U759 ( .A1(G224), .A2(G953), .ZN(n708) );
  XNOR2_X1 U760 ( .A(n708), .B(KEYINPUT122), .ZN(n709) );
  XNOR2_X1 U761 ( .A(KEYINPUT61), .B(n709), .ZN(n710) );
  NAND2_X1 U762 ( .A1(n710), .A2(G898), .ZN(n711) );
  NAND2_X1 U763 ( .A1(n712), .A2(n711), .ZN(n719) );
  XOR2_X1 U764 ( .A(n713), .B(G101), .Z(n714) );
  XNOR2_X1 U765 ( .A(G110), .B(n714), .ZN(n717) );
  NOR2_X1 U766 ( .A1(G898), .A2(n715), .ZN(n716) );
  NOR2_X1 U767 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U768 ( .A(n719), .B(n718), .ZN(n720) );
  XOR2_X1 U769 ( .A(KEYINPUT123), .B(n720), .Z(G69) );
  XOR2_X1 U770 ( .A(n722), .B(n721), .Z(n727) );
  XOR2_X1 U771 ( .A(n723), .B(n727), .Z(n724) );
  XNOR2_X1 U772 ( .A(KEYINPUT124), .B(n724), .ZN(n725) );
  NOR2_X1 U773 ( .A1(G953), .A2(n725), .ZN(n726) );
  XNOR2_X1 U774 ( .A(KEYINPUT125), .B(n726), .ZN(n731) );
  XNOR2_X1 U775 ( .A(G227), .B(n727), .ZN(n728) );
  NAND2_X1 U776 ( .A1(n728), .A2(G900), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n729), .A2(G953), .ZN(n730) );
  NAND2_X1 U778 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U779 ( .A(n732), .B(KEYINPUT126), .ZN(G72) );
  XNOR2_X1 U780 ( .A(n733), .B(G122), .ZN(G24) );
  XOR2_X1 U781 ( .A(G137), .B(n734), .Z(G39) );
  XNOR2_X1 U782 ( .A(G131), .B(KEYINPUT127), .ZN(n736) );
  XNOR2_X1 U783 ( .A(n736), .B(n735), .ZN(G33) );
  XNOR2_X1 U784 ( .A(G134), .B(n737), .ZN(G36) );
  XNOR2_X1 U785 ( .A(n738), .B(G119), .ZN(G21) );
endmodule

