//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973;
  NAND2_X1  g000(.A1(G211gat), .A2(G218gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT22), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205));
  AND2_X1   g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT78), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n202), .ZN(new_n210));
  NOR2_X1   g009(.A1(G211gat), .A2(G218gat), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT77), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G211gat), .ZN(new_n213));
  INV_X1    g012(.A(G218gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT77), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(new_n216), .A3(new_n202), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n204), .B(KEYINPUT78), .C1(new_n205), .C2(new_n206), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n209), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n206), .ZN(new_n221));
  INV_X1    g020(.A(new_n205), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n221), .A2(new_n222), .B1(new_n203), .B2(new_n202), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n223), .A2(KEYINPUT78), .A3(new_n212), .A4(new_n217), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT79), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT79), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n220), .A2(new_n227), .A3(new_n224), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT29), .ZN(new_n229));
  XOR2_X1   g028(.A(G141gat), .B(G148gat), .Z(new_n230));
  INV_X1    g029(.A(G155gat), .ZN(new_n231));
  INV_X1    g030(.A(G162gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G155gat), .A2(G162gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(KEYINPUT2), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n230), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G141gat), .B(G148gat), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n234), .B(new_n233), .C1(new_n238), .C2(KEYINPUT2), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  AOI22_X1  g040(.A1(new_n226), .A2(new_n228), .B1(new_n229), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G228gat), .A2(G233gat), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n237), .A2(new_n239), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n220), .A2(new_n229), .A3(new_n224), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n244), .B1(new_n245), .B2(new_n240), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n242), .A2(new_n243), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n243), .ZN(new_n248));
  INV_X1    g047(.A(new_n228), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n227), .B1(new_n220), .B2(new_n224), .ZN(new_n250));
  INV_X1    g049(.A(new_n241), .ZN(new_n251));
  OAI22_X1  g050(.A1(new_n249), .A2(new_n250), .B1(KEYINPUT29), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n246), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n248), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n247), .A2(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(G78gat), .B(G106gat), .Z(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT87), .B(G50gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT86), .B(KEYINPUT31), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G22gat), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n260), .B1(new_n247), .B2(new_n254), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT88), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n243), .B1(new_n242), .B2(new_n246), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n252), .A2(new_n253), .A3(new_n248), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n261), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NOR3_X1   g068(.A1(new_n269), .A2(KEYINPUT88), .A3(G22gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n262), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n264), .A2(new_n265), .A3(new_n263), .ZN(new_n272));
  OAI21_X1  g071(.A(G22gat), .B1(new_n269), .B2(KEYINPUT88), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n272), .A2(new_n273), .A3(new_n255), .A4(new_n261), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G8gat), .B(G36gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(G64gat), .B(G92gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G226gat), .A2(G233gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT27), .B(G183gat), .ZN(new_n282));
  INV_X1    g081(.A(G190gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(KEYINPUT28), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT66), .B(G183gat), .ZN(new_n286));
  AOI21_X1  g085(.A(G190gat), .B1(new_n286), .B2(KEYINPUT27), .ZN(new_n287));
  AND2_X1   g086(.A1(KEYINPUT67), .A2(KEYINPUT27), .ZN(new_n288));
  NOR2_X1   g087(.A1(KEYINPUT67), .A2(KEYINPUT27), .ZN(new_n289));
  OAI21_X1  g088(.A(G183gat), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT68), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g091(.A(KEYINPUT68), .B(G183gat), .C1(new_n288), .C2(new_n289), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n287), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n285), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT26), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g101(.A(KEYINPUT70), .B(new_n297), .C1(new_n298), .C2(new_n299), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n298), .A2(new_n299), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  XOR2_X1   g106(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n308));
  INV_X1    g107(.A(G169gat), .ZN(new_n309));
  INV_X1    g108(.A(G176gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(new_n310), .A3(KEYINPUT23), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n312), .B1(G169gat), .B2(G176gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n313), .A3(new_n297), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT24), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n306), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G183gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(new_n283), .ZN(new_n318));
  NAND3_X1  g117(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n314), .B1(KEYINPUT65), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT65), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n316), .A2(new_n318), .A3(new_n322), .A4(new_n319), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n308), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n286), .A2(new_n283), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n316), .A2(new_n319), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT25), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n314), .A2(new_n328), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  OAI22_X1  g129(.A1(new_n296), .A2(new_n307), .B1(new_n324), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n281), .B1(new_n331), .B2(new_n229), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n294), .A2(new_n295), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n284), .ZN(new_n334));
  INV_X1    g133(.A(new_n307), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n320), .A2(KEYINPUT65), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n311), .A2(new_n313), .A3(new_n297), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n323), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n308), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n339), .A2(new_n340), .B1(new_n327), .B2(new_n329), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n280), .B1(new_n336), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n249), .A2(new_n250), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n332), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n344), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n341), .B1(new_n334), .B2(new_n335), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n280), .B1(new_n347), .B2(KEYINPUT29), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n281), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n346), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n279), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT37), .B1(new_n345), .B2(new_n350), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n348), .A2(new_n346), .A3(new_n349), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n344), .B1(new_n332), .B2(new_n343), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT37), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n279), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT38), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n351), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n355), .B1(new_n353), .B2(new_n354), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n278), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n362), .A2(KEYINPUT38), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n240), .B1(new_n237), .B2(new_n239), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n251), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G120gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(G113gat), .ZN(new_n368));
  INV_X1    g167(.A(G113gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G120gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G127gat), .B(G134gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT72), .B(KEYINPUT1), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT73), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n372), .A2(new_n371), .A3(new_n373), .A4(KEYINPUT73), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n371), .A2(KEYINPUT71), .ZN(new_n379));
  XNOR2_X1  g178(.A(G113gat), .B(G120gat), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT71), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT1), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n379), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n372), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n378), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n366), .A2(new_n387), .ZN(new_n388));
  AND2_X1   g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n389), .A2(KEYINPUT5), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n376), .A2(new_n377), .B1(new_n384), .B2(new_n385), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n391), .B1(new_n392), .B2(new_n244), .ZN(new_n393));
  AND4_X1   g192(.A1(new_n391), .A2(new_n378), .A3(new_n386), .A4(new_n244), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n388), .B(new_n390), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT83), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n378), .A2(new_n386), .A3(new_n244), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT4), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n378), .A2(new_n386), .A3(new_n244), .A4(new_n391), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n400), .A2(new_n401), .A3(new_n388), .A4(new_n390), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n396), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(KEYINPUT82), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT82), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n392), .A2(new_n405), .A3(new_n391), .A4(new_n244), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(new_n406), .A3(new_n398), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n389), .B1(new_n366), .B2(new_n387), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n244), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n387), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n397), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n389), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n409), .A2(KEYINPUT5), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n403), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G1gat), .B(G29gat), .ZN(new_n416));
  INV_X1    g215(.A(G85gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT0), .B(G57gat), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n418), .B(new_n419), .Z(new_n420));
  NAND2_X1  g219(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n420), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n403), .A2(new_n414), .A3(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT84), .B(KEYINPUT6), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n421), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n415), .A2(new_n420), .A3(new_n424), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT85), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n415), .A2(KEYINPUT85), .A3(new_n420), .A4(new_n424), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n426), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n275), .B1(new_n364), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT80), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n278), .B1(new_n353), .B2(new_n354), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT81), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n433), .B(KEYINPUT30), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n345), .A2(new_n350), .A3(new_n279), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT80), .B1(new_n351), .B2(KEYINPUT81), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT30), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n440), .B1(new_n351), .B2(KEYINPUT80), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n436), .B(new_n438), .C1(new_n439), .C2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n388), .B1(new_n393), .B2(new_n394), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n389), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n444), .B(KEYINPUT39), .C1(new_n389), .C2(new_n412), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT39), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n443), .A2(new_n446), .A3(new_n389), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n445), .A2(KEYINPUT40), .A3(new_n422), .A4(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT40), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT39), .B1(new_n412), .B2(new_n389), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n450), .B1(new_n389), .B2(new_n443), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n447), .A2(new_n422), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n421), .A2(new_n448), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n442), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT89), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT89), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n458), .A3(new_n455), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n432), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n426), .A2(new_n429), .A3(new_n430), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT30), .B1(new_n434), .B2(new_n433), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n437), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n461), .A2(new_n436), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT34), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT74), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n336), .A2(new_n467), .A3(new_n387), .A4(new_n342), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n392), .A2(KEYINPUT74), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n387), .A2(new_n467), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n331), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(G227gat), .ZN(new_n473));
  INV_X1    g272(.A(G233gat), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n466), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  AOI211_X1 g276(.A(KEYINPUT34), .B(new_n475), .C1(new_n468), .C2(new_n471), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n468), .A2(new_n471), .A3(new_n475), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT32), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT33), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(G15gat), .B(G43gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(G71gat), .B(G99gat), .ZN(new_n485));
  XOR2_X1   g284(.A(new_n484), .B(new_n485), .Z(new_n486));
  NAND3_X1  g285(.A1(new_n481), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n486), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n480), .B(KEYINPUT32), .C1(new_n482), .C2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n479), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT76), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n487), .A2(new_n489), .ZN(new_n493));
  INV_X1    g292(.A(new_n479), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n479), .A2(new_n487), .A3(KEYINPUT76), .A4(new_n489), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n492), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT75), .ZN(new_n500));
  INV_X1    g299(.A(new_n477), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n472), .A2(new_n466), .A3(new_n476), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n493), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n489), .B(new_n487), .C1(new_n479), .C2(new_n500), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT36), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n465), .A2(new_n275), .B1(new_n499), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n497), .A2(new_n275), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT35), .ZN(new_n509));
  INV_X1    g308(.A(new_n442), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n508), .A2(new_n509), .A3(new_n461), .A4(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n504), .A2(new_n271), .A3(new_n505), .A4(new_n274), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT35), .B1(new_n465), .B2(new_n512), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n460), .A2(new_n507), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT99), .ZN(new_n515));
  NAND2_X1  g314(.A1(G99gat), .A2(G106gat), .ZN(new_n516));
  INV_X1    g315(.A(G92gat), .ZN(new_n517));
  AOI22_X1  g316(.A1(KEYINPUT8), .A2(new_n516), .B1(new_n417), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G85gat), .A2(G92gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT7), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n518), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G99gat), .B(G106gat), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n515), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n525), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n521), .A2(new_n522), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n528), .A2(KEYINPUT99), .A3(new_n524), .A4(new_n518), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G43gat), .B(G50gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT15), .ZN(new_n534));
  OR2_X1    g333(.A1(KEYINPUT93), .A2(G43gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(KEYINPUT93), .A2(G43gat), .ZN(new_n536));
  AOI21_X1  g335(.A(G50gat), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT15), .ZN(new_n538));
  INV_X1    g337(.A(G43gat), .ZN(new_n539));
  INV_X1    g338(.A(G50gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n534), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(G29gat), .A2(G36gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT91), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT91), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(G29gat), .B2(G36gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(new_n546), .A3(KEYINPUT14), .ZN(new_n547));
  INV_X1    g346(.A(G36gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT92), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT92), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(G36gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n551), .A3(G29gat), .ZN(new_n552));
  OR3_X1    g351(.A1(new_n543), .A2(KEYINPUT91), .A3(KEYINPUT14), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n542), .A2(new_n547), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n547), .A2(new_n553), .A3(new_n552), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n534), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n532), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT41), .ZN(new_n559));
  NAND2_X1  g358(.A1(G232gat), .A2(G233gat), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G134gat), .B(G162gat), .Z(new_n562));
  NOR2_X1   g361(.A1(new_n532), .A2(new_n557), .ZN(new_n563));
  OR3_X1    g362(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(G190gat), .B(G218gat), .Z(new_n565));
  NAND2_X1  g364(.A1(new_n560), .A2(new_n559), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n562), .B1(new_n561), .B2(new_n563), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n567), .B1(new_n564), .B2(new_n568), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G15gat), .B(G22gat), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n573), .A2(G1gat), .ZN(new_n574));
  INV_X1    g373(.A(G1gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT16), .ZN(new_n576));
  INV_X1    g375(.A(G15gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(G22gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n263), .A2(G15gat), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(G8gat), .B1(new_n574), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n573), .A2(new_n576), .ZN(new_n582));
  INV_X1    g381(.A(G8gat), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n582), .B(new_n583), .C1(G1gat), .C2(new_n573), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT21), .ZN(new_n587));
  XNOR2_X1  g386(.A(G57gat), .B(G64gat), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  OR2_X1    g388(.A1(G71gat), .A2(G78gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT9), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n589), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n591), .B(new_n590), .C1(new_n588), .C2(new_n593), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n586), .B1(new_n587), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n595), .A2(new_n596), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT21), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n598), .B1(new_n600), .B2(new_n586), .ZN(new_n601));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT98), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(new_n317), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(G211gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n601), .B(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G127gat), .B(G155gat), .Z(new_n607));
  XOR2_X1   g406(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n606), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n572), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n514), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT94), .B1(new_n557), .B2(new_n586), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT94), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n554), .A2(new_n585), .A3(new_n614), .A4(new_n556), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n557), .A2(KEYINPUT17), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n554), .A2(new_n531), .A3(new_n556), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(new_n586), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G229gat), .A2(G233gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT18), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n621), .B1(KEYINPUT96), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n616), .A2(new_n619), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT96), .B1(new_n625), .B2(new_n622), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n557), .A2(new_n586), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n616), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n620), .B(KEYINPUT13), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n616), .A2(new_n619), .A3(new_n626), .A4(new_n623), .ZN(new_n634));
  XNOR2_X1  g433(.A(G113gat), .B(G141gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G197gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT11), .B(G169gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n638), .B(KEYINPUT12), .Z(new_n639));
  NAND4_X1  g438(.A1(new_n628), .A2(new_n633), .A3(new_n634), .A4(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT97), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI22_X1  g441(.A1(new_n624), .A2(new_n627), .B1(new_n630), .B2(new_n632), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n643), .A2(KEYINPUT97), .A3(new_n634), .A4(new_n639), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n634), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n639), .B(KEYINPUT90), .ZN(new_n646));
  AOI22_X1  g445(.A1(new_n642), .A2(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n648));
  NAND2_X1  g447(.A1(G230gat), .A2(G233gat), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT10), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n525), .B1(new_n523), .B2(KEYINPUT100), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n523), .A2(KEYINPUT100), .A3(new_n525), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n653), .A2(new_n599), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT101), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n597), .A2(new_n652), .ZN(new_n658));
  AOI22_X1  g457(.A1(new_n654), .A2(new_n658), .B1(new_n530), .B2(new_n597), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n651), .B(new_n657), .C1(new_n659), .C2(new_n656), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n530), .A2(new_n651), .A3(new_n597), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n650), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n530), .A2(new_n597), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n656), .B1(new_n664), .B2(new_n655), .ZN(new_n665));
  AOI21_X1  g464(.A(KEYINPUT101), .B1(new_n658), .B2(new_n654), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(new_n649), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n648), .B1(new_n663), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(G176gat), .B(G204gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT102), .ZN(new_n671));
  XNOR2_X1  g470(.A(G120gat), .B(G148gat), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n671), .B(new_n672), .Z(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n648), .B(new_n673), .C1(new_n663), .C2(new_n668), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n647), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n612), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(new_n461), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(new_n575), .ZN(G1324gat));
  INV_X1    g480(.A(new_n679), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n442), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT16), .B(G8gat), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OR3_X1    g484(.A1(new_n685), .A2(KEYINPUT104), .A3(KEYINPUT42), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT104), .B1(new_n685), .B2(KEYINPUT42), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n683), .A2(G8gat), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n685), .A2(KEYINPUT42), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n686), .A2(new_n687), .A3(new_n688), .A4(new_n689), .ZN(G1325gat));
  NAND2_X1  g489(.A1(new_n499), .A2(new_n506), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n679), .A2(new_n577), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n497), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n682), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n692), .B1(new_n577), .B2(new_n694), .ZN(G1326gat));
  INV_X1    g494(.A(new_n275), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n679), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT43), .B(G22gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  INV_X1    g498(.A(new_n610), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n678), .A2(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n514), .A2(new_n572), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n703), .A2(G29gat), .A3(new_n461), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n704), .B(KEYINPUT45), .Z(new_n705));
  OAI21_X1  g504(.A(KEYINPUT44), .B1(new_n514), .B2(new_n572), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n431), .A2(new_n512), .A3(new_n442), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n693), .A2(new_n696), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n461), .A2(new_n509), .A3(new_n436), .A4(new_n464), .ZN(new_n709));
  OAI22_X1  g508(.A1(new_n707), .A2(new_n509), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n357), .A2(new_n358), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n362), .A2(KEYINPUT38), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n712), .A3(new_n351), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n696), .B1(new_n713), .B2(new_n461), .ZN(new_n714));
  AOI211_X1 g513(.A(KEYINPUT89), .B(new_n454), .C1(new_n464), .C2(new_n436), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n458), .B1(new_n442), .B2(new_n455), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n465), .A2(new_n275), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n691), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n710), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n721), .A3(new_n571), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n701), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n726), .A2(KEYINPUT105), .A3(new_n431), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G29gat), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT105), .B1(new_n726), .B2(new_n431), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n705), .B1(new_n728), .B2(new_n729), .ZN(G1328gat));
  AND2_X1   g529(.A1(new_n549), .A2(new_n551), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n703), .A2(new_n731), .A3(new_n510), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT46), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(new_n725), .B2(new_n510), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(G1329gat));
  NAND2_X1  g534(.A1(new_n535), .A2(new_n536), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n702), .A2(new_n736), .A3(new_n693), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n725), .A2(new_n691), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n738), .B2(new_n736), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(KEYINPUT47), .Z(G1330gat));
  NOR3_X1   g539(.A1(new_n514), .A2(KEYINPUT44), .A3(new_n572), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n721), .B1(new_n720), .B2(new_n571), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n275), .B(new_n724), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G50gat), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n696), .A2(G50gat), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n702), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n744), .A2(KEYINPUT48), .A3(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n748));
  INV_X1    g547(.A(new_n746), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n744), .B2(KEYINPUT106), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n743), .A2(new_n751), .A3(G50gat), .ZN(new_n752));
  AOI211_X1 g551(.A(new_n748), .B(KEYINPUT48), .C1(new_n750), .C2(new_n752), .ZN(new_n753));
  AOI211_X1 g552(.A(new_n696), .B(new_n701), .C1(new_n706), .C2(new_n722), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT106), .B1(new_n754), .B2(new_n540), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n755), .A2(new_n752), .A3(new_n746), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT48), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT107), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n747), .B1(new_n753), .B2(new_n758), .ZN(G1331gat));
  NAND2_X1  g558(.A1(new_n642), .A2(new_n644), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n645), .A2(new_n646), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n677), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n612), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n431), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G57gat), .ZN(G1332gat));
  INV_X1    g566(.A(KEYINPUT49), .ZN(new_n768));
  INV_X1    g567(.A(G64gat), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n765), .B(new_n442), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT108), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n769), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n771), .B(new_n772), .ZN(G1333gat));
  INV_X1    g572(.A(G71gat), .ZN(new_n774));
  INV_X1    g573(.A(new_n691), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n774), .B1(new_n765), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n612), .A2(new_n693), .A3(new_n764), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT109), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n776), .B1(new_n778), .B2(new_n774), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n275), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g581(.A1(new_n762), .A2(new_n610), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n723), .A2(new_n677), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(G85gat), .B1(new_n784), .B2(new_n461), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n514), .A2(new_n572), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n786), .A2(KEYINPUT51), .A3(new_n783), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT51), .B1(new_n786), .B2(new_n783), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n431), .A2(new_n417), .A3(new_n677), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n785), .B1(new_n789), .B2(new_n790), .ZN(G1336gat));
  INV_X1    g590(.A(new_n784), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n517), .B1(new_n792), .B2(new_n442), .ZN(new_n793));
  INV_X1    g592(.A(new_n789), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n442), .A2(new_n517), .A3(new_n677), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT110), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT111), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n793), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n799), .B1(new_n789), .B2(new_n796), .ZN(new_n800));
  OAI22_X1  g599(.A1(new_n798), .A2(new_n799), .B1(new_n793), .B2(new_n800), .ZN(G1337gat));
  OAI21_X1  g600(.A(G99gat), .B1(new_n784), .B2(new_n691), .ZN(new_n802));
  OR3_X1    g601(.A1(new_n497), .A2(G99gat), .A3(new_n763), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n789), .B2(new_n803), .ZN(G1338gat));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805));
  OAI21_X1  g604(.A(G106gat), .B1(new_n784), .B2(new_n696), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n805), .B1(new_n806), .B2(KEYINPUT112), .ZN(new_n807));
  OR3_X1    g606(.A1(new_n696), .A2(G106gat), .A3(new_n763), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n806), .B1(new_n789), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n807), .B(new_n809), .ZN(G1339gat));
  AOI21_X1  g609(.A(new_n620), .B1(new_n616), .B2(new_n619), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n616), .A2(new_n629), .A3(new_n631), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(KEYINPUT113), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n630), .B2(new_n632), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n638), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n760), .A2(new_n677), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n660), .A2(new_n650), .A3(new_n662), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n821), .A2(new_n663), .A3(new_n822), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n665), .A2(new_n666), .A3(KEYINPUT10), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n649), .B1(new_n824), .B2(new_n661), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n673), .B1(new_n825), .B2(KEYINPUT54), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n820), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n674), .B1(new_n663), .B2(new_n822), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(KEYINPUT54), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n828), .B(KEYINPUT55), .C1(new_n829), .C2(new_n821), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n825), .B(new_n674), .C1(new_n649), .C2(new_n667), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n827), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n572), .B(new_n819), .C1(new_n832), .C2(new_n647), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n760), .A2(new_n818), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n571), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n700), .A3(new_n835), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n572), .A2(new_n763), .A3(new_n647), .A4(new_n610), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n836), .A2(new_n837), .A3(KEYINPUT114), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT114), .B1(new_n836), .B2(new_n837), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n838), .A2(new_n839), .A3(new_n708), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n442), .A2(new_n461), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G113gat), .B1(new_n842), .B2(new_n647), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n838), .A2(new_n839), .A3(new_n512), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n841), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n762), .A2(new_n369), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT115), .ZN(G1340gat));
  OAI21_X1  g647(.A(G120gat), .B1(new_n842), .B2(new_n763), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n677), .A2(new_n367), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n849), .B1(new_n845), .B2(new_n850), .ZN(G1341gat));
  INV_X1    g650(.A(G127gat), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n842), .A2(new_n852), .A3(new_n700), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n845), .A2(new_n700), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(KEYINPUT116), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(G127gat), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(KEYINPUT116), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(G1342gat));
  NOR3_X1   g657(.A1(new_n845), .A2(G134gat), .A3(new_n572), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT56), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT117), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(KEYINPUT117), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n859), .A2(new_n860), .ZN(new_n864));
  OAI21_X1  g663(.A(G134gat), .B1(new_n842), .B2(new_n572), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n862), .A2(new_n863), .A3(new_n864), .A4(new_n865), .ZN(G1343gat));
  NOR3_X1   g665(.A1(new_n838), .A2(new_n839), .A3(new_n696), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n837), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n762), .A2(new_n827), .A3(new_n830), .A4(new_n831), .ZN(new_n871));
  AOI22_X1  g670(.A1(new_n642), .A2(new_n644), .B1(new_n816), .B2(new_n817), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n571), .B1(new_n872), .B2(new_n677), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n610), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n870), .B1(new_n874), .B2(new_n835), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT57), .B1(new_n875), .B2(new_n696), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n691), .A2(new_n841), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT118), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n869), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G141gat), .B1(new_n879), .B2(new_n647), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n867), .A2(new_n877), .ZN(new_n881));
  INV_X1    g680(.A(G141gat), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n882), .A3(new_n762), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g684(.A(G148gat), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n881), .A2(new_n886), .A3(new_n677), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n888), .B(G148gat), .C1(new_n879), .C2(new_n763), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT119), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n696), .B1(new_n836), .B2(new_n837), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(KEYINPUT57), .ZN(new_n893));
  OAI211_X1 g692(.A(KEYINPUT121), .B(new_n868), .C1(new_n875), .C2(new_n696), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n838), .A2(new_n839), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n896), .A2(new_n897), .A3(KEYINPUT57), .A4(new_n275), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n836), .A2(new_n837), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT114), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n836), .A2(new_n837), .A3(KEYINPUT114), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n901), .A2(KEYINPUT57), .A3(new_n275), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT120), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n895), .A2(new_n898), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n677), .A3(new_n878), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n888), .B1(new_n906), .B2(G148gat), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n887), .B1(new_n890), .B2(new_n907), .ZN(G1345gat));
  AOI21_X1  g707(.A(G155gat), .B1(new_n881), .B2(new_n610), .ZN(new_n909));
  INV_X1    g708(.A(new_n879), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n700), .A2(new_n231), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(G1346gat));
  AOI21_X1  g711(.A(G162gat), .B1(new_n881), .B2(new_n571), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n572), .A2(new_n232), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n910), .B2(new_n914), .ZN(G1347gat));
  NAND2_X1  g714(.A1(new_n442), .A2(new_n461), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n844), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n918), .A2(new_n309), .A3(new_n762), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n840), .A2(new_n917), .ZN(new_n920));
  OAI21_X1  g719(.A(G169gat), .B1(new_n920), .B2(new_n647), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1348gat));
  AOI21_X1  g721(.A(G176gat), .B1(new_n918), .B2(new_n677), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n920), .A2(new_n310), .A3(new_n763), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n923), .A2(new_n924), .ZN(G1349gat));
  INV_X1    g724(.A(new_n286), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n926), .B1(new_n920), .B2(new_n700), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n844), .A2(new_n610), .A3(new_n282), .A4(new_n917), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT122), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT122), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n931), .A2(new_n932), .A3(KEYINPUT60), .A4(new_n934), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n931), .A2(KEYINPUT60), .A3(new_n934), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT60), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT123), .B1(new_n930), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n935), .B1(new_n936), .B2(new_n938), .ZN(G1350gat));
  OAI21_X1  g738(.A(G190gat), .B1(new_n920), .B2(new_n572), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT61), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n918), .A2(new_n283), .A3(new_n571), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1351gat));
  NOR2_X1   g742(.A1(new_n775), .A2(new_n916), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n867), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(G197gat), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(new_n947), .A3(new_n762), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n944), .B(KEYINPUT124), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n905), .A2(new_n762), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n948), .B1(new_n950), .B2(new_n947), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT125), .ZN(G1352gat));
  NOR3_X1   g751(.A1(new_n945), .A2(G204gat), .A3(new_n763), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT62), .ZN(new_n954));
  OAI211_X1 g753(.A(new_n893), .B(new_n894), .C1(new_n903), .C2(KEYINPUT120), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n897), .B1(new_n867), .B2(KEYINPUT57), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n677), .B(new_n949), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n957), .A2(KEYINPUT126), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n905), .A2(new_n959), .A3(new_n677), .A4(new_n949), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(G204gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n954), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n954), .B(KEYINPUT127), .C1(new_n958), .C2(new_n961), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1353gat));
  NAND3_X1  g765(.A1(new_n946), .A2(new_n213), .A3(new_n610), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n905), .A2(new_n610), .A3(new_n944), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n968), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n969));
  AOI21_X1  g768(.A(KEYINPUT63), .B1(new_n968), .B2(G211gat), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(G1354gat));
  NAND3_X1  g770(.A1(new_n946), .A2(new_n214), .A3(new_n571), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n905), .A2(new_n571), .A3(new_n949), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n972), .B1(new_n973), .B2(new_n214), .ZN(G1355gat));
endmodule


