//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 0 0 0 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n191));
  OR3_X1    g005(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G146), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT73), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(G146), .B1(new_n191), .B2(new_n192), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  AOI211_X1 g011(.A(new_n194), .B(G146), .C1(new_n191), .C2(new_n192), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n200));
  INV_X1    g014(.A(G119), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(G128), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT23), .A3(G119), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n202), .B(new_n204), .C1(G119), .C2(new_n203), .ZN(new_n205));
  XNOR2_X1  g019(.A(G119), .B(G128), .ZN(new_n206));
  XOR2_X1   g020(.A(KEYINPUT24), .B(G110), .Z(new_n207));
  AOI22_X1  g021(.A1(new_n205), .A2(G110), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n199), .A2(new_n208), .ZN(new_n209));
  OAI22_X1  g023(.A1(new_n205), .A2(G110), .B1(new_n206), .B2(new_n207), .ZN(new_n210));
  AND2_X1   g024(.A1(KEYINPUT64), .A2(G146), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT64), .A2(G146), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(new_n188), .A3(new_n190), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n210), .A2(new_n193), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G953), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(G221), .A3(G234), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n217), .B(KEYINPUT74), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT22), .B(G137), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n218), .B(new_n219), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n209), .A2(new_n215), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n220), .B1(new_n209), .B2(new_n215), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G217), .ZN(new_n224));
  INV_X1    g038(.A(G902), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(G234), .B2(new_n225), .ZN(new_n226));
  NOR3_X1   g040(.A1(new_n223), .A2(G902), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n225), .B1(new_n221), .B2(new_n222), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n228), .B(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n227), .B1(new_n230), .B2(new_n226), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT26), .B(G101), .ZN(new_n233));
  NOR2_X1   g047(.A1(G237), .A2(G953), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G210), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n233), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT2), .A2(G113), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT2), .ZN(new_n241));
  INV_X1    g055(.A(G113), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n241), .A2(new_n242), .A3(KEYINPUT67), .ZN(new_n243));
  AOI21_X1  g057(.A(KEYINPUT67), .B1(new_n241), .B2(new_n242), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n240), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(G116), .B(G119), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n246), .B(new_n240), .C1(new_n243), .C2(new_n244), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  NOR3_X1   g065(.A1(new_n211), .A2(new_n212), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G146), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(G143), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n251), .A2(G146), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n258), .B1(new_n213), .B2(G143), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n255), .A2(new_n256), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT11), .ZN(new_n263));
  INV_X1    g077(.A(G134), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(G137), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT65), .ZN(new_n266));
  INV_X1    g080(.A(G137), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G134), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n269), .A3(new_n263), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G131), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n264), .A2(G137), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n273), .B1(new_n268), .B2(new_n263), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n271), .A2(new_n272), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n272), .B1(new_n271), .B2(new_n275), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n262), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NOR4_X1   g092(.A1(new_n252), .A2(KEYINPUT1), .A3(new_n203), .A4(new_n254), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT64), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n253), .ZN(new_n281));
  NAND2_X1  g095(.A1(KEYINPUT64), .A2(G146), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(G143), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n203), .B1(new_n283), .B2(KEYINPUT1), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT64), .B(G146), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n257), .B1(new_n285), .B2(new_n251), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT66), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT66), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT1), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n289), .B1(new_n213), .B2(G143), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n288), .B(new_n259), .C1(new_n290), .C2(new_n203), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n279), .B1(new_n287), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n274), .B1(new_n270), .B2(new_n266), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n272), .ZN(new_n294));
  INV_X1    g108(.A(new_n273), .ZN(new_n295));
  INV_X1    g109(.A(new_n268), .ZN(new_n296));
  OAI21_X1  g110(.A(G131), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n278), .B1(new_n292), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n250), .B1(new_n299), .B2(KEYINPUT70), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(KEYINPUT70), .B2(new_n299), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT28), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n299), .A2(new_n250), .ZN(new_n304));
  INV_X1    g118(.A(new_n250), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n278), .B(new_n305), .C1(new_n292), .C2(new_n298), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT69), .B1(new_n307), .B2(KEYINPUT28), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT69), .ZN(new_n309));
  AOI211_X1 g123(.A(new_n309), .B(new_n302), .C1(new_n304), .C2(new_n306), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n303), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT30), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n255), .A2(new_n289), .A3(G128), .ZN(new_n313));
  OAI21_X1  g127(.A(G128), .B1(new_n252), .B2(new_n289), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n288), .B1(new_n314), .B2(new_n259), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n284), .A2(new_n286), .A3(KEYINPUT66), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n298), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n312), .B1(new_n319), .B2(new_n278), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n312), .B(new_n278), .C1(new_n292), .C2(new_n298), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n250), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n238), .A3(new_n306), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT31), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n306), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n299), .A2(KEYINPUT30), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n321), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n327), .B1(new_n329), .B2(new_n250), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(KEYINPUT31), .A3(new_n238), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n239), .A2(new_n311), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(G472), .A2(G902), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(KEYINPUT71), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT32), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n311), .A2(new_n239), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n326), .A2(new_n331), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT32), .ZN(new_n339));
  INV_X1    g153(.A(new_n334), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n307), .A2(KEYINPUT28), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n238), .A2(KEYINPUT29), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n303), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT72), .ZN(new_n346));
  OR2_X1    g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n323), .A2(new_n306), .ZN(new_n348));
  AOI21_X1  g162(.A(KEYINPUT29), .B1(new_n348), .B2(new_n239), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n349), .B1(new_n311), .B2(new_n239), .ZN(new_n350));
  AOI21_X1  g164(.A(G902), .B1(new_n345), .B2(new_n346), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n347), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G472), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n232), .B1(new_n342), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(G210), .B1(G237), .B2(G902), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n189), .B(new_n313), .C1(new_n315), .C2(new_n316), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n262), .A2(new_n189), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G224), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(G953), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n359), .B(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n364));
  INV_X1    g178(.A(G104), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT3), .B1(new_n365), .B2(G107), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT3), .ZN(new_n367));
  INV_X1    g181(.A(G107), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n368), .A3(G104), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n365), .A2(G107), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n366), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n364), .B1(new_n371), .B2(G101), .ZN(new_n372));
  INV_X1    g186(.A(G101), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n366), .A2(new_n369), .A3(new_n373), .A4(new_n370), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n248), .A2(new_n249), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n364), .A3(G101), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT75), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT75), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n371), .A2(new_n378), .A3(new_n364), .A4(G101), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n201), .A2(G116), .ZN(new_n383));
  OAI21_X1  g197(.A(KEYINPUT80), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n246), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT80), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n381), .A2(new_n386), .A3(G116), .A4(new_n201), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n384), .A2(G113), .A3(new_n385), .A4(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n370), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n365), .A2(G107), .ZN(new_n390));
  OAI21_X1  g204(.A(G101), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n249), .A2(new_n374), .A3(new_n391), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n375), .A2(new_n380), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G110), .B(G122), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n393), .A2(KEYINPUT82), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(KEYINPUT82), .B1(new_n393), .B2(new_n394), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT6), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n388), .A2(new_n392), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n377), .A2(new_n379), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n372), .A2(new_n374), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n250), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n398), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT81), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT81), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n393), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n394), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n403), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n397), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n403), .A2(new_n405), .A3(KEYINPUT6), .A4(new_n406), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n363), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT82), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n411), .B1(new_n402), .B2(new_n406), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n393), .A2(KEYINPUT82), .A3(new_n394), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n362), .A2(KEYINPUT7), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n357), .A2(new_n358), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n415), .B1(new_n357), .B2(new_n358), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n394), .B(KEYINPUT8), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n391), .A2(new_n374), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n388), .B2(new_n249), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT83), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n384), .A2(G113), .A3(new_n387), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n246), .A2(KEYINPUT5), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n392), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n427), .B1(new_n422), .B2(new_n423), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n419), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n414), .A2(new_n418), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n225), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n356), .B1(new_n410), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n433), .B1(new_n412), .B2(new_n413), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n403), .A2(new_n405), .A3(new_n406), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n409), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n363), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n430), .A2(new_n225), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n439), .A3(new_n355), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n432), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G214), .B1(G237), .B2(G902), .ZN(new_n442));
  XOR2_X1   g256(.A(new_n442), .B(KEYINPUT78), .Z(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(G113), .B(G122), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(new_n365), .ZN(new_n447));
  INV_X1    g261(.A(G237), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n216), .A3(G214), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n251), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n234), .A2(G143), .A3(G214), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(KEYINPUT18), .A2(G131), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT84), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT84), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n450), .A2(new_n456), .A3(new_n451), .A4(new_n453), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n449), .A2(new_n251), .ZN(new_n459));
  AOI21_X1  g273(.A(G143), .B1(new_n234), .B2(G214), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n454), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n188), .A2(new_n190), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G146), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n214), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n458), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n452), .A2(KEYINPUT17), .A3(G131), .ZN(new_n466));
  OAI21_X1  g280(.A(G131), .B1(new_n459), .B2(new_n460), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n450), .A2(new_n272), .A3(new_n451), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n466), .B1(new_n469), .B2(KEYINPUT17), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n447), .B(new_n465), .C1(new_n199), .C2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n447), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n464), .A2(new_n461), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n473), .B1(new_n457), .B2(new_n455), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT19), .ZN(new_n475));
  AOI21_X1  g289(.A(KEYINPUT19), .B1(new_n188), .B2(new_n190), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n213), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n469), .A2(new_n193), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n472), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n471), .A2(new_n479), .A3(KEYINPUT85), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT85), .B1(new_n471), .B2(new_n479), .ZN(new_n481));
  NOR2_X1   g295(.A1(G475), .A2(G902), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT20), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT86), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n481), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n471), .A2(new_n479), .A3(KEYINPUT85), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n482), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT86), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT20), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n471), .A2(new_n479), .ZN(new_n492));
  AOI21_X1  g306(.A(KEYINPUT20), .B1(new_n483), .B2(KEYINPUT87), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n492), .B(new_n493), .C1(KEYINPUT87), .C2(new_n483), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n486), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G478), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(KEYINPUT15), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  XOR2_X1   g312(.A(KEYINPUT9), .B(G234), .Z(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(G217), .A3(new_n216), .ZN(new_n500));
  XOR2_X1   g314(.A(G116), .B(G122), .Z(new_n501));
  INV_X1    g315(.A(KEYINPUT88), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G116), .B(G122), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT88), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n368), .ZN(new_n507));
  XNOR2_X1  g321(.A(G128), .B(G143), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n264), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n251), .A2(G128), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n203), .A2(G143), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G134), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT14), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n504), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G122), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n516), .A2(G116), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n368), .B1(new_n517), .B2(KEYINPUT14), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n509), .A2(new_n513), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n510), .A2(KEYINPUT13), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(new_n264), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n508), .A2(KEYINPUT13), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT89), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n521), .A2(new_n522), .B1(new_n509), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n508), .A2(KEYINPUT89), .A3(new_n264), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n503), .A2(new_n505), .A3(G107), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n507), .A2(new_n527), .ZN(new_n528));
  AOI221_X4 g342(.A(new_n500), .B1(new_n507), .B2(new_n519), .C1(new_n526), .C2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n500), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(new_n528), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n507), .A2(new_n519), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n225), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT90), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g350(.A(KEYINPUT90), .B(new_n225), .C1(new_n529), .C2(new_n533), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n498), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n497), .B1(new_n534), .B2(new_n535), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n216), .A2(G952), .ZN(new_n540));
  NAND2_X1  g354(.A1(G234), .A2(G237), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(G902), .A3(G953), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT21), .B(G898), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n543), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR3_X1   g361(.A1(new_n538), .A2(new_n539), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n465), .B1(new_n199), .B2(new_n470), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(new_n447), .ZN(new_n550));
  OAI21_X1  g364(.A(G475), .B1(new_n550), .B2(G902), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n495), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(G221), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n553), .B1(new_n499), .B2(new_n225), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G469), .ZN(new_n556));
  XNOR2_X1  g370(.A(G110), .B(G140), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n216), .A2(G227), .ZN(new_n558));
  XOR2_X1   g372(.A(new_n557), .B(new_n558), .Z(new_n559));
  AOI21_X1  g373(.A(new_n289), .B1(G143), .B2(new_n253), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n203), .B1(new_n560), .B2(KEYINPUT76), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT1), .B1(new_n251), .B2(G146), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT76), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n254), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n561), .A2(new_n564), .B1(new_n283), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n421), .B1(new_n566), .B2(new_n279), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT10), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n380), .A2(new_n262), .A3(new_n400), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n421), .A2(KEYINPUT10), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n292), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n276), .A2(new_n277), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n559), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n575), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n571), .B2(new_n573), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT12), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n561), .A2(new_n564), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n283), .A2(new_n565), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n420), .B1(new_n583), .B2(new_n313), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n584), .B1(new_n292), .B2(new_n420), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n580), .B1(new_n585), .B2(new_n575), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n567), .B1(new_n317), .B2(new_n421), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(KEYINPUT12), .A3(new_n577), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n586), .A2(new_n588), .B1(new_n574), .B2(new_n575), .ZN(new_n589));
  INV_X1    g403(.A(new_n559), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n579), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n556), .B1(new_n591), .B2(new_n225), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n586), .A2(new_n588), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n317), .A2(KEYINPUT10), .A3(new_n421), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n594), .A2(new_n575), .A3(new_n569), .A4(new_n570), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n578), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n593), .A2(new_n576), .B1(new_n596), .B2(new_n559), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT77), .B(G469), .Z(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n597), .A2(G902), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n555), .B1(new_n592), .B2(new_n600), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n445), .A2(new_n552), .A3(new_n601), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n354), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(new_n373), .ZN(G3));
  INV_X1    g418(.A(KEYINPUT92), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n432), .A2(new_n605), .A3(new_n440), .ZN(new_n606));
  OAI211_X1 g420(.A(KEYINPUT92), .B(new_n356), .C1(new_n410), .C2(new_n431), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n534), .A2(G478), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n496), .A2(new_n225), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OR3_X1    g425(.A1(new_n529), .A2(new_n533), .A3(KEYINPUT33), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT33), .B1(new_n529), .B2(new_n533), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n613), .A3(G478), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  AOI211_X1 g429(.A(new_n547), .B(new_n615), .C1(new_n495), .C2(new_n551), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n608), .A2(KEYINPUT93), .A3(new_n444), .A4(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT93), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n606), .A2(new_n444), .A3(new_n607), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n495), .A2(new_n551), .ZN(new_n620));
  INV_X1    g434(.A(new_n547), .ZN(new_n621));
  INV_X1    g435(.A(new_n615), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n618), .B1(new_n619), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n617), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT91), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n626), .B1(new_n332), .B2(G902), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n338), .A2(KEYINPUT91), .A3(new_n225), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n628), .A3(G472), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n338), .A2(new_n340), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n231), .B(new_n555), .C1(new_n592), .C2(new_n600), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n625), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT94), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT34), .B(G104), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  NAND2_X1  g451(.A1(new_n484), .A2(new_n485), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n486), .A2(new_n638), .A3(new_n491), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n538), .A2(new_n539), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n639), .A2(new_n640), .A3(new_n551), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n621), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n619), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n633), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT35), .B(G107), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  NAND2_X1  g460(.A1(new_n230), .A2(new_n226), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n209), .A2(new_n215), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n220), .A2(KEYINPUT36), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n650), .B(new_n225), .C1(new_n224), .C2(G234), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n602), .A2(new_n630), .A3(new_n629), .A4(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  INV_X1    g469(.A(new_n652), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n656), .B1(new_n342), .B2(new_n353), .ZN(new_n657));
  INV_X1    g471(.A(new_n601), .ZN(new_n658));
  INV_X1    g472(.A(new_n619), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n542), .B(KEYINPUT95), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n661), .B1(new_n662), .B2(new_n545), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n641), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n657), .A2(new_n658), .A3(new_n659), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  XOR2_X1   g481(.A(new_n441), .B(KEYINPUT38), .Z(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n444), .B1(new_n538), .B2(new_n539), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n495), .B2(new_n551), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n663), .B(KEYINPUT39), .Z(new_n672));
  NAND2_X1  g486(.A1(new_n658), .A2(new_n672), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n669), .B(new_n671), .C1(KEYINPUT40), .C2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(KEYINPUT40), .B2(new_n673), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n330), .A2(new_n239), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n225), .B1(new_n307), .B2(new_n238), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n342), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n652), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  NAND3_X1  g497(.A1(new_n620), .A2(new_n622), .A3(new_n664), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n657), .A2(new_n658), .A3(new_n659), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  OAI21_X1  g501(.A(G469), .B1(new_n597), .B2(G902), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n595), .A2(new_n590), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n588), .B2(new_n586), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n590), .B1(new_n578), .B2(new_n595), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n225), .B(new_n598), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n688), .A2(new_n692), .A3(new_n555), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  AOI211_X1 g508(.A(new_n232), .B(new_n694), .C1(new_n342), .C2(new_n353), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n625), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT41), .B(G113), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT96), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n696), .B(new_n698), .ZN(G15));
  NAND2_X1  g513(.A1(new_n695), .A2(new_n643), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G116), .ZN(G18));
  INV_X1    g515(.A(new_n552), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n606), .A2(new_n693), .A3(new_n444), .A4(new_n607), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n703), .A2(KEYINPUT97), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(KEYINPUT97), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n702), .B(new_n657), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT98), .B(G119), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G21));
  OAI21_X1  g522(.A(G472), .B1(new_n332), .B2(G902), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n303), .A2(new_n343), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n239), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n337), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(KEYINPUT99), .A3(new_n340), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT99), .ZN(new_n714));
  AOI22_X1  g528(.A1(new_n326), .A2(new_n331), .B1(new_n710), .B2(new_n239), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n714), .B1(new_n715), .B2(new_n334), .ZN(new_n716));
  AND4_X1   g530(.A1(new_n231), .A2(new_n709), .A3(new_n713), .A4(new_n716), .ZN(new_n717));
  AND4_X1   g531(.A1(new_n621), .A2(new_n688), .A3(new_n555), .A4(new_n692), .ZN(new_n718));
  AND4_X1   g532(.A1(new_n607), .A2(new_n718), .A3(new_n606), .A4(new_n671), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  NAND4_X1  g535(.A1(new_n709), .A2(new_n716), .A3(new_n713), .A4(new_n652), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n684), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n723), .B1(new_n704), .B2(new_n705), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT100), .B(G125), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G27));
  NAND2_X1  g540(.A1(new_n342), .A2(new_n353), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n601), .A2(new_n441), .A3(new_n443), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n727), .A2(new_n231), .A3(new_n685), .A4(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT101), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(KEYINPUT42), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n731), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n354), .A2(new_n685), .A3(new_n728), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT102), .B(G131), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G33));
  NAND4_X1  g551(.A1(new_n727), .A2(new_n665), .A3(new_n231), .A4(new_n728), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G134), .ZN(G36));
  INV_X1    g553(.A(KEYINPUT45), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n556), .B1(new_n591), .B2(new_n740), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n579), .B(KEYINPUT45), .C1(new_n589), .C2(new_n590), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n741), .A2(new_n742), .B1(G469), .B2(G902), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n600), .B1(new_n743), .B2(KEYINPUT46), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n744), .A2(KEYINPUT103), .ZN(new_n745));
  OR3_X1    g559(.A1(new_n743), .A2(KEYINPUT104), .A3(KEYINPUT46), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(KEYINPUT103), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT104), .B1(new_n743), .B2(KEYINPUT46), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n745), .A2(new_n746), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n749), .A2(new_n555), .A3(new_n672), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n432), .A2(new_n444), .A3(new_n440), .ZN(new_n751));
  INV_X1    g565(.A(new_n620), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT105), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT43), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n622), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n754), .B(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n656), .B1(new_n629), .B2(new_n630), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n756), .A2(KEYINPUT44), .A3(new_n757), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n750), .A2(new_n751), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G137), .ZN(G39));
  NAND3_X1  g577(.A1(new_n685), .A2(new_n232), .A3(new_n751), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n727), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT106), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n749), .A2(KEYINPUT47), .A3(new_n555), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT47), .B1(new_n749), .B2(new_n555), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  NOR3_X1   g584(.A1(new_n232), .A2(new_n443), .A3(new_n554), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n688), .A2(new_n692), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n772), .A2(KEYINPUT49), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(KEYINPUT49), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  OR4_X1    g589(.A1(new_n679), .A2(new_n669), .A3(new_n755), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n756), .A2(new_n661), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n751), .A2(new_n693), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n680), .A2(new_n231), .A3(new_n543), .A4(new_n779), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n752), .A2(new_n615), .ZN(new_n782));
  OAI22_X1  g596(.A1(new_n780), .A2(new_n722), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n778), .A2(new_n717), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(new_n443), .A3(new_n668), .A4(new_n693), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n772), .A2(new_n555), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n767), .A2(new_n768), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n784), .A2(new_n751), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT114), .Z(new_n793));
  OAI21_X1  g607(.A(new_n789), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n789), .B(KEYINPUT51), .C1(new_n791), .C2(new_n793), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n620), .A2(new_n622), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n540), .B1(new_n781), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n778), .A2(new_n354), .A3(new_n779), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n800), .B(KEYINPUT48), .Z(new_n801));
  NOR2_X1   g615(.A1(new_n704), .A2(new_n705), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  AOI211_X1 g617(.A(new_n799), .B(new_n801), .C1(new_n803), .C2(new_n784), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n796), .A2(new_n797), .A3(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n538), .A2(new_n539), .A3(new_n663), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n639), .A2(new_n807), .A3(new_n551), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT110), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT110), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n639), .A2(new_n807), .A3(new_n810), .A4(new_n551), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n809), .A2(new_n751), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n809), .A2(KEYINPUT111), .A3(new_n751), .A4(new_n811), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n814), .A2(new_n657), .A3(new_n658), .A4(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n722), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n685), .A3(new_n728), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n816), .A2(KEYINPUT112), .A3(new_n738), .A4(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n819), .A2(new_n735), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n354), .A2(new_n602), .B1(new_n717), .B2(new_n719), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n696), .A2(new_n700), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n798), .A2(KEYINPUT107), .ZN(new_n823));
  AOI211_X1 g637(.A(new_n547), .B(new_n443), .C1(new_n432), .C2(new_n440), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT107), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n620), .A2(new_n825), .A3(new_n622), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n823), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT108), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n823), .A2(KEYINPUT108), .A3(new_n824), .A4(new_n826), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n633), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n706), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n822), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT109), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n443), .B1(new_n432), .B2(new_n440), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n752), .A2(new_n835), .A3(new_n640), .A4(new_n621), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(new_n629), .A3(new_n630), .A4(new_n632), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n834), .B1(new_n837), .B2(new_n653), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n837), .A2(new_n653), .A3(new_n834), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n842));
  INV_X1    g656(.A(new_n816), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n818), .A2(new_n738), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n820), .A2(new_n833), .A3(new_n841), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n658), .A2(new_n664), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n671), .A2(new_n606), .A3(new_n607), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n679), .A3(new_n656), .A4(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n724), .A2(new_n666), .A3(new_n686), .A4(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT52), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n806), .B1(new_n846), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT52), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n851), .B(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n837), .A2(new_n653), .A3(new_n834), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n838), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n857), .A2(new_n822), .A3(new_n832), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n819), .A2(new_n735), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n818), .A2(new_n738), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT112), .B1(new_n860), .B2(new_n816), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n855), .A2(new_n858), .A3(new_n862), .A4(KEYINPUT53), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n853), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT54), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT113), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n853), .A2(new_n866), .A3(new_n863), .ZN(new_n867));
  OAI211_X1 g681(.A(KEYINPUT113), .B(new_n806), .C1(new_n846), .C2(new_n852), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n865), .B1(new_n869), .B2(KEYINPUT54), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n805), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(G952), .A2(G953), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n776), .B1(new_n871), .B2(new_n872), .ZN(G75));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n869), .A2(G902), .ZN(new_n875));
  INV_X1    g689(.A(G210), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n436), .B(KEYINPUT115), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n363), .B(KEYINPUT55), .Z(new_n879));
  XNOR2_X1  g693(.A(new_n878), .B(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n877), .A2(new_n881), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n216), .A2(G952), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(G51));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n869), .B(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(G469), .A2(G902), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT57), .ZN(new_n889));
  OAI22_X1  g703(.A1(new_n887), .A2(new_n889), .B1(new_n691), .B2(new_n690), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n869), .A2(G902), .A3(new_n742), .A4(new_n741), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n884), .B1(new_n890), .B2(new_n891), .ZN(G54));
  NAND4_X1  g706(.A1(new_n869), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n480), .A2(new_n481), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n893), .A2(new_n895), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n896), .A2(new_n897), .A3(new_n884), .ZN(G60));
  NAND2_X1  g712(.A1(new_n612), .A2(new_n613), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n610), .B(KEYINPUT59), .Z(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n887), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n899), .B1(new_n870), .B2(new_n900), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n902), .A2(new_n884), .A3(new_n903), .ZN(G63));
  NAND2_X1  g718(.A1(G217), .A2(G902), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT117), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT60), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n869), .A2(KEYINPUT118), .A3(new_n650), .A4(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n867), .A2(new_n650), .A3(new_n868), .A4(new_n907), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT118), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n867), .A2(new_n868), .A3(new_n907), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n884), .B1(new_n912), .B2(new_n223), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n908), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT116), .ZN(new_n915));
  XNOR2_X1  g729(.A(KEYINPUT119), .B(KEYINPUT61), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n916), .B1(new_n914), .B2(new_n915), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(G66));
  NOR2_X1   g733(.A1(new_n546), .A2(new_n360), .ZN(new_n920));
  MUX2_X1   g734(.A(new_n920), .B(new_n858), .S(new_n216), .Z(new_n921));
  OAI21_X1  g735(.A(new_n878), .B1(G898), .B2(new_n216), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n921), .B(new_n922), .Z(G69));
  AOI21_X1  g737(.A(new_n216), .B1(G227), .B2(G900), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n475), .A2(new_n476), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT120), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n329), .B(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n769), .A2(new_n762), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n823), .A2(new_n826), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n752), .A2(new_n640), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n936), .A2(new_n354), .A3(new_n672), .A4(new_n728), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n724), .A2(new_n666), .A3(new_n686), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n938), .A2(KEYINPUT121), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(KEYINPUT121), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n682), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n933), .B(new_n937), .C1(KEYINPUT62), .C2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n942), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n945));
  OR3_X1    g759(.A1(new_n944), .A2(KEYINPUT122), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(KEYINPUT122), .B1(new_n944), .B2(new_n945), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n931), .B1(new_n948), .B2(G953), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n750), .A2(new_n354), .A3(new_n849), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n941), .A2(new_n735), .A3(new_n738), .A4(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n216), .B1(new_n951), .B2(new_n932), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(G900), .B2(new_n216), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n952), .B(KEYINPUT123), .C1(G900), .C2(new_n216), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n955), .A2(new_n930), .A3(new_n956), .ZN(new_n957));
  AOI211_X1 g771(.A(new_n926), .B(new_n927), .C1(new_n949), .C2(new_n957), .ZN(new_n958));
  AND4_X1   g772(.A1(new_n925), .A2(new_n949), .A3(new_n924), .A4(new_n957), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(G72));
  INV_X1    g774(.A(new_n951), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n961), .A2(new_n858), .A3(new_n933), .ZN(new_n962));
  XNOR2_X1  g776(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n963));
  NAND2_X1  g777(.A1(G472), .A2(G902), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n348), .A2(new_n238), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n884), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n948), .A2(new_n858), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n965), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n676), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n330), .A2(new_n238), .ZN(new_n974));
  INV_X1    g788(.A(new_n324), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n864), .B(new_n965), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n970), .A2(new_n973), .A3(new_n976), .ZN(G57));
endmodule


