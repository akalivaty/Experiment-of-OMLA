//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n550, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n591, new_n592, new_n595, new_n596, new_n598,
    new_n599, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168, new_n1169;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  NAND2_X1  g031(.A1(G113), .A2(G2104), .ZN(new_n457));
  INV_X1    g032(.A(G125), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n457), .B1(new_n463), .B2(KEYINPUT67), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(KEYINPUT67), .B(G125), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(G2105), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n460), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  OAI211_X1 g047(.A(G137), .B(new_n472), .C1(new_n465), .C2(new_n466), .ZN(new_n473));
  AND3_X1   g048(.A1(new_n469), .A2(new_n471), .A3(new_n473), .ZN(G160));
  NOR2_X1   g049(.A1(new_n465), .A2(new_n466), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n475), .A2(new_n472), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  OAI211_X1 g058(.A(G138), .B(new_n472), .C1(new_n465), .C2(new_n466), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n487), .A2(new_n472), .A3(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n486), .B1(new_n475), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n488), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n461), .A2(new_n462), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT68), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n485), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(G2105), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(new_n478), .B2(G126), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  XNOR2_X1  g074(.A(KEYINPUT5), .B(G543), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G651), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT69), .B(G651), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(new_n503), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT69), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT69), .A2(G651), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n507), .A2(new_n502), .A3(KEYINPUT6), .A4(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n501), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT71), .B(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n513), .B1(new_n506), .B2(new_n509), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(new_n505), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n512), .A2(new_n515), .A3(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND2_X1  g095(.A1(new_n514), .A2(G51), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n510), .A2(G89), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n525));
  AND2_X1   g100(.A1(G63), .A2(G651), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n524), .A2(new_n525), .B1(new_n500), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n521), .A2(new_n522), .A3(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  AOI22_X1  g104(.A1(new_n500), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n517), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n510), .A2(G90), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n514), .A2(G52), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT73), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n533), .A2(new_n538), .A3(new_n534), .A4(new_n535), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(G171));
  XNOR2_X1  g115(.A(KEYINPUT74), .B(G43), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n514), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n510), .A2(G81), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n500), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n517), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT75), .ZN(G188));
  NAND2_X1  g128(.A1(new_n506), .A2(new_n509), .ZN(new_n554));
  AND2_X1   g129(.A1(G53), .A2(G543), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n554), .A2(new_n558), .A3(new_n555), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n501), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n510), .A2(G91), .B1(G651), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n560), .A2(new_n564), .ZN(G299));
  AND2_X1   g140(.A1(new_n537), .A2(new_n539), .ZN(G301));
  NAND2_X1  g141(.A1(new_n514), .A2(G49), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n510), .A2(G87), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n500), .B2(G74), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(G288));
  NAND2_X1  g145(.A1(G73), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G61), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n501), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n514), .A2(G48), .B1(new_n505), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n510), .A2(G86), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(G305));
  NAND2_X1  g151(.A1(new_n514), .A2(G47), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n510), .A2(G85), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n579), .A2(new_n517), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(G290));
  NAND2_X1  g156(.A1(G79), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G66), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n501), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n514), .A2(G54), .B1(G651), .B2(new_n584), .ZN(new_n585));
  AND3_X1   g160(.A1(new_n510), .A2(KEYINPUT10), .A3(G92), .ZN(new_n586));
  AOI21_X1  g161(.A(KEYINPUT10), .B1(new_n510), .B2(G92), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  MUX2_X1   g163(.A(new_n588), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g164(.A(new_n588), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g165(.A1(G286), .A2(G868), .ZN(new_n591));
  INV_X1    g166(.A(G299), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(G868), .ZN(G297));
  OAI21_X1  g168(.A(new_n591), .B1(new_n592), .B2(G868), .ZN(G280));
  INV_X1    g169(.A(new_n588), .ZN(new_n595));
  INV_X1    g170(.A(G559), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(G860), .ZN(G148));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G868), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g175(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g176(.A1(new_n491), .A2(new_n470), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT12), .ZN(new_n603));
  XNOR2_X1  g178(.A(KEYINPUT76), .B(KEYINPUT13), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n603), .B(new_n604), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n605), .A2(G2100), .ZN(new_n606));
  AOI22_X1  g181(.A1(G123), .A2(new_n478), .B1(new_n476), .B2(G135), .ZN(new_n607));
  NOR3_X1   g182(.A1(new_n472), .A2(KEYINPUT77), .A3(G111), .ZN(new_n608));
  OAI21_X1  g183(.A(KEYINPUT77), .B1(new_n472), .B2(G111), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n609), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n607), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(G2096), .Z(new_n612));
  NAND2_X1  g187(.A1(new_n605), .A2(G2100), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n606), .A2(new_n612), .A3(new_n613), .ZN(G156));
  XNOR2_X1  g189(.A(G2427), .B(G2438), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2430), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT15), .B(G2435), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n618), .A2(KEYINPUT14), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(G1341), .B(G1348), .ZN(new_n621));
  XNOR2_X1  g196(.A(G2443), .B(G2446), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n620), .B(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(G2451), .B(G2454), .Z(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G14), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n624), .A2(new_n627), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n629), .A2(new_n630), .ZN(G401));
  XOR2_X1   g206(.A(G2072), .B(G2078), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT17), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2067), .B(G2678), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT79), .ZN(new_n637));
  XOR2_X1   g212(.A(G2084), .B(G2090), .Z(new_n638));
  AOI21_X1  g213(.A(new_n638), .B1(new_n635), .B2(new_n632), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n636), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n637), .B2(new_n639), .ZN(new_n641));
  INV_X1    g216(.A(new_n632), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n642), .A2(new_n638), .A3(new_n634), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT18), .Z(new_n644));
  NAND3_X1  g219(.A1(new_n633), .A2(new_n638), .A3(new_n635), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n641), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT80), .ZN(new_n647));
  XOR2_X1   g222(.A(G2096), .B(G2100), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(G227));
  XOR2_X1   g224(.A(G1971), .B(G1976), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT19), .ZN(new_n651));
  XOR2_X1   g226(.A(G1956), .B(G2474), .Z(new_n652));
  XOR2_X1   g227(.A(G1961), .B(G1966), .Z(new_n653));
  AND2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT20), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n652), .A2(new_n653), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n651), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n651), .B2(new_n657), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1991), .B(G1996), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1981), .B(G1986), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G229));
  AOI22_X1  g241(.A1(new_n491), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n667), .A2(new_n472), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n476), .A2(G139), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT87), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT86), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT25), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT88), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(KEYINPUT88), .B1(new_n671), .B2(new_n674), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n668), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  MUX2_X1   g254(.A(G33), .B(new_n679), .S(G29), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G2072), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(G5), .A2(G16), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT94), .Z(new_n684));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n684), .B1(G301), .B2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(G1961), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G1966), .ZN(new_n689));
  OAI21_X1  g264(.A(KEYINPUT90), .B1(G16), .B2(G21), .ZN(new_n690));
  NOR2_X1   g265(.A1(G286), .A2(new_n685), .ZN(new_n691));
  MUX2_X1   g266(.A(new_n690), .B(KEYINPUT90), .S(new_n691), .Z(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT91), .Z(new_n693));
  AOI21_X1  g268(.A(new_n688), .B1(new_n689), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(G4), .A2(G16), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n595), .B2(G16), .ZN(new_n696));
  INV_X1    g271(.A(G1348), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G35), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G162), .B2(new_n699), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT96), .ZN(new_n703));
  INV_X1    g278(.A(G2090), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n701), .B(new_n705), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n699), .A2(G32), .ZN(new_n707));
  NAND3_X1  g282(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT89), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT26), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n476), .A2(G141), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n478), .A2(G129), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n470), .A2(G105), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n707), .B1(new_n716), .B2(new_n699), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT27), .B(G1996), .Z(new_n718));
  AOI21_X1  g293(.A(new_n706), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G2078), .ZN(new_n720));
  NOR2_X1   g295(.A1(G164), .A2(new_n699), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G27), .B2(new_n699), .ZN(new_n722));
  OAI221_X1 g297(.A(new_n719), .B1(new_n720), .B2(new_n722), .C1(new_n717), .C2(new_n718), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n547), .A2(G16), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G16), .B2(G19), .ZN(new_n725));
  INV_X1    g300(.A(G1341), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT97), .B(G1956), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n685), .A2(G20), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT23), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n592), .B2(new_n685), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n727), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n725), .A2(new_n726), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n699), .A2(G26), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT28), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n476), .A2(G140), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT85), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n740));
  INV_X1    g315(.A(G116), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(G2105), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n478), .B2(G128), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n736), .B1(new_n744), .B2(G29), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G2067), .ZN(new_n746));
  AND2_X1   g321(.A1(KEYINPUT24), .A2(G34), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n699), .B1(KEYINPUT24), .B2(G34), .ZN(new_n748));
  OAI22_X1  g323(.A1(G160), .A2(new_n699), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G2084), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT93), .B(G28), .ZN(new_n751));
  AOI21_X1  g326(.A(G29), .B1(new_n751), .B2(KEYINPUT30), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(KEYINPUT30), .B2(new_n751), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT31), .B(G11), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n753), .B(new_n754), .C1(new_n611), .C2(new_n699), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n722), .B2(new_n720), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n749), .A2(G2084), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n746), .A2(new_n750), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n731), .A2(new_n728), .ZN(new_n759));
  NOR4_X1   g334(.A1(new_n723), .A2(new_n734), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  AND4_X1   g335(.A1(new_n682), .A2(new_n694), .A3(new_n698), .A4(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n693), .A2(new_n689), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT92), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n685), .A2(G22), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G166), .B2(new_n685), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(G1971), .Z(new_n767));
  MUX2_X1   g342(.A(G6), .B(G305), .S(G16), .Z(new_n768));
  XOR2_X1   g343(.A(KEYINPUT32), .B(G1981), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n685), .A2(G23), .ZN(new_n771));
  INV_X1    g346(.A(G288), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(new_n685), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT33), .B(G1976), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n767), .A2(new_n770), .A3(new_n775), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n776), .A2(KEYINPUT34), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(KEYINPUT34), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n685), .A2(G24), .ZN(new_n779));
  INV_X1    g354(.A(G290), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(new_n685), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT83), .B(G1986), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n699), .A2(G25), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n476), .A2(G131), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT81), .Z(new_n786));
  NOR2_X1   g361(.A1(G95), .A2(G2105), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT82), .ZN(new_n788));
  INV_X1    g363(.A(G107), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n460), .B1(new_n789), .B2(G2105), .ZN(new_n790));
  AOI22_X1  g365(.A1(G119), .A2(new_n478), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n786), .A2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n784), .B1(new_n793), .B2(new_n699), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT35), .B(G1991), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n777), .A2(new_n778), .A3(new_n783), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(KEYINPUT84), .A2(KEYINPUT36), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OR2_X1    g374(.A1(KEYINPUT84), .A2(KEYINPUT36), .ZN(new_n800));
  AND3_X1   g375(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n764), .A2(new_n799), .A3(new_n801), .ZN(G311));
  OR3_X1    g377(.A1(new_n764), .A2(new_n799), .A3(new_n801), .ZN(G150));
  NAND2_X1  g378(.A1(new_n595), .A2(G559), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT38), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n514), .A2(G55), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n510), .A2(G93), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n500), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n806), .B(new_n807), .C1(new_n517), .C2(new_n808), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(new_n546), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n546), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n805), .B(new_n813), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n814), .A2(KEYINPUT39), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(KEYINPUT39), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n815), .A2(new_n816), .A3(G860), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n809), .A2(G860), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT98), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT37), .Z(new_n820));
  OR2_X1    g395(.A1(new_n817), .A2(new_n820), .ZN(G145));
  XNOR2_X1  g396(.A(new_n744), .B(new_n498), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n476), .A2(G142), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n478), .A2(G130), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n472), .A2(G118), .ZN(new_n825));
  OAI21_X1  g400(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n823), .B(new_n824), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n822), .B(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n792), .B(new_n603), .Z(new_n830));
  INV_X1    g405(.A(new_n716), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n679), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n668), .B(new_n716), .C1(new_n677), .C2(new_n678), .ZN(new_n833));
  AND3_X1   g408(.A1(new_n830), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n830), .B1(new_n833), .B2(new_n832), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n829), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n832), .A2(new_n833), .ZN(new_n837));
  INV_X1    g412(.A(new_n830), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n830), .A2(new_n832), .A3(new_n833), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n839), .A2(new_n828), .A3(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(G160), .B(new_n611), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G162), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n836), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(G37), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n843), .B1(new_n836), .B2(new_n841), .ZN(new_n847));
  OAI21_X1  g422(.A(KEYINPUT99), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n836), .A2(new_n841), .ZN(new_n849));
  INV_X1    g424(.A(new_n843), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT99), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n851), .A2(new_n852), .A3(new_n845), .A4(new_n844), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n848), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g430(.A(new_n812), .B(new_n598), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n592), .A2(new_n595), .ZN(new_n857));
  NAND2_X1  g432(.A1(G299), .A2(new_n588), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT41), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n857), .A2(KEYINPUT41), .A3(new_n858), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n861), .B1(new_n856), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(G166), .B(G305), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(KEYINPUT101), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(KEYINPUT101), .ZN(new_n871));
  XNOR2_X1  g446(.A(G288), .B(KEYINPUT100), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n872), .A2(new_n780), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n780), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n870), .B(new_n871), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  OR3_X1    g450(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT42), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n866), .A2(new_n867), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n868), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n878), .A2(new_n867), .A3(new_n866), .ZN(new_n882));
  OAI21_X1  g457(.A(G868), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(G868), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n809), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(G295));
  NAND2_X1  g461(.A1(new_n883), .A2(new_n885), .ZN(G331));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n537), .A2(G286), .A3(new_n539), .ZN(new_n889));
  AOI21_X1  g464(.A(G286), .B1(new_n537), .B2(new_n539), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n812), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(G171), .A2(G168), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n537), .A2(G286), .A3(new_n539), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(new_n813), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n863), .A2(new_n864), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT103), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n891), .A2(new_n894), .A3(new_n860), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT103), .B1(new_n895), .B2(new_n896), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n899), .A2(new_n877), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n898), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n865), .B1(new_n894), .B2(new_n891), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n877), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n845), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT43), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n877), .B1(new_n899), .B2(new_n900), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n895), .A2(new_n896), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT103), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n877), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n910), .A2(new_n911), .A3(new_n898), .A4(new_n897), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n907), .A2(new_n912), .A3(new_n913), .A4(new_n845), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n888), .B1(new_n906), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n905), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n901), .A2(KEYINPUT43), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n907), .A2(new_n912), .A3(new_n845), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n916), .A2(new_n917), .B1(new_n918), .B2(KEYINPUT43), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n915), .B1(new_n919), .B2(new_n888), .ZN(G397));
  INV_X1    g495(.A(new_n457), .ZN(new_n921));
  OAI21_X1  g496(.A(G125), .B1(new_n465), .B2(new_n466), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT67), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n472), .B1(new_n924), .B2(new_n467), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n473), .A2(G40), .A3(new_n471), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT104), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n928));
  INV_X1    g503(.A(new_n926), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n469), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(G1384), .B1(new_n493), .B2(new_n497), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n931), .A2(KEYINPUT45), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(G1996), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT46), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT126), .ZN(new_n938));
  INV_X1    g513(.A(new_n933), .ZN(new_n939));
  INV_X1    g514(.A(G2067), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n744), .B(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n939), .B1(new_n941), .B2(new_n716), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n936), .B2(new_n935), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n938), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT127), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT47), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n716), .B(G1996), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n941), .A2(new_n947), .A3(new_n795), .A4(new_n793), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n739), .A2(new_n940), .A3(new_n743), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n939), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  XOR2_X1   g525(.A(new_n792), .B(new_n795), .Z(new_n951));
  NAND2_X1  g526(.A1(new_n941), .A2(new_n947), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  OR3_X1    g529(.A1(new_n939), .A2(G1986), .A3(G290), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n954), .A2(new_n933), .B1(new_n956), .B2(KEYINPUT48), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n956), .A2(KEYINPUT48), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n950), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n946), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n945), .A2(KEYINPUT47), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT63), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n927), .A2(new_n930), .A3(new_n932), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(G8), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1976), .ZN(new_n967));
  NOR2_X1   g542(.A1(G288), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT52), .B1(G288), .B2(new_n967), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n966), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT52), .B1(new_n965), .B2(new_n968), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(KEYINPUT109), .B(G1981), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n574), .A2(new_n575), .A3(new_n974), .ZN(new_n975));
  XOR2_X1   g550(.A(KEYINPUT110), .B(G86), .Z(new_n976));
  NAND2_X1  g551(.A1(new_n510), .A2(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n574), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G1981), .ZN(new_n979));
  OAI211_X1 g554(.A(KEYINPUT49), .B(new_n975), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT49), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n574), .A2(new_n575), .A3(new_n974), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n979), .B1(new_n574), .B2(new_n977), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n966), .A2(new_n980), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT111), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n980), .A2(new_n966), .A3(new_n984), .A4(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n973), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(G303), .A2(G8), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n991));
  OR3_X1    g566(.A1(new_n990), .A2(KEYINPUT107), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT107), .B1(new_n990), .B2(new_n991), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n990), .A2(new_n991), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1384), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n498), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT50), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n932), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n999), .A2(new_n927), .A3(new_n930), .A4(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(G2090), .B1(new_n1002), .B2(KEYINPUT112), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1000), .B1(new_n498), .B2(new_n997), .ZN(new_n1004));
  AOI211_X1 g579(.A(KEYINPUT50), .B(G1384), .C1(new_n493), .C2(new_n497), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n931), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n928), .B1(new_n469), .B2(new_n929), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n922), .A2(new_n923), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1010), .A2(new_n467), .A3(new_n457), .ZN(new_n1011));
  AOI211_X1 g586(.A(KEYINPUT104), .B(new_n926), .C1(new_n1011), .C2(G2105), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT105), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n998), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n997), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT105), .B1(new_n932), .B2(KEYINPUT45), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1013), .A2(new_n1016), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT106), .B(G1971), .Z(new_n1020));
  AOI22_X1  g595(.A1(new_n1003), .A2(new_n1008), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G8), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n996), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1006), .A2(new_n704), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1022), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1026), .A2(KEYINPUT108), .A3(new_n995), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT108), .B1(new_n1026), .B2(new_n995), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n989), .B(new_n1023), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G2084), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1013), .A2(new_n1030), .A3(new_n999), .A4(new_n1001), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n932), .A2(KEYINPUT45), .ZN(new_n1032));
  AOI211_X1 g607(.A(new_n1015), .B(G1384), .C1(new_n493), .C2(new_n497), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n931), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1031), .B1(new_n1034), .B2(G1966), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1035), .A2(G8), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G168), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n963), .B1(new_n1029), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT113), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n986), .A2(new_n988), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1040), .A2(new_n972), .A3(new_n971), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1026), .A2(new_n995), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1039), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1036), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1026), .A2(new_n995), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT108), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1026), .A2(KEYINPUT108), .A3(new_n995), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1044), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n989), .B(KEYINPUT113), .C1(new_n995), .C2(new_n1026), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1043), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1038), .A2(new_n1051), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1041), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1040), .A2(new_n967), .A3(new_n772), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n965), .B1(new_n1054), .B2(new_n975), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1052), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1031), .B(G168), .C1(new_n1034), .C2(G1966), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n1059));
  AND2_X1   g634(.A1(KEYINPUT122), .A2(G8), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1035), .A2(G8), .A3(G286), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1059), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT123), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT51), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT123), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(new_n1062), .A4(new_n1061), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT62), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT62), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1065), .A2(new_n1072), .A3(new_n1069), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1074), .A2(G2078), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1034), .A2(new_n1075), .B1(new_n1002), .B2(new_n687), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1074), .B1(new_n1019), .B2(G2078), .ZN(new_n1077));
  AOI21_X1  g652(.A(G301), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1071), .A2(new_n1073), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n554), .A2(new_n558), .A3(new_n555), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n558), .B1(new_n554), .B2(new_n555), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n564), .B(new_n1081), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1081), .B1(new_n560), .B2(new_n564), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI22_X1  g664(.A1(new_n1085), .A2(new_n1086), .B1(new_n1089), .B2(KEYINPUT57), .ZN(new_n1090));
  INV_X1    g665(.A(new_n564), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT116), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT57), .B1(new_n560), .B2(KEYINPUT115), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1092), .A2(new_n1093), .A3(new_n1084), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1017), .A2(new_n927), .A3(new_n930), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1096), .A2(new_n1018), .A3(new_n1016), .A4(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT114), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1006), .B2(G1956), .ZN(new_n1100));
  INV_X1    g675(.A(G1956), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1002), .A2(KEYINPUT114), .A3(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1095), .A2(new_n1098), .A3(new_n1100), .A4(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1104));
  AOI211_X1 g679(.A(new_n1099), .B(G1956), .C1(new_n1104), .C2(new_n1013), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT114), .B1(new_n1002), .B2(new_n1101), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1095), .B1(new_n1107), .B2(new_n1098), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1002), .A2(new_n697), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n927), .A2(new_n930), .A3(new_n940), .A4(new_n932), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1110), .A2(KEYINPUT117), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(KEYINPUT117), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1109), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1113), .A2(new_n595), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1080), .B(new_n1103), .C1(new_n1108), .C2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1100), .A2(new_n1098), .A3(new_n1102), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1092), .A2(new_n1093), .A3(new_n1084), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1093), .B1(new_n1092), .B2(new_n1084), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1116), .A2(new_n1119), .B1(new_n595), .B2(new_n1113), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT118), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1115), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1103), .B1(new_n1108), .B2(KEYINPUT121), .ZN(new_n1124));
  OR3_X1    g699(.A1(new_n1116), .A2(new_n1119), .A3(KEYINPUT121), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1124), .A2(KEYINPUT61), .A3(new_n1125), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n1127));
  NAND2_X1  g702(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1127), .B1(new_n1128), .B2(new_n1103), .ZN(new_n1129));
  OR2_X1    g704(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1096), .A2(new_n934), .A3(new_n1018), .A4(new_n1016), .ZN(new_n1131));
  XOR2_X1   g706(.A(KEYINPUT58), .B(G1341), .Z(new_n1132));
  NAND2_X1  g707(.A1(new_n964), .A2(new_n1132), .ZN(new_n1133));
  AOI211_X1 g708(.A(new_n546), .B(new_n1130), .C1(new_n1131), .C2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1135));
  NAND2_X1  g710(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1135), .A2(new_n547), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1134), .B1(new_n1130), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT60), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n588), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1109), .A2(new_n1111), .A3(new_n1112), .A4(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n595), .A2(KEYINPUT60), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1141), .B(new_n1143), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n1129), .A2(new_n1138), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1123), .B1(new_n1126), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1076), .A2(new_n1077), .A3(G301), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n469), .A2(new_n929), .A3(new_n1075), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1002), .A2(new_n687), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1077), .A2(new_n1150), .ZN(new_n1151));
  OAI211_X1 g726(.A(KEYINPUT54), .B(new_n1147), .C1(new_n1151), .C2(G301), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT54), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1077), .A2(G301), .A3(new_n1150), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1153), .B1(new_n1154), .B2(new_n1078), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1070), .B(new_n1152), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1079), .B1(new_n1146), .B2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1029), .B(KEYINPUT125), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1057), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  XOR2_X1   g737(.A(G290), .B(G1986), .Z(new_n1163));
  AOI21_X1  g738(.A(new_n939), .B1(new_n953), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n962), .B1(new_n1162), .B2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g740(.A(G319), .B1(new_n629), .B2(new_n630), .ZN(new_n1167));
  NOR3_X1   g741(.A1(G229), .A2(G227), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g742(.A1(new_n854), .A2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g743(.A1(new_n919), .A2(new_n1169), .ZN(G308));
  OR2_X1    g744(.A1(new_n919), .A2(new_n1169), .ZN(G225));
endmodule


