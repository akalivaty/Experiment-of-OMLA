//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  XNOR2_X1  g000(.A(KEYINPUT71), .B(G953), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XOR2_X1   g002(.A(KEYINPUT70), .B(G237), .Z(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G101), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT11), .A3(G134), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G137), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT11), .ZN(new_n200));
  OAI211_X1 g014(.A(KEYINPUT65), .B(new_n200), .C1(new_n197), .C2(G137), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n195), .A2(G134), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT65), .B1(new_n203), .B2(new_n200), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n199), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G131), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n199), .B(new_n207), .C1(new_n202), .C2(new_n204), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(KEYINPUT66), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n205), .A2(new_n210), .A3(G131), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT64), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(new_n217), .B2(KEYINPUT64), .ZN(new_n221));
  OAI22_X1  g035(.A1(new_n219), .A2(new_n221), .B1(new_n220), .B2(new_n216), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n209), .A2(new_n211), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT67), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n214), .A2(KEYINPUT1), .A3(G146), .ZN(new_n226));
  XNOR2_X1  g040(.A(G143), .B(G146), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n226), .B1(new_n227), .B2(G128), .ZN(new_n228));
  INV_X1    g042(.A(G128), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT69), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n227), .A2(new_n233), .A3(new_n230), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n228), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n203), .A2(new_n198), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G131), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n208), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n235), .B1(KEYINPUT68), .B2(new_n238), .ZN(new_n239));
  OR2_X1    g053(.A1(new_n238), .A2(KEYINPUT68), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n209), .A2(new_n242), .A3(new_n211), .A4(new_n223), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n225), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G119), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G116), .ZN(new_n246));
  INV_X1    g060(.A(G116), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G119), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT2), .B(G113), .ZN(new_n250));
  OR2_X1    g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n250), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n244), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n253), .ZN(new_n255));
  OR2_X1    g069(.A1(new_n235), .A2(new_n238), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n224), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT28), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT28), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n224), .A2(new_n259), .A3(new_n256), .A4(new_n255), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n194), .B1(new_n254), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT31), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n224), .A2(KEYINPUT30), .A3(new_n256), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n253), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT30), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(new_n244), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n194), .A2(new_n257), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n263), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n268), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n224), .A2(KEYINPUT67), .B1(new_n239), .B2(new_n240), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT30), .B1(new_n271), .B2(new_n243), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n270), .B(KEYINPUT31), .C1(new_n272), .C2(new_n265), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n262), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(G472), .A2(G902), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT32), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n254), .A2(new_n261), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n194), .B1(new_n279), .B2(KEYINPUT29), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n224), .A2(new_n256), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n253), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n261), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n280), .B1(KEYINPUT29), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n244), .A2(new_n266), .ZN(new_n286));
  INV_X1    g100(.A(new_n265), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n194), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n257), .A3(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n285), .B1(new_n290), .B2(KEYINPUT29), .ZN(new_n291));
  OAI21_X1  g105(.A(G472), .B1(new_n284), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n278), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n262), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT31), .B1(new_n288), .B2(new_n270), .ZN(new_n295));
  AOI211_X1 g109(.A(new_n263), .B(new_n268), .C1(new_n286), .C2(new_n287), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(new_n275), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT73), .B1(new_n274), .B2(new_n276), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT74), .B(KEYINPUT32), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n299), .A2(new_n300), .A3(KEYINPUT75), .A4(new_n301), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n293), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT22), .B(G137), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(KEYINPUT79), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n308), .B(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(G125), .B(G140), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT16), .ZN(new_n312));
  INV_X1    g126(.A(G125), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n313), .A2(G140), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n312), .B(G146), .C1(KEYINPUT16), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n311), .A2(new_n212), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n229), .A2(KEYINPUT23), .A3(G119), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(KEYINPUT76), .ZN(new_n318));
  INV_X1    g132(.A(G110), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n320));
  AOI22_X1  g134(.A1(KEYINPUT77), .A2(new_n320), .B1(new_n229), .B2(G119), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(KEYINPUT77), .B2(new_n320), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n245), .A2(G128), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n318), .A2(new_n319), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n229), .A2(G119), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n323), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT24), .B(G110), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n324), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n325), .B1(new_n324), .B2(new_n329), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n315), .B(new_n316), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n327), .A2(new_n328), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n318), .A2(new_n322), .A3(new_n323), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n334), .B1(new_n335), .B2(G110), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n312), .B1(KEYINPUT16), .B2(new_n314), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n212), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n315), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n310), .B1(new_n333), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n315), .A2(new_n316), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n324), .A2(new_n329), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT78), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n342), .B1(new_n344), .B2(new_n330), .ZN(new_n345));
  INV_X1    g159(.A(new_n340), .ZN(new_n346));
  INV_X1    g160(.A(new_n310), .ZN(new_n347));
  NOR3_X1   g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n285), .B1(new_n341), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n333), .A2(new_n340), .A3(new_n310), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n347), .B1(new_n345), .B2(new_n346), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(KEYINPUT25), .A3(new_n285), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G217), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(G234), .B2(new_n285), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(G902), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n354), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n306), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(KEYINPUT9), .B(G234), .ZN(new_n364));
  OAI21_X1  g178(.A(G221), .B1(new_n364), .B2(G902), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n209), .A2(new_n211), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT83), .ZN(new_n368));
  INV_X1    g182(.A(G107), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G104), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT82), .ZN(new_n371));
  INV_X1    g185(.A(G104), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G107), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT82), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(new_n369), .A3(G104), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G101), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT3), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT80), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n378), .A2(KEYINPUT80), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n379), .B1(new_n380), .B2(new_n370), .ZN(new_n381));
  INV_X1    g195(.A(G101), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT80), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(KEYINPUT3), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n372), .A2(G107), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n381), .A2(new_n382), .A3(new_n373), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n377), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n235), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n368), .B1(new_n389), .B2(KEYINPUT10), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT10), .ZN(new_n391));
  OAI211_X1 g205(.A(KEYINPUT83), .B(new_n391), .C1(new_n235), .C2(new_n388), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n388), .A2(KEYINPUT84), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT84), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n377), .A2(new_n387), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n235), .A2(new_n391), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n390), .A2(new_n392), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n383), .A2(KEYINPUT3), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n384), .B1(new_n385), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n373), .B1(new_n379), .B2(new_n370), .ZN(new_n401));
  OAI21_X1  g215(.A(G101), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(KEYINPUT4), .A3(new_n387), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT81), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n402), .A2(new_n387), .A3(KEYINPUT81), .A4(KEYINPUT4), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT4), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n408), .B(G101), .C1(new_n400), .C2(new_n401), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n407), .A2(new_n223), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n367), .B1(new_n398), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n390), .A2(new_n392), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n396), .A2(new_n397), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n412), .A2(new_n410), .A3(new_n413), .A4(new_n367), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n188), .A2(G227), .ZN(new_n415));
  XOR2_X1   g229(.A(G110), .B(G140), .Z(new_n416));
  XNOR2_X1  g230(.A(new_n415), .B(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT86), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n411), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n414), .A2(KEYINPUT86), .A3(new_n418), .ZN(new_n422));
  INV_X1    g236(.A(new_n389), .ZN(new_n423));
  INV_X1    g237(.A(new_n235), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n423), .B1(new_n396), .B2(new_n424), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n209), .A2(KEYINPUT85), .A3(new_n211), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT12), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT12), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n425), .A2(new_n429), .A3(new_n426), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n414), .A3(new_n430), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n421), .A2(new_n422), .B1(new_n431), .B2(new_n417), .ZN(new_n432));
  OAI21_X1  g246(.A(G469), .B1(new_n432), .B2(G902), .ZN(new_n433));
  INV_X1    g247(.A(new_n414), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n417), .B1(new_n434), .B2(new_n411), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n428), .A2(new_n414), .A3(new_n430), .A4(new_n418), .ZN(new_n436));
  AOI21_X1  g250(.A(G902), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT87), .B(G469), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n366), .B1(new_n433), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n285), .B1(G234), .B2(G237), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n187), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(G898), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G952), .ZN(new_n446));
  AOI211_X1 g260(.A(G953), .B(new_n446), .C1(G234), .C2(G237), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(G214), .B1(G237), .B2(G902), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT89), .B1(new_n223), .B2(new_n313), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n235), .A2(new_n313), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT89), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n222), .A2(new_n454), .A3(G125), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n452), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G224), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT7), .B1(new_n457), .B2(G953), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n456), .B(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n246), .A2(new_n248), .A3(KEYINPUT5), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n460), .B(G113), .C1(KEYINPUT5), .C2(new_n246), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n251), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n462), .B1(new_n393), .B2(new_n395), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n463), .B1(new_n388), .B2(new_n462), .ZN(new_n464));
  XNOR2_X1  g278(.A(G110), .B(G122), .ZN(new_n465));
  XOR2_X1   g279(.A(new_n465), .B(KEYINPUT8), .Z(new_n466));
  NOR2_X1   g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n459), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n253), .A2(new_n409), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(new_n405), .B2(new_n406), .ZN(new_n470));
  INV_X1    g284(.A(new_n465), .ZN(new_n471));
  OR3_X1    g285(.A1(new_n470), .A2(new_n463), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(G902), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n471), .B1(new_n470), .B2(new_n463), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n472), .A2(new_n474), .A3(KEYINPUT6), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n457), .A2(G953), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n456), .B(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n478), .B(new_n471), .C1(new_n470), .C2(new_n463), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT88), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n479), .A2(new_n480), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n475), .B(new_n477), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n473), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(G210), .B1(G237), .B2(G902), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n473), .A2(new_n485), .A3(new_n483), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n451), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT20), .ZN(new_n490));
  NOR2_X1   g304(.A1(G475), .A2(G902), .ZN(new_n491));
  XNOR2_X1  g305(.A(G113), .B(G122), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(new_n372), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n214), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT70), .B(G237), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n187), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(G143), .A3(G214), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n495), .A2(new_n207), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n207), .B1(new_n495), .B2(new_n498), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT90), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n494), .A2(new_n214), .ZN(new_n503));
  AOI21_X1  g317(.A(G143), .B1(new_n497), .B2(G214), .ZN(new_n504));
  OAI21_X1  g318(.A(G131), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT90), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n506), .A3(new_n499), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT19), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n311), .B(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT91), .B1(new_n509), .B2(G146), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n311), .B(KEYINPUT19), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT91), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n512), .A3(new_n212), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(new_n315), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n502), .A2(new_n507), .A3(new_n515), .ZN(new_n516));
  OAI211_X1 g330(.A(KEYINPUT18), .B(G131), .C1(new_n503), .C2(new_n504), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n311), .B(new_n212), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT18), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n495), .B(new_n498), .C1(new_n519), .C2(new_n207), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n493), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n339), .B1(new_n501), .B2(KEYINPUT17), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT17), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n505), .A2(new_n524), .A3(new_n499), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n526), .A2(new_n493), .A3(new_n521), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n490), .B(new_n491), .C1(new_n522), .C2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n526), .A2(new_n493), .A3(new_n521), .ZN(new_n530));
  INV_X1    g344(.A(new_n521), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n505), .A2(new_n499), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n514), .B1(new_n532), .B2(KEYINPUT90), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n531), .B1(new_n533), .B2(new_n507), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n530), .B1(new_n534), .B2(new_n493), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n490), .B1(new_n535), .B2(new_n491), .ZN(new_n536));
  INV_X1    g350(.A(G475), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n526), .A2(new_n521), .ZN(new_n538));
  INV_X1    g352(.A(new_n493), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(G902), .B1(new_n540), .B2(new_n530), .ZN(new_n541));
  OAI22_X1  g355(.A1(new_n529), .A2(new_n536), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n364), .A2(new_n357), .A3(G953), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(G128), .B(G143), .ZN(new_n545));
  OR2_X1    g359(.A1(new_n545), .A2(G134), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(G134), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(G116), .B(G122), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT92), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n549), .A2(KEYINPUT92), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n369), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n247), .A2(KEYINPUT14), .A3(G122), .ZN(new_n554));
  INV_X1    g368(.A(new_n549), .ZN(new_n555));
  OAI211_X1 g369(.A(G107), .B(new_n554), .C1(new_n555), .C2(KEYINPUT14), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n548), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n552), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(new_n550), .A3(G107), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT13), .B1(new_n229), .B2(G143), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(new_n197), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n561), .A2(new_n545), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n545), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n553), .A2(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n544), .B1(new_n557), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n553), .A2(new_n559), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n562), .A2(new_n563), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n553), .A2(new_n556), .A3(new_n546), .A4(new_n547), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n569), .A3(new_n543), .ZN(new_n570));
  AOI21_X1  g384(.A(G902), .B1(new_n565), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(G478), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(KEYINPUT15), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  AOI211_X1 g389(.A(G902), .B(new_n573), .C1(new_n565), .C2(new_n570), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n542), .A2(new_n578), .ZN(new_n579));
  AND4_X1   g393(.A1(new_n441), .A2(new_n449), .A3(new_n489), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n363), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(G101), .ZN(G3));
  AND3_X1   g396(.A1(new_n473), .A2(new_n485), .A3(new_n483), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n485), .B1(new_n473), .B2(new_n483), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n449), .B(new_n450), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(new_n362), .ZN(new_n586));
  OAI21_X1  g400(.A(G472), .B1(new_n274), .B2(G902), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n299), .A2(new_n300), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n586), .A2(new_n589), .A3(new_n441), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n540), .A2(new_n530), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n537), .B1(new_n591), .B2(new_n285), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n522), .A2(new_n527), .ZN(new_n593));
  INV_X1    g407(.A(new_n491), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT20), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n592), .B1(new_n595), .B2(new_n528), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT93), .B1(new_n565), .B2(new_n570), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT33), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n572), .A2(G902), .ZN(new_n599));
  INV_X1    g413(.A(new_n571), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n598), .A2(new_n599), .B1(new_n572), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n590), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT34), .B(G104), .Z(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G6));
  NAND3_X1  g419(.A1(new_n590), .A2(new_n578), .A3(new_n596), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT35), .B(G107), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G9));
  NOR3_X1   g422(.A1(new_n345), .A2(new_n346), .A3(KEYINPUT94), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n310), .A2(KEYINPUT36), .ZN(new_n611));
  OAI21_X1  g425(.A(KEYINPUT94), .B1(new_n345), .B2(new_n346), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT94), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n333), .B2(new_n340), .ZN(new_n615));
  OAI22_X1  g429(.A1(new_n615), .A2(new_n609), .B1(KEYINPUT36), .B2(new_n310), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n356), .A2(new_n358), .B1(new_n360), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n589), .A2(KEYINPUT95), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT95), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n621), .B1(new_n588), .B2(new_n618), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n580), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT37), .B(G110), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G12));
  INV_X1    g439(.A(G900), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n447), .B1(new_n443), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n596), .A2(new_n578), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT96), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n631), .A3(new_n489), .ZN(new_n632));
  AOI211_X1 g446(.A(new_n366), .B(new_n618), .C1(new_n433), .C2(new_n440), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n450), .B1(new_n583), .B2(new_n584), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT96), .B1(new_n634), .B2(new_n629), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n304), .A2(new_n305), .ZN(new_n637));
  INV_X1    g451(.A(new_n293), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G128), .ZN(G30));
  XOR2_X1   g455(.A(KEYINPUT98), .B(KEYINPUT39), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n627), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n441), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT40), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT99), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT40), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n644), .B(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT99), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n487), .A2(new_n488), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n542), .A2(new_n578), .ZN(new_n654));
  NOR4_X1   g468(.A1(new_n653), .A2(new_n451), .A3(new_n619), .A4(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n288), .A2(new_n257), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n194), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n289), .A2(new_n257), .ZN(new_n658));
  AOI21_X1  g472(.A(G902), .B1(new_n658), .B2(new_n282), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  AOI22_X1  g474(.A1(new_n277), .A2(KEYINPUT32), .B1(G472), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n637), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n646), .A2(new_n650), .A3(new_n655), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G143), .ZN(G45));
  INV_X1    g478(.A(new_n601), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n542), .A2(new_n665), .A3(new_n628), .ZN(new_n666));
  OAI21_X1  g480(.A(KEYINPUT100), .B1(new_n634), .B2(new_n666), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n596), .A2(new_n601), .A3(new_n627), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT100), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n489), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n633), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n639), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  INV_X1    g487(.A(KEYINPUT101), .ZN(new_n674));
  INV_X1    g488(.A(new_n436), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n412), .A2(new_n410), .A3(new_n413), .ZN(new_n676));
  INV_X1    g490(.A(new_n367), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n418), .B1(new_n678), .B2(new_n414), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n674), .B(new_n285), .C1(new_n675), .C2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(G469), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n437), .A2(new_n674), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n365), .B(new_n440), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n602), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n683), .A2(new_n684), .A3(new_n585), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n363), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT41), .B(G113), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G15));
  INV_X1    g502(.A(new_n683), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n585), .A2(new_n577), .A3(new_n542), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n363), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  OAI21_X1  g506(.A(KEYINPUT102), .B1(new_n683), .B2(new_n634), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n285), .B1(new_n675), .B2(new_n679), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n694), .A2(new_n438), .ZN(new_n695));
  INV_X1    g509(.A(G469), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n696), .B1(new_n437), .B2(new_n674), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n694), .A2(KEYINPUT101), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n695), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT102), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n699), .A2(new_n700), .A3(new_n365), .A4(new_n489), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n693), .A2(new_n701), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n579), .A2(new_n449), .A3(new_n619), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n639), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  NOR2_X1   g519(.A1(new_n295), .A2(new_n296), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n194), .B1(new_n261), .B2(new_n282), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n275), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n587), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n362), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n634), .A2(new_n654), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n689), .A2(new_n710), .A3(new_n449), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G122), .ZN(G24));
  NAND4_X1  g527(.A1(new_n668), .A2(new_n587), .A3(new_n619), .A4(new_n708), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n693), .B2(new_n701), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT103), .B(G125), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G27));
  NAND3_X1  g531(.A1(new_n487), .A2(new_n450), .A3(new_n488), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n366), .ZN(new_n719));
  INV_X1    g533(.A(new_n362), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n421), .A2(new_n422), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n431), .A2(new_n417), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OR3_X1    g537(.A1(new_n696), .A2(KEYINPUT104), .A3(G902), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(KEYINPUT104), .B2(new_n433), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n719), .B(new_n720), .C1(new_n726), .C2(new_n695), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n306), .A2(new_n727), .A3(new_n666), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n638), .B1(KEYINPUT32), .B2(new_n277), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(KEYINPUT42), .A3(new_n668), .ZN(new_n730));
  OAI22_X1  g544(.A1(new_n728), .A2(KEYINPUT42), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G131), .ZN(G33));
  NOR3_X1   g546(.A1(new_n306), .A2(new_n727), .A3(new_n629), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n197), .ZN(G36));
  AND2_X1   g548(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n735));
  NOR2_X1   g549(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n736));
  OAI22_X1  g550(.A1(new_n542), .A2(new_n601), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n596), .A2(new_n665), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n737), .B1(new_n738), .B2(new_n736), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n588), .A3(new_n619), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n583), .A2(new_n584), .A3(new_n451), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n742), .A2(KEYINPUT106), .A3(new_n743), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(G469), .A2(G902), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n432), .A2(KEYINPUT45), .ZN(new_n750));
  OAI21_X1  g564(.A(G469), .B1(new_n432), .B2(KEYINPUT45), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT46), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n695), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n754), .B1(new_n753), .B2(new_n752), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n755), .A2(new_n365), .A3(new_n643), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n740), .A2(new_n741), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n748), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G137), .ZN(G39));
  NAND2_X1  g574(.A1(new_n755), .A2(new_n365), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(KEYINPUT47), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NOR4_X1   g577(.A1(new_n639), .A2(new_n720), .A3(new_n666), .A4(new_n718), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G140), .ZN(G42));
  NAND2_X1  g580(.A1(new_n729), .A2(new_n720), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n719), .A2(new_n447), .A3(new_n699), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n739), .A3(new_n769), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(KEYINPUT48), .Z(new_n771));
  AND3_X1   g585(.A1(new_n710), .A2(new_n739), .A3(new_n447), .ZN(new_n772));
  AOI211_X1 g586(.A(new_n446), .B(G953), .C1(new_n772), .C2(new_n702), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n769), .A2(new_n720), .ZN(new_n774));
  INV_X1    g588(.A(new_n662), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n775), .A3(new_n602), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(KEYINPUT114), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n771), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(KEYINPUT114), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n772), .A2(new_n451), .A3(new_n653), .A4(new_n689), .ZN(new_n781));
  XOR2_X1   g595(.A(new_n781), .B(KEYINPUT50), .Z(new_n782));
  NAND4_X1  g596(.A1(new_n774), .A2(new_n775), .A3(new_n596), .A4(new_n601), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n709), .A2(new_n618), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n769), .A2(new_n784), .A3(new_n739), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n782), .A2(KEYINPUT51), .A3(new_n783), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n772), .A2(new_n743), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n699), .A2(new_n366), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n787), .B1(new_n762), .B2(new_n788), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n779), .B(new_n780), .C1(new_n786), .C2(new_n789), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n762), .A2(KEYINPUT113), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n762), .A2(KEYINPUT113), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n792), .A3(new_n788), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n743), .A3(new_n772), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n794), .A2(new_n783), .A3(new_n785), .A4(new_n782), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n790), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n639), .B(new_n720), .C1(new_n685), .C2(new_n580), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n691), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n600), .A2(new_n573), .ZN(new_n800));
  INV_X1    g614(.A(new_n576), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(new_n801), .A3(KEYINPUT108), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT108), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(new_n575), .B2(new_n576), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n596), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n684), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n586), .A2(new_n807), .A3(new_n589), .A4(new_n441), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n712), .A2(new_n808), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n704), .A2(new_n809), .A3(new_n623), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT109), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n802), .A2(new_n628), .A3(new_n804), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n811), .B1(new_n542), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n805), .A2(new_n627), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n596), .A3(KEYINPUT109), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n743), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT110), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n743), .A2(new_n813), .A3(new_n815), .A4(KEYINPUT110), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n633), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n719), .B1(new_n726), .B2(new_n695), .ZN(new_n821));
  OAI22_X1  g635(.A1(new_n820), .A2(new_n306), .B1(new_n821), .B2(new_n714), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n733), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n799), .A2(new_n810), .A3(new_n823), .A4(new_n731), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT52), .ZN(new_n825));
  INV_X1    g639(.A(new_n654), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n627), .A2(new_n366), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n826), .A2(new_n489), .A3(new_n618), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n433), .A2(KEYINPUT104), .ZN(new_n829));
  INV_X1    g643(.A(new_n725), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n695), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n662), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n714), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n702), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n640), .A2(new_n672), .A3(new_n833), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT111), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n824), .B1(new_n825), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n836), .A2(KEYINPUT111), .A3(KEYINPUT52), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT53), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n823), .A2(new_n731), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n623), .A2(new_n712), .A3(new_n808), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n691), .A3(new_n704), .A4(new_n798), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n836), .A2(new_n825), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n715), .B1(new_n639), .B2(new_n636), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(KEYINPUT52), .A3(new_n672), .A4(new_n833), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT54), .B1(new_n840), .B2(new_n851), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n845), .A2(new_n847), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n850), .B1(new_n853), .B2(new_n824), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n837), .A2(new_n825), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n844), .A2(KEYINPUT53), .A3(new_n839), .A4(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(KEYINPUT112), .B(new_n850), .C1(new_n853), .C2(new_n824), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n856), .A2(new_n857), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n797), .A2(new_n852), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n862), .B1(G952), .B2(G953), .ZN(new_n863));
  INV_X1    g677(.A(new_n699), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n864), .A2(KEYINPUT49), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT107), .ZN(new_n866));
  NOR4_X1   g680(.A1(new_n738), .A2(new_n362), .A3(new_n366), .A4(new_n451), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n653), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n868), .B1(KEYINPUT49), .B2(new_n864), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n775), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n863), .A2(new_n870), .ZN(G75));
  NOR2_X1   g685(.A1(new_n188), .A2(G952), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT115), .Z(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT56), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n856), .A2(new_n859), .A3(new_n860), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(G902), .ZN(new_n877));
  INV_X1    g691(.A(G210), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n475), .B1(new_n481), .B2(new_n482), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(new_n477), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT55), .Z(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n879), .A2(new_n883), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n874), .B1(new_n884), .B2(new_n885), .ZN(G51));
  NOR2_X1   g700(.A1(new_n750), .A2(new_n751), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n876), .A2(G902), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n435), .A2(new_n436), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n860), .A2(new_n859), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT112), .B1(new_n849), .B2(new_n850), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT54), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n861), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n749), .B(KEYINPUT57), .Z(new_n896));
  AOI21_X1  g710(.A(new_n891), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT116), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n889), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n896), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n894), .B2(new_n861), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT116), .B1(new_n901), .B2(new_n891), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n872), .B1(new_n899), .B2(new_n902), .ZN(G54));
  NAND2_X1  g717(.A1(KEYINPUT58), .A2(G475), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n593), .B1(new_n877), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n905), .B1(G952), .B2(new_n188), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n877), .A2(new_n593), .A3(new_n904), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(G60));
  NAND2_X1  g722(.A1(G478), .A2(G902), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT59), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n895), .A2(new_n598), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n852), .A2(new_n861), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n598), .B1(new_n912), .B2(new_n910), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n911), .A2(new_n913), .A3(new_n874), .ZN(G63));
  NAND2_X1  g728(.A1(G217), .A2(G902), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT60), .Z(new_n916));
  NAND3_X1  g730(.A1(new_n876), .A2(new_n617), .A3(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT117), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT61), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n354), .B1(new_n876), .B2(new_n916), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n917), .A2(new_n873), .ZN(new_n921));
  OR3_X1    g735(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(G66));
  NAND2_X1  g738(.A1(new_n843), .A2(new_n188), .ZN(new_n925));
  OAI21_X1  g739(.A(G953), .B1(new_n444), .B2(new_n457), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT118), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n880), .B1(G898), .B2(new_n188), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(G69));
  AND2_X1   g744(.A1(new_n846), .A2(new_n672), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n663), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n932), .A2(KEYINPUT62), .ZN(new_n933));
  AOI22_X1  g747(.A1(new_n763), .A2(new_n764), .B1(new_n748), .B2(new_n758), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(KEYINPUT62), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n718), .B1(new_n807), .B2(KEYINPUT119), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(KEYINPUT119), .B2(new_n807), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n937), .A2(new_n644), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n363), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n933), .A2(new_n934), .A3(new_n935), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n188), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n286), .A2(new_n264), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(new_n511), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT120), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n941), .A2(KEYINPUT120), .A3(new_n943), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n945), .A2(KEYINPUT121), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n943), .B1(G900), .B2(new_n187), .ZN(new_n948));
  INV_X1    g762(.A(new_n733), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n756), .A2(new_n711), .A3(new_n768), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n931), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n934), .A2(new_n731), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n948), .B1(new_n952), .B2(new_n187), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n945), .A2(new_n946), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n947), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n946), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n957), .A2(new_n944), .ZN(new_n958));
  INV_X1    g772(.A(new_n955), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n958), .B(new_n953), .C1(KEYINPUT121), .C2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n956), .A2(new_n960), .ZN(G72));
  NAND2_X1  g775(.A1(G472), .A2(G902), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT123), .ZN(new_n963));
  XOR2_X1   g777(.A(KEYINPUT122), .B(KEYINPUT63), .Z(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT124), .Z(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(new_n940), .B2(new_n843), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n967), .A2(new_n194), .A3(new_n656), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n966), .B1(new_n952), .B2(new_n843), .ZN(new_n969));
  INV_X1    g783(.A(new_n290), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n872), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n973));
  INV_X1    g787(.A(new_n656), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n973), .B1(new_n974), .B2(new_n194), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n267), .B2(new_n268), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n974), .A2(new_n973), .A3(new_n194), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n965), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT126), .Z(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(new_n840), .B2(new_n851), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n981), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n972), .B1(new_n982), .B2(new_n983), .ZN(G57));
endmodule


