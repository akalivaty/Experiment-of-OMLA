//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n557,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1139, new_n1140, new_n1141, new_n1143;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(G173));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n456), .A2(G2106), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n458), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(KEYINPUT67), .A3(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G113), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(new_n466), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n473), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n479));
  OR2_X1    g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  INV_X1    g057(.A(G2105), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n470), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n470), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(new_n483), .B2(G112), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n485), .B(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND3_X1  g066(.A1(new_n467), .A2(new_n469), .A3(G126), .ZN(new_n492));
  NAND2_X1  g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n483), .A2(G102), .A3(G2104), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n467), .A2(new_n469), .A3(G138), .A4(new_n483), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n473), .A2(KEYINPUT4), .A3(G138), .A4(new_n483), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n495), .A2(new_n496), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  XOR2_X1   g078(.A(KEYINPUT68), .B(KEYINPUT6), .Z(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT69), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n504), .A2(new_n509), .A3(G651), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n506), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n503), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT5), .B(G543), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT70), .B(G88), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(G62), .A2(G651), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n515), .A2(new_n521), .ZN(G166));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n511), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n506), .A2(KEYINPUT71), .A3(new_n508), .A4(new_n510), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n524), .A2(G51), .A3(G543), .A4(new_n525), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n506), .A2(G89), .A3(new_n508), .A4(new_n510), .ZN(new_n527));
  NAND2_X1  g102(.A1(G63), .A2(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(new_n516), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n526), .A2(new_n530), .A3(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND4_X1  g109(.A1(new_n506), .A2(new_n508), .A3(new_n510), .A4(new_n516), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n517), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n536), .A2(G90), .B1(G651), .B2(new_n539), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n524), .A2(G52), .A3(G543), .A4(new_n525), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(G171));
  AND3_X1   g118(.A1(new_n524), .A2(G543), .A3(new_n525), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G43), .ZN(new_n545));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n517), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n536), .A2(G81), .B1(G651), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(KEYINPUT72), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT72), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(new_n544), .A2(G53), .ZN(new_n562));
  NAND2_X1  g137(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n562), .A2(new_n563), .B1(G91), .B2(new_n536), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n565), .A2(new_n507), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n544), .A2(KEYINPUT73), .A3(KEYINPUT9), .A4(G53), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(G299));
  XNOR2_X1  g143(.A(new_n542), .B(KEYINPUT74), .ZN(G301));
  INV_X1    g144(.A(G166), .ZN(G303));
  INV_X1    g145(.A(G87), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n535), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT75), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n544), .A2(G49), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(G48), .A2(G543), .ZN(new_n577));
  OR3_X1    g152(.A1(new_n511), .A2(KEYINPUT76), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT76), .B1(new_n511), .B2(new_n577), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n536), .A2(G86), .ZN(new_n581));
  AND2_X1   g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n583), .A2(new_n507), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(new_n544), .A2(G47), .ZN(new_n586));
  NAND2_X1  g161(.A1(G72), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G60), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n517), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n536), .A2(G85), .B1(G651), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n536), .A2(G92), .ZN(new_n593));
  XOR2_X1   g168(.A(new_n593), .B(KEYINPUT10), .Z(new_n594));
  NAND2_X1  g169(.A1(new_n544), .A2(G54), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n516), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n507), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n592), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n592), .B1(new_n599), .B2(G868), .ZN(G321));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(G299), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n602), .B2(G168), .ZN(G297));
  OAI21_X1  g179(.A(new_n603), .B1(new_n602), .B2(G168), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n599), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n486), .A2(G135), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT77), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n612), .A2(new_n613), .B1(G123), .B2(new_n484), .ZN(new_n614));
  NOR2_X1   g189(.A1(G99), .A2(G2105), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(new_n483), .B2(G111), .ZN(new_n616));
  OAI221_X1 g191(.A(new_n614), .B1(new_n613), .B2(new_n612), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT78), .Z(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2096), .Z(new_n619));
  NAND3_X1  g194(.A1(new_n483), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2100), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n619), .A2(new_n623), .ZN(G156));
  XNOR2_X1  g199(.A(G2427), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2430), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT15), .B(G2435), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(KEYINPUT14), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2443), .B(G2446), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT80), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n631), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G14), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT81), .ZN(G401));
  XNOR2_X1  g215(.A(G2072), .B(G2078), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT83), .Z(new_n642));
  XOR2_X1   g217(.A(G2067), .B(G2678), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT84), .B(KEYINPUT17), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n641), .B(new_n647), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n644), .B(new_n646), .C1(new_n643), .C2(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(new_n643), .A3(new_n645), .ZN(new_n650));
  INV_X1    g225(.A(new_n643), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n651), .A2(new_n641), .A3(new_n645), .ZN(new_n652));
  XOR2_X1   g227(.A(KEYINPUT82), .B(KEYINPUT18), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n649), .A2(new_n650), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2096), .B(G2100), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT86), .ZN(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT87), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(KEYINPUT87), .B1(new_n660), .B2(new_n661), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n666), .B(new_n667), .Z(new_n668));
  NOR3_X1   g243(.A1(new_n664), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT20), .Z(new_n670));
  NOR2_X1   g245(.A1(new_n660), .A2(new_n661), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n672), .A2(new_n662), .A3(new_n668), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n670), .B(new_n673), .C1(new_n668), .C2(new_n672), .ZN(new_n674));
  XOR2_X1   g249(.A(G1986), .B(G1996), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  INV_X1    g252(.A(G1981), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G1991), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n676), .B(new_n680), .ZN(G229));
  NAND2_X1  g256(.A1(new_n484), .A2(G128), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n486), .A2(G140), .ZN(new_n683));
  NOR2_X1   g258(.A1(G104), .A2(G2105), .ZN(new_n684));
  OAI21_X1  g259(.A(G2104), .B1(new_n483), .B2(G116), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n682), .B(new_n683), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G29), .ZN(new_n687));
  AND2_X1   g262(.A1(KEYINPUT88), .A2(G29), .ZN(new_n688));
  NOR2_X1   g263(.A1(KEYINPUT88), .A2(G29), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n691), .A2(KEYINPUT28), .A3(G26), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(KEYINPUT28), .B1(new_n691), .B2(G26), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT94), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G2067), .ZN(new_n697));
  NAND2_X1  g272(.A1(G171), .A2(G16), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G5), .B2(G16), .ZN(new_n699));
  INV_X1    g274(.A(G1961), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT97), .Z(new_n702));
  NAND2_X1  g277(.A1(G168), .A2(G16), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G16), .B2(G21), .ZN(new_n704));
  INV_X1    g279(.A(G1966), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n707), .A2(G32), .ZN(new_n708));
  AOI22_X1  g283(.A1(G129), .A2(new_n484), .B1(new_n486), .B2(G141), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n483), .A2(G105), .A3(G2104), .ZN(new_n710));
  NAND3_X1  g285(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT26), .Z(new_n712));
  NAND3_X1  g287(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n708), .B1(new_n713), .B2(G29), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT95), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT27), .B(G1996), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n707), .A2(G33), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n483), .A2(G103), .A3(G2104), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT25), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n486), .A2(G139), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n720), .B(new_n721), .C1(new_n483), .C2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n718), .B1(new_n723), .B2(G29), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(G2072), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT24), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(G34), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(G34), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n691), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n481), .B2(new_n707), .ZN(new_n731));
  INV_X1    g306(.A(G2084), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n725), .A2(G2072), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n717), .A2(new_n726), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT96), .ZN(new_n736));
  OAI22_X1  g311(.A1(new_n735), .A2(new_n736), .B1(new_n705), .B2(new_n704), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n700), .B2(new_n699), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT30), .B(G28), .Z(new_n739));
  OAI22_X1  g314(.A1(new_n618), .A2(new_n691), .B1(G29), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n731), .A2(new_n732), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n715), .B2(new_n716), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n691), .A2(G27), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G164), .B2(new_n691), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G2078), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n740), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT31), .B(G11), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n735), .A2(new_n736), .ZN(new_n748));
  AND3_X1   g323(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n702), .A2(new_n706), .A3(new_n738), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT98), .ZN(new_n751));
  NAND2_X1  g326(.A1(G299), .A2(G16), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(KEYINPUT23), .ZN(new_n753));
  INV_X1    g328(.A(G16), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G20), .ZN(new_n755));
  MUX2_X1   g330(.A(KEYINPUT23), .B(new_n753), .S(new_n755), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G1956), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(G1956), .ZN(new_n758));
  NOR2_X1   g333(.A1(G16), .A2(G19), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n555), .B2(G16), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(G1341), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n754), .A2(G4), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n599), .B2(new_n754), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n763), .A2(G1348), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(G1348), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n691), .A2(G35), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G162), .B2(new_n691), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT29), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G2090), .ZN(new_n769));
  NOR3_X1   g344(.A1(new_n764), .A2(new_n765), .A3(new_n769), .ZN(new_n770));
  AND3_X1   g345(.A1(new_n758), .A2(new_n761), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n751), .A2(new_n757), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G22), .ZN(new_n773));
  OAI21_X1  g348(.A(KEYINPUT92), .B1(new_n773), .B2(G16), .ZN(new_n774));
  OR3_X1    g349(.A1(new_n773), .A2(KEYINPUT92), .A3(G16), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n774), .B(new_n775), .C1(G166), .C2(new_n754), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1971), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n754), .A2(G23), .ZN(new_n778));
  INV_X1    g353(.A(G288), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(new_n754), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT33), .Z(new_n781));
  AOI21_X1  g356(.A(new_n777), .B1(new_n781), .B2(G1976), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n754), .A2(G6), .ZN(new_n783));
  INV_X1    g358(.A(G305), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n754), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT32), .B(G1981), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n782), .B(new_n787), .C1(G1976), .C2(new_n781), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(KEYINPUT34), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n690), .A2(G25), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n484), .A2(G119), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n486), .A2(G131), .ZN(new_n792));
  NOR2_X1   g367(.A1(G95), .A2(G2105), .ZN(new_n793));
  OAI21_X1  g368(.A(G2104), .B1(new_n483), .B2(G107), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n791), .B(new_n792), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT89), .Z(new_n796));
  AOI21_X1  g371(.A(new_n790), .B1(new_n796), .B2(new_n690), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT91), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT35), .B(G1991), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT90), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n798), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n754), .A2(G24), .ZN(new_n802));
  INV_X1    g377(.A(G290), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(new_n754), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1986), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n788), .B2(KEYINPUT34), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n789), .A2(new_n801), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n807), .A2(KEYINPUT93), .A3(KEYINPUT36), .ZN(new_n808));
  NAND2_X1  g383(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n789), .A2(new_n806), .A3(new_n809), .A4(new_n801), .ZN(new_n810));
  AOI211_X1 g385(.A(new_n697), .B(new_n772), .C1(new_n808), .C2(new_n810), .ZN(G311));
  AOI21_X1  g386(.A(new_n772), .B1(new_n808), .B2(new_n810), .ZN(new_n812));
  INV_X1    g387(.A(new_n697), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(G150));
  XOR2_X1   g389(.A(KEYINPUT100), .B(G55), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n544), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(G80), .A2(G543), .ZN(new_n817));
  INV_X1    g392(.A(G67), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n517), .B2(new_n818), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n536), .A2(G93), .B1(G651), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G860), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT101), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT37), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n599), .A2(G559), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT39), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n555), .A2(new_n821), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n551), .A2(new_n821), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n826), .B(new_n830), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n824), .B1(new_n833), .B2(G860), .ZN(G145));
  XNOR2_X1  g409(.A(new_n686), .B(new_n501), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n723), .B(new_n621), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n713), .B(new_n795), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n486), .A2(G142), .ZN(new_n840));
  OAI21_X1  g415(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT102), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n842), .ZN(new_n844));
  OAI211_X1 g419(.A(new_n843), .B(new_n844), .C1(G118), .C2(new_n483), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n484), .A2(G130), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n840), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n839), .B(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n618), .B(new_n481), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G162), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT103), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(G37), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n848), .A2(new_n850), .A3(KEYINPUT103), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n852), .B(new_n853), .C1(new_n850), .C2(new_n848), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g430(.A(KEYINPUT104), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n830), .B(new_n608), .Z(new_n857));
  OR2_X1    g432(.A1(G299), .A2(new_n598), .ZN(new_n858));
  NAND2_X1  g433(.A1(G299), .A2(new_n598), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT41), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(KEYINPUT41), .B1(new_n858), .B2(new_n859), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n861), .B1(new_n857), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n803), .A2(G303), .ZN(new_n867));
  NAND2_X1  g442(.A1(G290), .A2(G166), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(G288), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(G288), .B1(new_n867), .B2(new_n868), .ZN(new_n871));
  OAI21_X1  g446(.A(G305), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n871), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n873), .A2(new_n784), .A3(new_n869), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n875), .A2(KEYINPUT42), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(KEYINPUT42), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n866), .A2(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n857), .A2(new_n865), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n880), .A2(new_n861), .B1(new_n877), .B2(new_n876), .ZN(new_n881));
  OAI21_X1  g456(.A(G868), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n821), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n883), .A2(G868), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n856), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n866), .A2(new_n878), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n880), .A2(new_n861), .A3(new_n877), .A4(new_n876), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n602), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n889), .A2(KEYINPUT104), .A3(new_n884), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n886), .A2(new_n890), .ZN(G295));
  NAND2_X1  g466(.A1(new_n882), .A2(new_n885), .ZN(G331));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n893));
  INV_X1    g468(.A(G37), .ZN(new_n894));
  NAND2_X1  g469(.A1(G301), .A2(G168), .ZN(new_n895));
  NAND2_X1  g470(.A1(G171), .A2(G286), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n827), .A2(new_n829), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n883), .B1(new_n552), .B2(new_n554), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n895), .B(new_n896), .C1(new_n899), .C2(new_n828), .ZN(new_n900));
  AOI22_X1  g475(.A1(new_n898), .A2(new_n900), .B1(new_n859), .B2(new_n858), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n860), .B(new_n862), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n898), .A2(new_n900), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n901), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n875), .A2(KEYINPUT105), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n875), .A2(KEYINPUT105), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n898), .B(new_n900), .C1(new_n863), .C2(new_n864), .ZN(new_n910));
  INV_X1    g485(.A(new_n901), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n909), .B1(new_n912), .B2(new_n875), .ZN(new_n913));
  INV_X1    g488(.A(new_n875), .ZN(new_n914));
  AOI211_X1 g489(.A(KEYINPUT106), .B(new_n914), .C1(new_n910), .C2(new_n911), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n894), .B(new_n908), .C1(new_n913), .C2(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT106), .B1(new_n905), .B2(new_n914), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n912), .A2(new_n909), .A3(new_n875), .ZN(new_n920));
  AOI21_X1  g495(.A(G37), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n918), .B1(new_n921), .B2(new_n908), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n893), .B1(new_n917), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n918), .A3(new_n908), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n925), .A3(KEYINPUT44), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(G397));
  INV_X1    g502(.A(G1996), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n713), .B(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G2067), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n686), .B(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(G40), .B1(new_n479), .B2(G2105), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n933), .B1(new_n477), .B2(G2105), .ZN(new_n934));
  INV_X1    g509(.A(G1384), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT45), .B1(new_n501), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n932), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n799), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n795), .B(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n939), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(G290), .B(G1986), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n942), .B1(new_n943), .B2(new_n938), .ZN(new_n944));
  INV_X1    g519(.A(new_n493), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n945), .B1(new_n473), .B2(G126), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n496), .B1(new_n946), .B2(new_n483), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n499), .A2(new_n500), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n935), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n934), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G8), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G1976), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n954), .B1(G288), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT52), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT107), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(new_n959), .A3(KEYINPUT52), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT49), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n582), .A2(new_n678), .A3(new_n584), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n678), .B1(new_n582), .B2(new_n584), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n965), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n967), .A2(KEYINPUT49), .A3(new_n963), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n966), .A2(new_n968), .A3(new_n954), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n949), .A2(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(KEYINPUT45), .B(new_n935), .C1(new_n947), .C2(new_n948), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n934), .ZN(new_n974));
  INV_X1    g549(.A(G1971), .ZN(new_n975));
  INV_X1    g550(.A(G2090), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n949), .A2(KEYINPUT50), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n501), .A2(new_n978), .A3(new_n935), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n977), .A2(new_n934), .A3(new_n979), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n974), .A2(new_n975), .B1(new_n976), .B2(new_n980), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n981), .A2(new_n953), .ZN(new_n982));
  OAI21_X1  g557(.A(G8), .B1(new_n515), .B2(new_n521), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT55), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT52), .B1(G288), .B2(new_n955), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n986), .B(new_n954), .C1(new_n955), .C2(G288), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n961), .A2(new_n969), .A3(new_n985), .A4(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G2078), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n971), .A2(new_n934), .A3(new_n989), .A4(new_n972), .ZN(new_n990));
  XOR2_X1   g565(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n991));
  NAND3_X1  g566(.A1(new_n977), .A2(new_n934), .A3(new_n979), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n990), .A2(new_n991), .B1(new_n992), .B2(new_n700), .ZN(new_n993));
  INV_X1    g568(.A(new_n933), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n472), .A2(new_n474), .B1(G113), .B2(G2104), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n995), .A2(KEYINPUT119), .ZN(new_n996));
  OAI21_X1  g571(.A(G2105), .B1(new_n995), .B2(KEYINPUT119), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n994), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT120), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n989), .A2(KEYINPUT53), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n998), .A2(new_n999), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n1000), .A2(new_n973), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(G301), .A2(new_n993), .A3(new_n1003), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1004), .A2(KEYINPUT121), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT74), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n542), .B(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n936), .B1(new_n1008), .B2(new_n972), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n501), .A2(KEYINPUT109), .A3(KEYINPUT45), .A4(new_n935), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n934), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(new_n1011), .A3(new_n1001), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n993), .A2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n1004), .A2(KEYINPUT121), .B1(new_n1007), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT54), .B1(new_n1005), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n984), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n974), .A2(new_n975), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n980), .A2(KEYINPUT108), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n976), .B1(new_n980), .B2(KEYINPUT108), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1016), .B1(G8), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1007), .A2(new_n1013), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n542), .B1(new_n1003), .B2(new_n993), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  NOR4_X1   g600(.A1(new_n988), .A2(new_n1015), .A3(new_n1021), .A4(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n972), .A2(new_n1008), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1027), .A2(new_n971), .A3(new_n934), .A4(new_n1010), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n732), .A2(new_n980), .B1(new_n1028), .B2(new_n705), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT115), .B1(new_n1029), .B2(new_n953), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n1031));
  AND3_X1   g606(.A1(G286), .A2(new_n1031), .A3(G8), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1031), .B1(G286), .B2(G8), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1966), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n992), .A2(G2084), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1035), .B(G8), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1030), .A2(new_n1034), .A3(new_n1038), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1039), .A2(KEYINPUT116), .A3(KEYINPUT51), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT116), .B1(new_n1039), .B2(KEYINPUT51), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1034), .A2(new_n1029), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1034), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1029), .A2(new_n953), .ZN(new_n1046));
  NOR3_X1   g621(.A1(new_n1045), .A2(KEYINPUT51), .A3(new_n1046), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n1043), .A2(new_n1044), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1041), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1042), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1039), .A2(KEYINPUT116), .A3(KEYINPUT51), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1047), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT117), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1026), .B1(new_n1048), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT122), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT61), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n1059));
  NAND2_X1  g634(.A1(G299), .A2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n564), .A2(KEYINPUT57), .A3(new_n566), .A4(new_n567), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT56), .B(G2072), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  OAI22_X1  g638(.A1(new_n974), .A2(new_n1063), .B1(G1956), .B2(new_n980), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1060), .A2(new_n1061), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1064), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1058), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT111), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n973), .A2(new_n928), .A3(new_n934), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT110), .B(KEYINPUT58), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1071), .B(G1341), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n951), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1069), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n555), .A2(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1075), .B(KEYINPUT59), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1064), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1079), .A2(KEYINPUT61), .A3(new_n1065), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1068), .A2(new_n1076), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT112), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT113), .ZN(new_n1083));
  INV_X1    g658(.A(G1348), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n952), .A2(new_n930), .B1(new_n992), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT60), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n599), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1083), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1087), .B(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(KEYINPUT60), .B2(new_n1085), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT112), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1068), .A2(new_n1076), .A3(new_n1080), .A4(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1082), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n598), .A2(new_n1085), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1079), .B1(new_n1066), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1026), .B(KEYINPUT122), .C1(new_n1048), .C2(new_n1054), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1057), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1046), .A2(G168), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1099), .A2(KEYINPUT63), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n985), .B1(new_n1021), .B2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1101), .A2(new_n987), .A3(new_n961), .A4(new_n969), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n969), .A2(new_n955), .A3(new_n779), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n954), .B1(new_n1103), .B2(new_n964), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n982), .A2(new_n984), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n961), .A2(new_n969), .A3(new_n987), .A4(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT63), .B1(new_n1106), .B2(new_n1099), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1102), .A2(new_n1104), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1098), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1044), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1052), .A2(KEYINPUT117), .A3(new_n1053), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1007), .A2(new_n1013), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n988), .A2(new_n1114), .A3(new_n1021), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1113), .A2(KEYINPUT123), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT123), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1111), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n944), .B1(new_n1109), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n937), .A2(G1996), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT46), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1121), .B(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n931), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n938), .B1(new_n1125), .B2(new_n713), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1124), .B(new_n1126), .C1(new_n1122), .C2(KEYINPUT46), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT47), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n796), .A2(new_n940), .ZN(new_n1129));
  OAI22_X1  g704(.A1(new_n932), .A2(new_n1129), .B1(G2067), .B2(new_n686), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n938), .ZN(new_n1131));
  NOR3_X1   g706(.A1(G290), .A2(G1986), .A3(new_n937), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1132), .B(KEYINPUT125), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT48), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1128), .B(new_n1131), .C1(new_n1134), .C2(new_n942), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT126), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1120), .A2(new_n1136), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g712(.A1(G229), .A2(new_n463), .ZN(new_n1139));
  NAND2_X1  g713(.A1(new_n854), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g714(.A1(new_n639), .A2(new_n657), .ZN(new_n1141));
  AOI211_X1 g715(.A(new_n1140), .B(new_n1141), .C1(new_n924), .C2(new_n925), .ZN(G308));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n924), .B2(new_n925), .ZN(new_n1143));
  NAND3_X1  g717(.A1(new_n1143), .A2(new_n854), .A3(new_n1139), .ZN(G225));
endmodule


