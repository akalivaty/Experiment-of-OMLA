//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n868, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991, new_n992;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT66), .B(G190gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT27), .B(G183gat), .ZN(new_n204));
  AOI21_X1  g003(.A(KEYINPUT68), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(KEYINPUT28), .ZN(new_n206));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G169gat), .ZN(new_n210));
  INV_X1    g009(.A(G176gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT69), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n212), .A2(KEYINPUT26), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n212), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n205), .A2(KEYINPUT28), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G183gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n218), .B1(new_n203), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT24), .B1(new_n207), .B2(KEYINPUT65), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(KEYINPUT65), .B2(new_n207), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT23), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G169gat), .B2(G176gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n223), .A2(KEYINPUT25), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n230));
  INV_X1    g029(.A(G190gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n219), .A2(new_n231), .A3(KEYINPUT64), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT24), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n207), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(G183gat), .B2(G190gat), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n232), .A2(new_n234), .A3(new_n236), .A4(new_n217), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT25), .B1(new_n228), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  AND3_X1   g038(.A1(new_n229), .A2(new_n230), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n230), .B1(new_n229), .B2(new_n239), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n216), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G127gat), .B(G134gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT70), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n245));
  INV_X1    g044(.A(G127gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n246), .A3(G134gat), .ZN(new_n247));
  INV_X1    g046(.A(G113gat), .ZN(new_n248));
  INV_X1    g047(.A(G120gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G113gat), .A2(G120gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n244), .B(new_n247), .C1(KEYINPUT1), .C2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT71), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n250), .A2(KEYINPUT71), .A3(new_n251), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n255), .A2(new_n256), .A3(new_n243), .A4(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT72), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT72), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n253), .A2(new_n258), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n242), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n228), .A2(KEYINPUT25), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n265), .B1(new_n222), .B2(new_n220), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT67), .B1(new_n266), .B2(new_n238), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n229), .A2(new_n230), .A3(new_n239), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n260), .A2(new_n262), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n270), .A3(new_n216), .ZN(new_n271));
  NAND2_X1  g070(.A1(G227gat), .A2(G233gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n264), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT34), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT34), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n264), .A2(new_n271), .A3(new_n275), .A4(new_n272), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(G15gat), .B(G43gat), .Z(new_n278));
  XNOR2_X1  g077(.A(G71gat), .B(G99gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n272), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n242), .A2(new_n263), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n270), .B1(new_n269), .B2(new_n216), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT73), .B(KEYINPUT33), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n281), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n277), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n272), .B1(new_n264), .B2(new_n271), .ZN(new_n289));
  INV_X1    g088(.A(new_n286), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n280), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(new_n274), .A3(new_n276), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n285), .A2(KEYINPUT32), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n288), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n294), .B1(new_n288), .B2(new_n292), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n202), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n288), .A2(new_n292), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n293), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n288), .A2(new_n292), .A3(new_n294), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(KEYINPUT36), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G1gat), .B(G29gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT0), .ZN(new_n304));
  XNOR2_X1  g103(.A(G57gat), .B(G85gat), .ZN(new_n305));
  XOR2_X1   g104(.A(new_n304), .B(new_n305), .Z(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G225gat), .A2(G233gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT81), .B(G141gat), .ZN(new_n310));
  INV_X1    g109(.A(G148gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n311), .A2(G141gat), .ZN(new_n313));
  INV_X1    g112(.A(G155gat), .ZN(new_n314));
  INV_X1    g113(.A(G162gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NOR3_X1   g115(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n317));
  OAI22_X1  g116(.A1(new_n312), .A2(new_n313), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n311), .A2(G141gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT2), .ZN(new_n320));
  OAI22_X1  g119(.A1(new_n313), .A2(new_n319), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT79), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(G155gat), .B2(G162gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n314), .A2(new_n315), .A3(KEYINPUT79), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n316), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT80), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n321), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI211_X1 g126(.A(KEYINPUT80), .B(new_n316), .C1(new_n323), .C2(new_n324), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n318), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n253), .A2(new_n258), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n329), .A2(new_n259), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n309), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT5), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT4), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n330), .A2(new_n260), .A3(new_n262), .ZN(new_n338));
  AOI22_X1  g137(.A1(KEYINPUT82), .A2(new_n337), .B1(new_n338), .B2(KEYINPUT4), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n333), .A2(new_n340), .A3(new_n336), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n331), .B1(KEYINPUT3), .B2(new_n329), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n330), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n309), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n335), .B1(new_n342), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT5), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n338), .A2(new_n336), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n333), .A2(KEYINPUT4), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n346), .A2(new_n348), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n307), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n346), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n354), .B1(new_n339), .B2(new_n341), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n351), .B(new_n306), .C1(new_n355), .C2(new_n335), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT6), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n353), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  OAI211_X1 g157(.A(KEYINPUT6), .B(new_n307), .C1(new_n347), .C2(new_n352), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n267), .A2(new_n268), .B1(new_n209), .B2(new_n215), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n361), .B1(new_n362), .B2(KEYINPUT29), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n364));
  XOR2_X1   g163(.A(G211gat), .B(G218gat), .Z(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  XOR2_X1   g165(.A(KEYINPUT74), .B(G197gat), .Z(new_n367));
  INV_X1    g166(.A(G204gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT74), .B(G197gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G204gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G211gat), .A2(G218gat), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT22), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n366), .B1(new_n376), .B2(KEYINPUT75), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n369), .A2(new_n371), .B1(new_n374), .B2(new_n373), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT75), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n378), .A2(new_n379), .A3(new_n365), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n364), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n376), .A2(KEYINPUT75), .A3(new_n366), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n365), .B1(new_n378), .B2(new_n379), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(new_n383), .A3(KEYINPUT76), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n209), .A2(new_n215), .B1(new_n229), .B2(new_n239), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n386), .B1(new_n387), .B2(new_n361), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n229), .A2(new_n239), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n216), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n361), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(KEYINPUT77), .A3(new_n391), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n363), .A2(new_n385), .A3(new_n388), .A4(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n391), .A2(KEYINPUT29), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n362), .A2(new_n391), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n381), .A2(new_n384), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  XOR2_X1   g196(.A(G8gat), .B(G36gat), .Z(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(KEYINPUT78), .ZN(new_n399));
  XNOR2_X1  g198(.A(G64gat), .B(G92gat), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n399), .B(new_n400), .Z(new_n401));
  NAND3_X1  g200(.A1(new_n393), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n401), .B1(new_n393), .B2(new_n397), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n402), .B1(new_n403), .B2(KEYINPUT30), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n393), .A2(new_n397), .ZN(new_n405));
  INV_X1    g204(.A(new_n401), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n405), .A2(KEYINPUT30), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n360), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G78gat), .B(G106gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT31), .B(G50gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(new_n412), .B(KEYINPUT83), .Z(new_n413));
  INV_X1    g212(.A(G228gat), .ZN(new_n414));
  INV_X1    g213(.A(G233gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT29), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n382), .A2(new_n383), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n344), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n417), .B1(new_n420), .B2(new_n329), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n418), .B1(new_n329), .B2(KEYINPUT3), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT85), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n385), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n422), .A2(new_n423), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n421), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT84), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n381), .A2(new_n422), .A3(new_n384), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n376), .A2(new_n366), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n418), .B1(new_n378), .B2(new_n365), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n344), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n329), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n428), .B1(new_n434), .B2(new_n417), .ZN(new_n435));
  AOI211_X1 g234(.A(KEYINPUT84), .B(new_n416), .C1(new_n429), .C2(new_n433), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n427), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT86), .B(G22gat), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n427), .B(new_n438), .C1(new_n435), .C2(new_n436), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n413), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n437), .A2(G22gat), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n444), .A2(new_n441), .A3(new_n412), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n409), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n343), .A2(new_n345), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n349), .A2(new_n447), .A3(new_n350), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n309), .ZN(new_n449));
  OR2_X1    g248(.A1(new_n332), .A2(new_n333), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n449), .B(KEYINPUT39), .C1(new_n309), .C2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT39), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n448), .A2(new_n452), .A3(new_n309), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT87), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n453), .A2(new_n454), .A3(new_n306), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n454), .B1(new_n453), .B2(new_n306), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n451), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT40), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n353), .ZN(new_n460));
  OAI22_X1  g259(.A1(new_n404), .A2(new_n407), .B1(new_n457), .B2(new_n458), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n444), .A2(new_n441), .A3(new_n412), .ZN(new_n462));
  OAI22_X1  g261(.A1(new_n460), .A2(new_n461), .B1(new_n462), .B2(new_n442), .ZN(new_n463));
  INV_X1    g262(.A(new_n403), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n392), .A2(new_n388), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n385), .B1(new_n465), .B2(new_n363), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT37), .B1(new_n395), .B2(new_n396), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT88), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT38), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n391), .B1(new_n242), .B2(new_n418), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n392), .A2(new_n388), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n396), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT37), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n390), .A2(new_n394), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(new_n242), .B2(new_n361), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n473), .B1(new_n475), .B2(new_n385), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT88), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n472), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n468), .A2(new_n469), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n405), .A2(new_n473), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n401), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n464), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n406), .B1(new_n405), .B2(new_n473), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n393), .A2(KEYINPUT37), .A3(new_n397), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n469), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n482), .A2(new_n360), .A3(new_n485), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n302), .B(new_n446), .C1(new_n463), .C2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT35), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(KEYINPUT89), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n409), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(KEYINPUT89), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n443), .A2(new_n445), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n295), .A2(new_n296), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n490), .A2(new_n491), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n300), .B(new_n299), .C1(new_n462), .C2(new_n442), .ZN(new_n495));
  OAI211_X1 g294(.A(KEYINPUT89), .B(new_n488), .C1(new_n495), .C2(new_n409), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n487), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(new_n314), .ZN(new_n499));
  XNOR2_X1  g298(.A(G183gat), .B(G211gat), .ZN(new_n500));
  XOR2_X1   g299(.A(new_n499), .B(new_n500), .Z(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(G71gat), .A2(G78gat), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT100), .ZN(new_n505));
  NAND2_X1  g304(.A1(G71gat), .A2(G78gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n506), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT100), .B1(new_n508), .B2(new_n503), .ZN(new_n509));
  AND2_X1   g308(.A1(G57gat), .A2(G64gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(G57gat), .A2(G64gat), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT9), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n507), .A2(new_n509), .A3(new_n512), .A4(new_n514), .ZN(new_n515));
  OR2_X1    g314(.A1(G57gat), .A2(G64gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(G57gat), .A2(G64gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(KEYINPUT99), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT99), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n519), .B1(new_n510), .B2(new_n511), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n518), .A2(new_n520), .A3(new_n514), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT98), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n504), .A2(new_n522), .A3(new_n506), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT98), .B1(new_n508), .B2(new_n503), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n515), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n527), .A2(KEYINPUT21), .ZN(new_n528));
  NAND2_X1  g327(.A1(G231gat), .A2(G233gat), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n528), .B(new_n529), .Z(new_n530));
  OR2_X1    g329(.A1(new_n530), .A2(new_n246), .ZN(new_n531));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT16), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n532), .B1(new_n533), .B2(G1gat), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(G1gat), .B2(new_n532), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(G8gat), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n536), .B1(KEYINPUT21), .B2(new_n527), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n530), .A2(new_n246), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n531), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n538), .B1(new_n531), .B2(new_n539), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n502), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n542), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n544), .A2(new_n540), .A3(new_n501), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  AND2_X1   g345(.A1(G232gat), .A2(G233gat), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(KEYINPUT41), .ZN(new_n548));
  XNOR2_X1  g347(.A(G134gat), .B(G162gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT93), .ZN(new_n552));
  XNOR2_X1  g351(.A(KEYINPUT92), .B(G36gat), .ZN(new_n553));
  INV_X1    g352(.A(G29gat), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(G36gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT92), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT92), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(G36gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(KEYINPUT93), .A3(G29gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G43gat), .A2(G50gat), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(G43gat), .A2(G50gat), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT15), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(G43gat), .ZN(new_n567));
  INV_X1    g366(.A(G50gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT15), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n570), .A3(new_n563), .ZN(new_n571));
  NOR2_X1   g370(.A1(G29gat), .A2(G36gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT91), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT14), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(KEYINPUT91), .A2(KEYINPUT14), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n572), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n572), .A2(new_n576), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n566), .B(new_n571), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  AND2_X1   g378(.A1(KEYINPUT91), .A2(KEYINPUT14), .ZN(new_n580));
  NOR2_X1   g379(.A1(KEYINPUT91), .A2(KEYINPUT14), .ZN(new_n581));
  OAI22_X1  g380(.A1(new_n580), .A2(new_n581), .B1(G29gat), .B2(G36gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n572), .A2(new_n576), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n582), .A2(new_n583), .B1(new_n560), .B2(G29gat), .ZN(new_n584));
  OAI22_X1  g383(.A1(new_n562), .A2(new_n579), .B1(new_n584), .B2(new_n566), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT94), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT17), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n566), .A2(new_n571), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n582), .A2(new_n583), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n588), .A2(new_n589), .A3(new_n555), .A4(new_n561), .ZN(new_n590));
  INV_X1    g389(.A(new_n566), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n577), .A2(new_n578), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n553), .A2(new_n554), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT94), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n590), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n586), .A2(new_n587), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT95), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT95), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n586), .A2(new_n596), .A3(new_n599), .A4(new_n587), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT101), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(G85gat), .A3(G92gat), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT7), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  INV_X1    g405(.A(G85gat), .ZN(new_n607));
  INV_X1    g406(.A(G92gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n602), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n605), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G99gat), .B(G106gat), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n605), .A2(new_n609), .A3(new_n612), .A4(new_n610), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT96), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(new_n585), .B2(new_n587), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n590), .A2(new_n594), .A3(KEYINPUT96), .A4(KEYINPUT17), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n601), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G190gat), .B(G218gat), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n586), .A2(new_n596), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  AOI22_X1  g425(.A1(new_n626), .A2(new_n617), .B1(KEYINPUT41), .B2(new_n547), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n622), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n624), .B1(new_n622), .B2(new_n627), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n551), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n630), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n632), .A2(new_n550), .A3(new_n628), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G230gat), .A2(G233gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n526), .A2(new_n616), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT10), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n518), .A2(new_n520), .A3(new_n514), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n639), .A2(new_n524), .A3(new_n523), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n640), .A2(new_n515), .A3(new_n615), .A4(new_n614), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n637), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n527), .A2(KEYINPUT10), .A3(new_n617), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n636), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n637), .A2(new_n641), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n644), .B1(new_n645), .B2(new_n636), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G120gat), .B(G148gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(G176gat), .B(G204gat), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n648), .B(new_n649), .Z(new_n650));
  NAND3_X1  g449(.A1(new_n647), .A2(KEYINPUT102), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n650), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n652), .B1(new_n646), .B2(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n546), .A2(new_n634), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G113gat), .B(G141gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT90), .B(G197gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT11), .B(G169gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT12), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n536), .B1(new_n619), .B2(new_n620), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n601), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT97), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(KEYINPUT18), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(G229gat), .A2(G233gat), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n626), .A2(new_n536), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n666), .A2(new_n669), .A3(new_n670), .A4(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n536), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n625), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n670), .B(KEYINPUT13), .Z(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n625), .A2(new_n673), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n678), .B1(new_n601), .B2(new_n665), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n669), .B1(new_n679), .B2(new_n670), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n664), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n670), .A3(new_n671), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n668), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n683), .A2(new_n676), .A3(new_n672), .A4(new_n663), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n657), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n497), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n360), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G1gat), .ZN(G1324gat));
  INV_X1    g490(.A(new_n408), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT104), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G8gat), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT42), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT16), .B(G8gat), .ZN(new_n697));
  OR3_X1    g496(.A1(new_n693), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n694), .A2(new_n697), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n700));
  OAI211_X1 g499(.A(new_n695), .B(new_n698), .C1(new_n699), .C2(new_n700), .ZN(G1325gat));
  INV_X1    g500(.A(new_n688), .ZN(new_n702));
  OAI21_X1  g501(.A(G15gat), .B1(new_n702), .B2(new_n302), .ZN(new_n703));
  INV_X1    g502(.A(new_n493), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n704), .A2(G15gat), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n702), .B2(new_n705), .ZN(G1326gat));
  INV_X1    g505(.A(new_n492), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n688), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT105), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT43), .B(G22gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1327gat));
  INV_X1    g510(.A(new_n634), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n497), .A2(new_n712), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n546), .A2(new_n686), .A3(new_n655), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n716), .A2(new_n554), .A3(new_n689), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT45), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(KEYINPUT44), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n713), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n723));
  NAND3_X1  g522(.A1(new_n497), .A2(new_n712), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n715), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT107), .B1(new_n726), .B2(new_n360), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G29gat), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n726), .A2(KEYINPUT107), .A3(new_n360), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n718), .B1(new_n728), .B2(new_n729), .ZN(G1328gat));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n408), .A2(new_n560), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT46), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n553), .B1(new_n725), .B2(new_n692), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n731), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n733), .B(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n735), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(new_n739), .A3(KEYINPUT108), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n736), .A2(new_n740), .ZN(G1329gat));
  INV_X1    g540(.A(new_n302), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G43gat), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n713), .A2(new_n704), .A3(new_n715), .ZN(new_n744));
  OAI22_X1  g543(.A1(new_n726), .A2(new_n743), .B1(G43gat), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g545(.A(new_n568), .B1(new_n725), .B2(new_n707), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT48), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n707), .A2(new_n568), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT109), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n716), .A2(new_n750), .ZN(new_n751));
  OR3_X1    g550(.A1(new_n747), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n748), .B1(new_n747), .B2(new_n751), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(G1331gat));
  INV_X1    g553(.A(new_n546), .ZN(new_n755));
  NOR4_X1   g554(.A1(new_n755), .A2(new_n685), .A3(new_n712), .A4(new_n656), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n497), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n689), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g558(.A(new_n408), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n761), .B(new_n762), .Z(G1333gat));
  NAND2_X1  g562(.A1(new_n757), .A2(new_n742), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n704), .A2(G71gat), .ZN(new_n765));
  AOI22_X1  g564(.A1(new_n764), .A2(G71gat), .B1(new_n757), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g566(.A1(new_n757), .A2(new_n707), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G78gat), .ZN(G1335gat));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n546), .A2(new_n685), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n497), .A2(new_n712), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n497), .A2(KEYINPUT51), .A3(new_n712), .A4(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n776), .A2(new_n607), .A3(new_n689), .A4(new_n655), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n771), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(new_n656), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n722), .B2(new_n724), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n607), .B1(new_n782), .B2(new_n689), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n770), .B1(new_n778), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n783), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n785), .A2(KEYINPUT110), .A3(new_n777), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(G1336gat));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n497), .A2(new_n712), .A3(new_n723), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n720), .B1(new_n497), .B2(new_n712), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n692), .B(new_n780), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G92gat), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n408), .A2(G92gat), .A3(new_n656), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n795));
  AND4_X1   g594(.A1(new_n788), .A2(new_n792), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n791), .A2(G92gat), .B1(new_n776), .B2(new_n793), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n788), .B1(new_n797), .B2(new_n795), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n796), .B1(new_n799), .B2(new_n800), .ZN(G1337gat));
  INV_X1    g600(.A(G99gat), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n782), .A2(new_n742), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n805), .B1(new_n804), .B2(new_n803), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n776), .A2(new_n802), .A3(new_n493), .A4(new_n655), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(G1338gat));
  NOR2_X1   g607(.A1(new_n492), .A2(new_n656), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n776), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(G106gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT53), .ZN(new_n814));
  OR2_X1    g613(.A1(new_n813), .A2(KEYINPUT53), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n492), .A2(new_n811), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n780), .B(new_n816), .C1(new_n789), .C2(new_n790), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n812), .A2(new_n814), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(G106gat), .B1(new_n776), .B2(new_n809), .ZN(new_n819));
  INV_X1    g618(.A(new_n817), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n813), .B(KEYINPUT53), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n818), .A2(new_n821), .ZN(G1339gat));
  NOR2_X1   g621(.A1(new_n657), .A2(new_n685), .ZN(new_n823));
  OAI22_X1  g622(.A1(new_n679), .A2(new_n670), .B1(new_n674), .B2(new_n675), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n662), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n684), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n642), .A2(new_n643), .A3(new_n636), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n642), .A2(new_n643), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n635), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT115), .A4(new_n636), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n829), .A2(new_n831), .A3(KEYINPUT54), .A4(new_n832), .ZN(new_n833));
  XOR2_X1   g632(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n834));
  AOI21_X1  g633(.A(new_n650), .B1(new_n644), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(KEYINPUT55), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n646), .A2(new_n650), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n833), .A2(new_n835), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n837), .B1(new_n836), .B2(new_n838), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n712), .A2(new_n826), .A3(new_n845), .ZN(new_n846));
  AOI22_X1  g645(.A1(new_n655), .A2(new_n826), .B1(new_n845), .B2(new_n685), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(new_n712), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n823), .B1(new_n848), .B2(new_n755), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(new_n707), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n692), .A2(new_n360), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n493), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(G113gat), .B1(new_n852), .B2(new_n686), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n849), .A2(new_n360), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n495), .A2(new_n692), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n856), .B(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n685), .A2(new_n248), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n853), .B1(new_n858), .B2(new_n859), .ZN(G1340gat));
  OAI21_X1  g659(.A(G120gat), .B1(new_n852), .B2(new_n656), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n655), .A2(new_n249), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n861), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT119), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n865), .B(new_n861), .C1(new_n858), .C2(new_n862), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(new_n866), .ZN(G1341gat));
  NOR3_X1   g666(.A1(new_n852), .A2(new_n246), .A3(new_n755), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n856), .A2(new_n755), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n869), .A2(KEYINPUT120), .ZN(new_n870));
  AOI21_X1  g669(.A(G127gat), .B1(new_n869), .B2(KEYINPUT120), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(G1342gat));
  INV_X1    g671(.A(new_n856), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n634), .A2(G134gat), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT121), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n873), .A2(new_n877), .A3(new_n874), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT56), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(G134gat), .B1(new_n852), .B2(new_n634), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n876), .A2(KEYINPUT56), .A3(new_n878), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(G1343gat));
  NOR3_X1   g683(.A1(new_n742), .A2(new_n492), .A3(new_n692), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n854), .A2(new_n885), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n886), .A2(G141gat), .A3(new_n686), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n845), .A2(new_n685), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n684), .A2(new_n825), .A3(new_n655), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n712), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n712), .A2(new_n826), .A3(new_n845), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n755), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n657), .A2(new_n685), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n492), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT122), .B1(new_n894), .B2(KEYINPUT57), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n896), .B(new_n897), .C1(new_n849), .C2(new_n492), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n889), .A2(new_n899), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n842), .A2(new_n838), .A3(new_n836), .ZN(new_n901));
  INV_X1    g700(.A(new_n676), .ZN(new_n902));
  INV_X1    g701(.A(new_n670), .ZN(new_n903));
  AOI211_X1 g702(.A(new_n903), .B(new_n678), .C1(new_n601), .C2(new_n665), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n902), .B1(new_n904), .B2(new_n669), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n663), .B1(new_n905), .B2(new_n683), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n677), .A2(new_n680), .A3(new_n664), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n901), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n684), .A2(new_n655), .A3(KEYINPUT123), .A4(new_n825), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n900), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n634), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n546), .B1(new_n911), .B2(new_n846), .ZN(new_n912));
  OAI211_X1 g711(.A(KEYINPUT57), .B(new_n707), .C1(new_n912), .C2(new_n823), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n895), .A2(new_n898), .A3(new_n913), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n302), .A2(new_n851), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(new_n685), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n887), .B1(new_n916), .B2(new_n310), .ZN(new_n917));
  XNOR2_X1  g716(.A(KEYINPUT124), .B(KEYINPUT58), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n917), .B(new_n919), .ZN(G1344gat));
  INV_X1    g719(.A(KEYINPUT126), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n886), .A2(G148gat), .A3(new_n656), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n914), .A2(new_n655), .A3(new_n915), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n311), .A2(KEYINPUT59), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n707), .A2(KEYINPUT57), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n927), .B1(new_n892), .B2(new_n893), .ZN(new_n928));
  INV_X1    g727(.A(new_n844), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(new_n839), .A3(new_n842), .ZN(new_n930));
  OAI21_X1  g729(.A(KEYINPUT125), .B1(new_n930), .B2(new_n634), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n712), .A2(new_n845), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n931), .A2(new_n933), .A3(new_n826), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n546), .B1(new_n911), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n707), .B1(new_n935), .B2(new_n823), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n928), .B1(new_n936), .B2(new_n897), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n915), .A2(new_n655), .ZN(new_n938));
  OAI21_X1  g737(.A(G148gat), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n939), .A2(KEYINPUT59), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n921), .B(new_n923), .C1(new_n926), .C2(new_n940), .ZN(new_n941));
  AOI22_X1  g740(.A1(new_n924), .A2(new_n925), .B1(new_n939), .B2(KEYINPUT59), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT126), .B1(new_n942), .B2(new_n922), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1345gat));
  NAND2_X1  g743(.A1(new_n914), .A2(new_n915), .ZN(new_n945));
  OAI21_X1  g744(.A(G155gat), .B1(new_n945), .B2(new_n755), .ZN(new_n946));
  INV_X1    g745(.A(new_n886), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n947), .A2(new_n314), .A3(new_n546), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(G1346gat));
  NOR3_X1   g748(.A1(new_n945), .A2(new_n315), .A3(new_n634), .ZN(new_n950));
  AOI21_X1  g749(.A(G162gat), .B1(new_n947), .B2(new_n712), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n950), .A2(new_n951), .ZN(G1347gat));
  NOR4_X1   g751(.A1(new_n849), .A2(new_n689), .A3(new_n495), .A4(new_n408), .ZN(new_n953));
  AOI21_X1  g752(.A(G169gat), .B1(new_n953), .B2(new_n685), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n689), .A2(new_n408), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  NOR4_X1   g755(.A1(new_n849), .A2(new_n707), .A3(new_n704), .A4(new_n956), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n686), .A2(new_n210), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(G1348gat));
  AOI21_X1  g758(.A(G176gat), .B1(new_n953), .B2(new_n655), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n656), .A2(new_n211), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n960), .B1(new_n957), .B2(new_n961), .ZN(G1349gat));
  AOI21_X1  g761(.A(new_n219), .B1(new_n957), .B2(new_n546), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n546), .A2(new_n204), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n963), .B1(new_n953), .B2(new_n964), .ZN(new_n965));
  XOR2_X1   g764(.A(new_n965), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g765(.A(new_n231), .B1(new_n957), .B2(new_n712), .ZN(new_n967));
  XOR2_X1   g766(.A(new_n967), .B(KEYINPUT61), .Z(new_n968));
  NAND3_X1  g767(.A1(new_n953), .A2(new_n203), .A3(new_n712), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(G1351gat));
  NOR2_X1   g769(.A1(new_n849), .A2(new_n689), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n971), .A2(new_n707), .A3(new_n692), .A4(new_n302), .ZN(new_n972));
  OR2_X1    g771(.A1(new_n972), .A2(KEYINPUT127), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(KEYINPUT127), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n973), .A2(new_n685), .A3(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(G197gat), .ZN(new_n976));
  NOR3_X1   g775(.A1(new_n937), .A2(new_n742), .A3(new_n956), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n686), .A2(new_n976), .ZN(new_n978));
  AOI22_X1  g777(.A1(new_n975), .A2(new_n976), .B1(new_n977), .B2(new_n978), .ZN(G1352gat));
  NOR3_X1   g778(.A1(new_n972), .A2(G204gat), .A3(new_n656), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT62), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n977), .A2(new_n655), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n982), .B2(new_n368), .ZN(G1353gat));
  NOR2_X1   g782(.A1(new_n755), .A2(G211gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n973), .A2(new_n974), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n977), .A2(new_n546), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n986), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT63), .B1(new_n986), .B2(G211gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(G1354gat));
  INV_X1    g788(.A(G218gat), .ZN(new_n990));
  NAND4_X1  g789(.A1(new_n973), .A2(new_n990), .A3(new_n712), .A4(new_n974), .ZN(new_n991));
  AND2_X1   g790(.A1(new_n977), .A2(new_n712), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n991), .B1(new_n992), .B2(new_n990), .ZN(G1355gat));
endmodule


