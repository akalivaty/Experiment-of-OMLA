//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n623,
    new_n626, new_n627, new_n629, new_n630, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT65), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n458));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n458), .B1(G2104), .B2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR3_X1   g036(.A1(new_n461), .A2(KEYINPUT66), .A3(G2105), .ZN(new_n462));
  OAI21_X1  g037(.A(G101), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(G137), .A3(new_n459), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n459), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n466), .A2(new_n471), .ZN(G160));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(new_n461), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n459), .B1(new_n474), .B2(new_n475), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n459), .A2(G112), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n477), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT67), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  OAI211_X1 g059(.A(G126), .B(G2105), .C1(new_n467), .C2(new_n468), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n485), .A2(new_n488), .A3(KEYINPUT68), .ZN(new_n492));
  OAI211_X1 g067(.A(G138), .B(new_n459), .C1(new_n467), .C2(new_n468), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n464), .A2(new_n495), .A3(G138), .A4(new_n459), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n491), .A2(new_n492), .B1(new_n494), .B2(new_n496), .ZN(G164));
  OR2_X1    g072(.A1(KEYINPUT6), .A2(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT6), .A2(G651), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n498), .A2(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n501), .B1(new_n498), .B2(new_n499), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n504), .A2(G88), .B1(new_n505), .B2(G50), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  XOR2_X1   g084(.A(new_n509), .B(KEYINPUT69), .Z(new_n510));
  NAND2_X1  g085(.A1(new_n502), .A2(new_n503), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G62), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n508), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n507), .A2(new_n513), .ZN(G166));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT7), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n498), .A2(new_n499), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G51), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n517), .A2(G89), .ZN(new_n524));
  NAND2_X1  g099(.A1(G63), .A2(G651), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n520), .A2(new_n526), .ZN(G168));
  AOI22_X1  g102(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n508), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT70), .B(G52), .Z(new_n530));
  AND2_X1   g105(.A1(KEYINPUT6), .A2(G651), .ZN(new_n531));
  NOR2_X1   g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n522), .A2(new_n521), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n518), .A2(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n529), .A2(new_n535), .ZN(G171));
  INV_X1    g111(.A(G56), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(new_n502), .B2(new_n503), .ZN(new_n538));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g115(.A(KEYINPUT71), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n542), .B(new_n539), .C1(new_n523), .C2(new_n537), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n541), .A2(G651), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n541), .A2(new_n543), .A3(KEYINPUT72), .A4(G651), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n504), .A2(G81), .B1(new_n505), .B2(G43), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G860), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT73), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n505), .A2(new_n557), .A3(G53), .ZN(new_n558));
  OAI211_X1 g133(.A(G53), .B(G543), .C1(new_n531), .C2(new_n532), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT74), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n558), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n567), .B2(new_n508), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n523), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n571), .A2(KEYINPUT75), .A3(G651), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n568), .A2(new_n572), .B1(G91), .B2(new_n504), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n565), .A2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  INV_X1    g150(.A(G168), .ZN(G286));
  INV_X1    g151(.A(G166), .ZN(G303));
  OAI21_X1  g152(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g155(.A(KEYINPUT76), .B(G651), .C1(new_n511), .C2(G74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G49), .ZN(new_n583));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n518), .A2(new_n583), .B1(new_n533), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(G288));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  INV_X1    g163(.A(G73), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n523), .A2(new_n588), .B1(new_n589), .B2(new_n501), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G651), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(KEYINPUT77), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n588), .B1(new_n502), .B2(new_n503), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n589), .A2(new_n501), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n593), .B(G651), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n504), .A2(G86), .B1(new_n505), .B2(G48), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n592), .A2(new_n596), .A3(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n508), .ZN(new_n600));
  INV_X1    g175(.A(G47), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n518), .A2(new_n601), .B1(new_n533), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  XOR2_X1   g180(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n533), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n504), .A2(G92), .A3(new_n606), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n505), .A2(G54), .ZN(new_n611));
  INV_X1    g186(.A(G66), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(new_n502), .B2(new_n503), .ZN(new_n613));
  AND2_X1   g188(.A1(G79), .A2(G543), .ZN(new_n614));
  OAI21_X1  g189(.A(G651), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND4_X1  g190(.A1(new_n609), .A2(new_n610), .A3(new_n611), .A4(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(new_n617), .B2(G171), .ZN(G284));
  OAI21_X1  g194(.A(new_n618), .B1(new_n617), .B2(G171), .ZN(G321));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT79), .ZN(new_n622));
  INV_X1    g197(.A(G299), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(G868), .B2(new_n623), .ZN(G297));
  OAI21_X1  g199(.A(new_n622), .B1(G868), .B2(new_n623), .ZN(G280));
  INV_X1    g200(.A(new_n616), .ZN(new_n626));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n549), .A2(new_n617), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n616), .A2(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n617), .B2(new_n630), .ZN(G323));
  XNOR2_X1  g206(.A(KEYINPUT80), .B(KEYINPUT11), .ZN(new_n632));
  XNOR2_X1  g207(.A(G323), .B(new_n632), .ZN(G282));
  OR2_X1    g208(.A1(new_n460), .A2(new_n462), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(new_n464), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  INV_X1    g212(.A(G2100), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n476), .A2(G135), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n478), .A2(G123), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n459), .A2(G111), .ZN(new_n643));
  OAI21_X1  g218(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n641), .B(new_n642), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2096), .Z(new_n646));
  NAND3_X1  g221(.A1(new_n639), .A2(new_n640), .A3(new_n646), .ZN(G156));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT83), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2427), .B(G2430), .Z(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT82), .B(KEYINPUT14), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n659), .B(new_n660), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  OR3_X1    g237(.A1(new_n657), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n662), .B1(new_n657), .B2(new_n658), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n667), .A2(G14), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n663), .A2(new_n666), .ZN(new_n669));
  AND3_X1   g244(.A1(new_n669), .A2(KEYINPUT84), .A3(new_n664), .ZN(new_n670));
  AOI21_X1  g245(.A(KEYINPUT84), .B1(new_n669), .B2(new_n664), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n668), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G401));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2072), .B(G2078), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT87), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT88), .B(G2100), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n677), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT86), .B(KEYINPUT17), .Z(new_n685));
  NAND2_X1  g260(.A1(new_n676), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n674), .A2(new_n675), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G2096), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n683), .A2(new_n689), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(G227));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  XNOR2_X1  g268(.A(G1971), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT19), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1956), .B(G2474), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT89), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1961), .B(G1966), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(new_n695), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n698), .A2(new_n699), .ZN(new_n702));
  MUX2_X1   g277(.A(new_n695), .B(new_n701), .S(new_n702), .Z(new_n703));
  NOR2_X1   g278(.A1(new_n700), .A2(new_n695), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT20), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n703), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n707), .B1(new_n703), .B2(new_n706), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n693), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(new_n693), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n712), .A2(new_n713), .A3(new_n708), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(G1981), .B(G1986), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n711), .A2(new_n714), .A3(new_n716), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(G229));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G35), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G162), .B2(new_n722), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT29), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G2090), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G20), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT23), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n623), .B2(new_n727), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(G1956), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT100), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n727), .A2(G19), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT92), .Z(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n549), .B2(G16), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1341), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT93), .B(KEYINPUT25), .Z(new_n738));
  NAND3_X1  g313(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n476), .A2(G139), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(new_n459), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(new_n722), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n722), .B2(G33), .ZN(new_n747));
  INV_X1    g322(.A(G2072), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT94), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n722), .A2(G27), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G164), .B2(new_n722), .ZN(new_n752));
  INV_X1    g327(.A(G2078), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G168), .A2(new_n727), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n727), .B2(G21), .ZN(new_n756));
  INV_X1    g331(.A(G1966), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT98), .Z(new_n759));
  NAND3_X1  g334(.A1(new_n750), .A2(new_n754), .A3(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G2084), .ZN(new_n761));
  NAND2_X1  g336(.A1(G160), .A2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT95), .B(KEYINPUT24), .ZN(new_n763));
  INV_X1    g338(.A(G34), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(G29), .B1(new_n763), .B2(new_n764), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT96), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n767), .B2(new_n766), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n762), .A2(new_n769), .ZN(new_n770));
  OAI22_X1  g345(.A1(new_n747), .A2(new_n748), .B1(new_n761), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n761), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n727), .A2(G5), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G171), .B2(new_n727), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n772), .B1(new_n774), .B2(G1961), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n626), .A2(G16), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G4), .B2(G16), .ZN(new_n778));
  INV_X1    g353(.A(G1348), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G28), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n781), .A2(KEYINPUT30), .ZN(new_n782));
  AOI21_X1  g357(.A(G29), .B1(new_n781), .B2(KEYINPUT30), .ZN(new_n783));
  OR2_X1    g358(.A1(KEYINPUT31), .A2(G11), .ZN(new_n784));
  NAND2_X1  g359(.A1(KEYINPUT31), .A2(G11), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n782), .A2(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n645), .B2(new_n722), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n756), .B2(new_n757), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n778), .A2(new_n779), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n722), .A2(G26), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT28), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n476), .A2(G140), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n478), .A2(G128), .ZN(new_n793));
  OR2_X1    g368(.A1(G104), .A2(G2105), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n794), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n792), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n791), .B1(new_n797), .B2(new_n722), .ZN(new_n798));
  INV_X1    g373(.A(G2067), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  AND4_X1   g375(.A1(new_n780), .A2(new_n788), .A3(new_n789), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n774), .A2(G1961), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT99), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n776), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n722), .A2(G32), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n634), .A2(G105), .B1(G141), .B2(new_n476), .ZN(new_n806));
  NAND3_X1  g381(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT26), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G129), .B2(new_n478), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n805), .B1(new_n811), .B2(new_n722), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT97), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT27), .B(G1996), .Z(new_n814));
  XOR2_X1   g389(.A(new_n813), .B(new_n814), .Z(new_n815));
  NOR2_X1   g390(.A1(new_n725), .A2(G2090), .ZN(new_n816));
  NOR4_X1   g391(.A1(new_n760), .A2(new_n804), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n733), .A2(new_n737), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n727), .A2(G23), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n585), .B1(new_n580), .B2(new_n581), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(new_n727), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT33), .B(G1976), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n821), .B(new_n822), .Z(new_n823));
  OR2_X1    g398(.A1(G6), .A2(G16), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G305), .B2(new_n727), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT32), .B(G1981), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n727), .A2(G22), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(G166), .B2(new_n727), .ZN(new_n831));
  INV_X1    g406(.A(G1971), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n829), .B1(new_n833), .B2(KEYINPUT91), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n828), .B(new_n834), .C1(KEYINPUT91), .C2(new_n833), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n835), .A2(KEYINPUT34), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT36), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(KEYINPUT34), .ZN(new_n838));
  NOR2_X1   g413(.A1(G16), .A2(G24), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n604), .B(KEYINPUT90), .Z(new_n840));
  AOI21_X1  g415(.A(new_n839), .B1(new_n840), .B2(G16), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G1986), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n722), .A2(G25), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n476), .A2(G131), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n478), .A2(G119), .ZN(new_n845));
  OR2_X1    g420(.A1(G95), .A2(G2105), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n846), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n844), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n843), .B1(new_n849), .B2(new_n722), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT35), .B(G1991), .Z(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n850), .B(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n842), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n836), .A2(new_n837), .A3(new_n838), .A4(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n836), .A2(new_n838), .A3(new_n854), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(KEYINPUT36), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n818), .B1(new_n855), .B2(new_n857), .ZN(G311));
  INV_X1    g433(.A(new_n818), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n855), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(G150));
  INV_X1    g436(.A(G67), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(new_n502), .B2(new_n503), .ZN(new_n863));
  NAND2_X1  g438(.A1(G80), .A2(G543), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(KEYINPUT102), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n867), .B(new_n864), .C1(new_n523), .C2(new_n862), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n866), .A2(G651), .A3(new_n868), .ZN(new_n869));
  AOI22_X1  g444(.A1(new_n504), .A2(G93), .B1(new_n505), .B2(G55), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n869), .A2(new_n870), .A3(KEYINPUT103), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n549), .A2(new_n873), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n546), .A2(new_n871), .A3(new_n547), .A4(new_n548), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n869), .A2(KEYINPUT103), .A3(new_n870), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT103), .B1(new_n869), .B2(new_n870), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n874), .B1(new_n881), .B2(new_n549), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n626), .A2(G559), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n887), .A2(KEYINPUT39), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(KEYINPUT39), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n550), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n881), .A2(new_n550), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT37), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(G145));
  NAND2_X1  g468(.A1(new_n476), .A2(G142), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT106), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT107), .ZN(new_n896));
  OAI21_X1  g471(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n897));
  INV_X1    g472(.A(G118), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n897), .B1(new_n898), .B2(G2105), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n899), .B1(G130), .B2(new_n478), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n895), .A2(new_n896), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n636), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n896), .B1(new_n895), .B2(new_n900), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n895), .A2(new_n900), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT107), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n636), .B1(new_n907), .B2(new_n901), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n849), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n903), .B1(new_n902), .B2(new_n904), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n907), .A2(new_n636), .A3(new_n901), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n848), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n745), .A2(KEYINPUT105), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n489), .B1(new_n494), .B2(new_n496), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n797), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n494), .A2(new_n496), .ZN(new_n917));
  INV_X1    g492(.A(new_n489), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n796), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n810), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n811), .A2(new_n916), .A3(new_n920), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n914), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n745), .A2(KEYINPUT105), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n914), .A2(new_n922), .A3(new_n925), .A4(new_n923), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n913), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n909), .A2(new_n927), .A3(new_n912), .A4(new_n928), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(G160), .B(new_n645), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(new_n483), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(G37), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n930), .A2(new_n934), .A3(new_n931), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(KEYINPUT108), .A3(new_n937), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n940), .A2(new_n941), .A3(KEYINPUT40), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT40), .B1(new_n940), .B2(new_n941), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(G395));
  XOR2_X1   g519(.A(new_n883), .B(new_n630), .Z(new_n945));
  INV_X1    g520(.A(KEYINPUT41), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n565), .A2(new_n626), .A3(new_n573), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n626), .B1(new_n565), .B2(new_n573), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(G299), .A2(new_n616), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n565), .A2(new_n626), .A3(new_n573), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(KEYINPUT41), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n945), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n945), .B1(new_n948), .B2(new_n947), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n604), .A2(KEYINPUT109), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n604), .A2(KEYINPUT109), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n820), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n957), .A2(G288), .A3(new_n958), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(G305), .B(G166), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n963), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n965), .A2(new_n961), .A3(new_n960), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n967), .B(KEYINPUT42), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n955), .A2(new_n956), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n968), .B1(new_n955), .B2(new_n956), .ZN(new_n970));
  OAI21_X1  g545(.A(G868), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(G868), .B2(new_n881), .ZN(G295));
  OAI21_X1  g547(.A(new_n971), .B1(G868), .B2(new_n881), .ZN(G331));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n975));
  XNOR2_X1  g550(.A(G171), .B(G168), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n878), .B2(new_n882), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n549), .A2(new_n873), .A3(new_n875), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT104), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n980), .A2(new_n877), .A3(new_n876), .A4(new_n976), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n954), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n947), .A2(new_n948), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n978), .A2(new_n984), .A3(new_n981), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(G37), .B1(new_n986), .B2(new_n967), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n978), .A2(new_n984), .A3(new_n981), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n953), .B1(new_n978), .B2(new_n981), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n964), .A2(new_n966), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NOR4_X1   g568(.A1(new_n989), .A2(new_n990), .A3(new_n967), .A4(KEYINPUT110), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n975), .B(new_n987), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n983), .A2(new_n992), .A3(new_n985), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT110), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n983), .A2(new_n992), .A3(new_n988), .A4(new_n985), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n975), .B1(new_n1000), .B2(new_n987), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n974), .B1(new_n996), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n987), .B1(new_n993), .B2(new_n994), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT43), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(KEYINPUT44), .A3(new_n995), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1002), .A2(new_n1005), .ZN(G397));
  AOI21_X1  g581(.A(G1384), .B1(new_n917), .B2(new_n918), .ZN(new_n1007));
  INV_X1    g582(.A(G125), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(new_n474), .B2(new_n475), .ZN(new_n1009));
  INV_X1    g584(.A(new_n470), .ZN(new_n1010));
  OAI21_X1  g585(.A(G2105), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1011), .A2(G40), .A3(new_n463), .A4(new_n465), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n1007), .A2(KEYINPUT45), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1996), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT112), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT46), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1013), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n796), .B(new_n799), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1018), .B1(new_n1019), .B2(new_n811), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1017), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT126), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1017), .A2(KEYINPUT126), .A3(new_n1021), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(KEYINPUT47), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1019), .B1(new_n1014), .B2(new_n811), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n1013), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n1016), .B2(new_n810), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n848), .B(new_n852), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1029), .B1(new_n1013), .B2(new_n1030), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1018), .A2(G1986), .A3(G290), .ZN(new_n1032));
  XOR2_X1   g607(.A(new_n1032), .B(KEYINPUT48), .Z(new_n1033));
  NAND2_X1  g608(.A1(new_n849), .A2(new_n851), .ZN(new_n1034));
  OAI22_X1  g609(.A1(new_n1029), .A2(new_n1034), .B1(G2067), .B2(new_n796), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n1031), .A2(new_n1033), .B1(new_n1035), .B2(new_n1013), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1026), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT47), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1981), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n592), .A2(new_n1040), .A3(new_n596), .A4(new_n597), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n597), .A2(new_n596), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n593), .B1(new_n590), .B2(G651), .ZN(new_n1044));
  OAI21_X1  g619(.A(G1981), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(new_n1041), .A3(KEYINPUT49), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT114), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1045), .A2(new_n1041), .A3(new_n1048), .A4(KEYINPUT49), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT49), .B1(new_n1045), .B2(new_n1041), .ZN(new_n1051));
  INV_X1    g626(.A(G8), .ZN(new_n1052));
  INV_X1    g627(.A(G40), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n466), .A2(new_n1053), .A3(new_n471), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1052), .B1(new_n1007), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1051), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1050), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(G288), .A2(G1976), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1042), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT113), .B1(new_n820), .B2(G1976), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n1055), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1007), .A2(new_n1054), .ZN(new_n1064));
  INV_X1    g639(.A(G1976), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1064), .A2(G8), .A3(new_n1065), .A4(G288), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1062), .A2(new_n1063), .A3(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n820), .A2(G1976), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1061), .B(new_n1055), .C1(new_n1068), .C2(KEYINPUT52), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1058), .A2(new_n1070), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n485), .A2(new_n488), .A3(KEYINPUT68), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT68), .B1(new_n485), .B2(new_n488), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n917), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1384), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT45), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT45), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(G1384), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1054), .B1(new_n915), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n832), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1082));
  INV_X1    g657(.A(G2090), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT50), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1012), .B1(new_n1007), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1081), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1088));
  NAND3_X1  g663(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1087), .B(G8), .C1(new_n1088), .C2(new_n1090), .ZN(new_n1091));
  OAI22_X1  g666(.A1(new_n1060), .A2(new_n1056), .B1(new_n1071), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT63), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1050), .A2(new_n1057), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1074), .A2(new_n1084), .A3(new_n1075), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT50), .B1(new_n915), .B2(G1384), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1095), .A2(new_n1083), .A3(new_n1096), .A4(new_n1054), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1081), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(G8), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1090), .A2(new_n1088), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1094), .A2(new_n1101), .A3(new_n1091), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n919), .A2(new_n1075), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1012), .B1(new_n1103), .B2(new_n1077), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1074), .A2(KEYINPUT115), .A3(new_n1078), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT115), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(G164), .B2(new_n1079), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1104), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n757), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n919), .A2(new_n1084), .A3(new_n1075), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n1054), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1084), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n761), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1109), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1115), .A2(G8), .A3(G168), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1093), .B1(new_n1102), .B2(new_n1116), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1108), .A2(new_n757), .B1(new_n1113), .B2(new_n761), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1118), .A2(new_n1052), .A3(G286), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1087), .A2(G8), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1093), .B1(new_n1120), .B2(new_n1100), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1119), .A2(new_n1121), .A3(new_n1091), .A4(new_n1094), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1092), .B1(new_n1117), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1076), .A2(new_n1080), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT53), .B1(new_n1124), .B2(new_n753), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT53), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1126), .A2(G2078), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1104), .A2(new_n1107), .A3(new_n1127), .A4(new_n1105), .ZN(new_n1128));
  INV_X1    g703(.A(G1961), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT120), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1128), .A2(new_n1130), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1125), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1135), .A2(G301), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1102), .ZN(new_n1137));
  NAND2_X1  g712(.A1(G286), .A2(G8), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1118), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT51), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(G8), .B(new_n1143), .C1(new_n1115), .C2(G286), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1138), .B(new_n1142), .C1(new_n1118), .C2(new_n1052), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1139), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1136), .B(new_n1137), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1148));
  AOI211_X1 g723(.A(KEYINPUT62), .B(new_n1139), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1123), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1007), .A2(new_n1054), .A3(KEYINPUT117), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT117), .B1(new_n1007), .B2(new_n1054), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n799), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1154), .B(new_n616), .C1(G1348), .C2(new_n1113), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT117), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1064), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(G2067), .B1(new_n1157), .B2(new_n1151), .ZN(new_n1158));
  AOI21_X1  g733(.A(G1348), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n626), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1155), .A2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n616), .A2(KEYINPUT60), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1161), .A2(KEYINPUT60), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT57), .B1(new_n558), .B2(new_n560), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n573), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT57), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1166), .B1(new_n623), .B2(new_n1167), .ZN(new_n1168));
  XOR2_X1   g743(.A(KEYINPUT116), .B(G1956), .Z(new_n1169));
  INV_X1    g744(.A(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1012), .B1(new_n1103), .B2(KEYINPUT50), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1170), .B1(new_n1171), .B2(new_n1095), .ZN(new_n1172));
  XOR2_X1   g747(.A(KEYINPUT56), .B(G2072), .Z(new_n1173));
  NOR3_X1   g748(.A1(new_n1076), .A2(new_n1080), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1168), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1174), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1095), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1096), .A2(new_n1054), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1169), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  AOI22_X1  g754(.A1(G299), .A2(KEYINPUT57), .B1(new_n573), .B2(new_n1165), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1176), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1175), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1176), .A2(new_n1179), .A3(KEYINPUT61), .A4(new_n1180), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n549), .ZN(new_n1186));
  XNOR2_X1  g761(.A(KEYINPUT58), .B(G1341), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1152), .A2(new_n1153), .A3(new_n1187), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1076), .A2(new_n1080), .A3(G1996), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1186), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT59), .ZN(new_n1192));
  OAI211_X1 g767(.A(new_n1192), .B(new_n1186), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1164), .A2(new_n1185), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1180), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n1196), .A2(KEYINPUT118), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1160), .B1(new_n1196), .B2(KEYINPUT118), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1181), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1012), .B1(new_n919), .B2(new_n1078), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n491), .A2(new_n492), .ZN(new_n1202));
  AOI21_X1  g777(.A(G1384), .B1(new_n1202), .B2(new_n917), .ZN(new_n1203));
  OAI211_X1 g778(.A(new_n1201), .B(new_n753), .C1(new_n1203), .C2(KEYINPUT45), .ZN(new_n1204));
  AOI211_X1 g779(.A(new_n1126), .B(G2078), .C1(new_n919), .C2(new_n1078), .ZN(new_n1205));
  AOI22_X1  g780(.A1(new_n1204), .A2(new_n1126), .B1(new_n1104), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT121), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1130), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1209), .A2(KEYINPUT121), .A3(new_n1129), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1206), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n1212));
  AOI21_X1  g787(.A(G301), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1213), .B1(new_n1212), .B2(new_n1211), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n1125), .A2(G171), .ZN(new_n1215));
  INV_X1    g790(.A(new_n1134), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1133), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1215), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1218), .A2(KEYINPUT124), .ZN(new_n1219));
  INV_X1    g794(.A(KEYINPUT124), .ZN(new_n1220));
  OAI211_X1 g795(.A(new_n1220), .B(new_n1215), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1221));
  NAND4_X1  g796(.A1(new_n1214), .A2(KEYINPUT54), .A3(new_n1219), .A4(new_n1221), .ZN(new_n1222));
  NOR2_X1   g797(.A1(new_n1146), .A2(new_n1102), .ZN(new_n1223));
  AND3_X1   g798(.A1(new_n1200), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  NAND4_X1  g799(.A1(new_n1206), .A2(new_n1208), .A3(G301), .A4(new_n1210), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1225), .A2(KEYINPUT122), .ZN(new_n1226));
  AOI21_X1  g801(.A(KEYINPUT121), .B1(new_n1209), .B2(new_n1129), .ZN(new_n1227));
  AOI211_X1 g802(.A(new_n1207), .B(G1961), .C1(new_n1082), .C2(new_n1085), .ZN(new_n1228));
  NOR2_X1   g803(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g804(.A(KEYINPUT122), .ZN(new_n1230));
  NAND4_X1  g805(.A1(new_n1229), .A2(new_n1230), .A3(G301), .A4(new_n1206), .ZN(new_n1231));
  OAI211_X1 g806(.A(new_n1226), .B(new_n1231), .C1(new_n1135), .C2(G301), .ZN(new_n1232));
  INV_X1    g807(.A(KEYINPUT54), .ZN(new_n1233));
  AND3_X1   g808(.A1(new_n1232), .A2(KEYINPUT123), .A3(new_n1233), .ZN(new_n1234));
  AOI21_X1  g809(.A(KEYINPUT123), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1235));
  NOR2_X1   g810(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g811(.A(new_n1150), .B1(new_n1224), .B2(new_n1236), .ZN(new_n1237));
  AND2_X1   g812(.A1(G290), .A2(G1986), .ZN(new_n1238));
  AOI21_X1  g813(.A(new_n1032), .B1(new_n1013), .B2(new_n1238), .ZN(new_n1239));
  XOR2_X1   g814(.A(new_n1239), .B(KEYINPUT111), .Z(new_n1240));
  NAND2_X1  g815(.A1(new_n1240), .A2(new_n1031), .ZN(new_n1241));
  OAI21_X1  g816(.A(new_n1039), .B1(new_n1237), .B2(new_n1241), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g817(.A1(new_n690), .A2(new_n456), .A3(new_n691), .ZN(new_n1244));
  INV_X1    g818(.A(KEYINPUT127), .ZN(new_n1245));
  NAND2_X1  g819(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND4_X1  g820(.A1(new_n690), .A2(KEYINPUT127), .A3(new_n456), .A4(new_n691), .ZN(new_n1247));
  NAND2_X1  g821(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  AND3_X1   g822(.A1(new_n720), .A2(new_n672), .A3(new_n1248), .ZN(new_n1249));
  AOI21_X1  g823(.A(KEYINPUT108), .B1(new_n936), .B2(new_n937), .ZN(new_n1250));
  INV_X1    g824(.A(new_n931), .ZN(new_n1251));
  AOI22_X1  g825(.A1(new_n909), .A2(new_n912), .B1(new_n927), .B2(new_n928), .ZN(new_n1252));
  OAI21_X1  g826(.A(new_n935), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g827(.A(G37), .ZN(new_n1254));
  AND4_X1   g828(.A1(KEYINPUT108), .A2(new_n1253), .A3(new_n1254), .A4(new_n937), .ZN(new_n1255));
  OAI21_X1  g829(.A(new_n1249), .B1(new_n1250), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g830(.A(new_n1256), .B1(new_n1004), .B2(new_n995), .ZN(G308));
  OAI221_X1 g831(.A(new_n1249), .B1(new_n1250), .B2(new_n1255), .C1(new_n996), .C2(new_n1001), .ZN(G225));
endmodule


