//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976;
  INV_X1    g000(.A(KEYINPUT78), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT76), .ZN(new_n203));
  INV_X1    g002(.A(G190gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT66), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT66), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G190gat), .ZN(new_n207));
  INV_X1    g006(.A(G183gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT27), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT27), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G183gat), .ZN(new_n211));
  NAND4_X1  g010(.A1(new_n205), .A2(new_n207), .A3(new_n209), .A4(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT28), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G190gat), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT28), .B1(new_n210), .B2(G183gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT67), .B1(new_n210), .B2(G183gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(new_n208), .A3(KEYINPUT27), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n215), .A2(new_n216), .A3(new_n217), .A4(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n213), .A2(new_n214), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT26), .ZN(new_n222));
  INV_X1    g021(.A(G169gat), .ZN(new_n223));
  INV_X1    g022(.A(G176gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT69), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT68), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n225), .A2(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NOR3_X1   g030(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(KEYINPUT69), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n227), .A2(new_n228), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n229), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n221), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT23), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(new_n223), .A3(new_n224), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n231), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n214), .A2(KEYINPUT24), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT24), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(G183gat), .A3(G190gat), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(G183gat), .A2(G190gat), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n240), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n247));
  INV_X1    g046(.A(new_n239), .ZN(new_n248));
  NOR3_X1   g047(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n230), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(KEYINPUT25), .A3(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n243), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n246), .A2(new_n247), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n203), .B1(new_n236), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n238), .A2(new_n239), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n253), .A2(KEYINPUT25), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n258), .A2(new_n261), .A3(new_n252), .A4(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n230), .B1(new_n248), .B2(new_n249), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n245), .B1(new_n241), .B2(new_n243), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n247), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n229), .A2(new_n233), .A3(new_n234), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n268), .A2(new_n214), .A3(new_n213), .A4(new_n220), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n269), .A3(KEYINPUT76), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT29), .B1(new_n260), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G226gat), .A2(G233gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n202), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G197gat), .B(G204gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT22), .ZN(new_n276));
  INV_X1    g075(.A(G211gat), .ZN(new_n277));
  INV_X1    g076(.A(G218gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G211gat), .B(G218gat), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(new_n275), .A3(new_n279), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT29), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n267), .A2(new_n269), .A3(KEYINPUT76), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT76), .B1(new_n267), .B2(new_n269), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(KEYINPUT78), .A3(new_n272), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n267), .A2(new_n269), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n272), .B(KEYINPUT75), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n274), .A2(new_n286), .A3(new_n291), .A4(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G8gat), .B(G36gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(G64gat), .B(G92gat), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n296), .B(new_n297), .Z(new_n298));
  INV_X1    g097(.A(KEYINPUT77), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n273), .B1(new_n288), .B2(new_n289), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n293), .B1(new_n292), .B2(new_n287), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n299), .B1(new_n303), .B2(new_n285), .ZN(new_n304));
  AOI211_X1 g103(.A(KEYINPUT77), .B(new_n286), .C1(new_n300), .C2(new_n302), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n295), .B(new_n298), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT79), .B(KEYINPUT30), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  XOR2_X1   g107(.A(G1gat), .B(G29gat), .Z(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G57gat), .B(G85gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT4), .ZN(new_n314));
  XOR2_X1   g113(.A(G127gat), .B(G134gat), .Z(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT71), .ZN(new_n316));
  XNOR2_X1  g115(.A(G113gat), .B(G120gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(KEYINPUT1), .ZN(new_n318));
  XNOR2_X1  g117(.A(G127gat), .B(G134gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT71), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n316), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT1), .ZN(new_n323));
  INV_X1    g122(.A(G113gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n324), .A2(G120gat), .ZN(new_n325));
  INV_X1    g124(.A(G120gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(G113gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n323), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G127gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n329), .A2(KEYINPUT70), .A3(G134gat), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n328), .B(new_n330), .C1(KEYINPUT70), .C2(new_n315), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n322), .A2(new_n331), .ZN(new_n332));
  XOR2_X1   g131(.A(G141gat), .B(G148gat), .Z(new_n333));
  INV_X1    g132(.A(G155gat), .ZN(new_n334));
  INV_X1    g133(.A(G162gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(KEYINPUT2), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n333), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G141gat), .B(G148gat), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n337), .B(new_n336), .C1(new_n341), .C2(KEYINPUT2), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n314), .B1(new_n332), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(KEYINPUT3), .ZN(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT80), .B(KEYINPUT3), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n340), .A2(new_n342), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n332), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G225gat), .A2(G233gat), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n340), .A2(new_n342), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n350), .A2(KEYINPUT4), .A3(new_n331), .A4(new_n322), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n344), .A2(new_n348), .A3(new_n349), .A4(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT5), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n332), .A2(new_n343), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n350), .A2(new_n331), .A3(new_n322), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n349), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n352), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n352), .A2(new_n353), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n313), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT6), .ZN(new_n361));
  INV_X1    g160(.A(new_n313), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n357), .B(new_n362), .C1(new_n353), .C2(new_n352), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n360), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n358), .A2(new_n359), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n365), .A2(KEYINPUT6), .A3(new_n362), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n295), .B1(new_n304), .B2(new_n305), .ZN(new_n368));
  INV_X1    g167(.A(new_n298), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n260), .A2(new_n270), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n301), .B1(new_n371), .B2(new_n273), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT77), .B1(new_n372), .B2(new_n286), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n303), .A2(new_n299), .A3(new_n285), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n298), .A2(KEYINPUT30), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n295), .A3(new_n376), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n308), .A2(new_n367), .A3(new_n370), .A4(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT34), .ZN(new_n379));
  INV_X1    g178(.A(new_n332), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n292), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n267), .A2(new_n269), .A3(new_n332), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G227gat), .A2(G233gat), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n379), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n267), .A2(new_n269), .A3(new_n332), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n332), .B1(new_n267), .B2(new_n269), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n379), .B(new_n384), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n384), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n381), .A2(new_n391), .A3(new_n382), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT32), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT72), .B(KEYINPUT33), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  XOR2_X1   g194(.A(G15gat), .B(G43gat), .Z(new_n396));
  XNOR2_X1  g195(.A(G71gat), .B(G99gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n393), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n398), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n392), .B(KEYINPUT32), .C1(new_n394), .C2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  OAI211_X1 g201(.A(KEYINPUT73), .B(new_n390), .C1(new_n399), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n383), .A2(new_n384), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT34), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(KEYINPUT73), .A3(new_n388), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT73), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n407), .B1(new_n385), .B2(new_n389), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n395), .A3(new_n398), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n406), .A2(new_n408), .A3(new_n401), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n403), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n347), .A2(new_n287), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n285), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT29), .B1(new_n283), .B2(new_n284), .ZN(new_n414));
  INV_X1    g213(.A(new_n346), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n343), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(G228gat), .A2(G233gat), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n412), .B2(new_n285), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n343), .B1(new_n414), .B2(KEYINPUT3), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n417), .A2(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G22gat), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT83), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT83), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n419), .A2(new_n420), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  AOI22_X1  g225(.A1(new_n413), .A2(new_n416), .B1(G228gat), .B2(G233gat), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n424), .B(G22gat), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G78gat), .B(G106gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT31), .B(G50gat), .ZN(new_n431));
  XOR2_X1   g230(.A(new_n430), .B(new_n431), .Z(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT82), .B(G22gat), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n432), .B1(new_n421), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n433), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n435), .B1(new_n426), .B2(new_n427), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n433), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n429), .A2(new_n434), .B1(new_n438), .B2(new_n432), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n411), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT35), .B1(new_n378), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT87), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(KEYINPUT87), .B(KEYINPUT35), .C1(new_n378), .C2(new_n441), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n308), .A2(new_n370), .A3(new_n377), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT84), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n375), .A2(new_n295), .A3(new_n376), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n298), .B1(new_n375), .B2(new_n295), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT84), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(new_n451), .A3(new_n308), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n441), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n367), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n454), .A2(KEYINPUT35), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n444), .A2(new_n445), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT74), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n403), .A2(new_n410), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT36), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n403), .A2(new_n410), .A3(new_n457), .A4(KEYINPUT36), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n378), .A2(new_n439), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n306), .A2(new_n366), .A3(new_n364), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n368), .A2(KEYINPUT37), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n298), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n467), .B1(new_n449), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n466), .B1(new_n470), .B2(KEYINPUT38), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n290), .A2(new_n272), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n472), .A2(new_n202), .B1(new_n292), .B2(new_n293), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n286), .B1(new_n473), .B2(new_n291), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT86), .ZN(new_n475));
  OAI22_X1  g274(.A1(new_n474), .A2(new_n475), .B1(new_n285), .B2(new_n303), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n274), .A2(new_n291), .A3(new_n294), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n285), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n478), .A2(KEYINPUT86), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT37), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n469), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT38), .B1(new_n370), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n439), .B1(new_n471), .B2(new_n483), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n344), .A2(new_n351), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n349), .B1(new_n485), .B2(new_n348), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT39), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n354), .A2(new_n355), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n487), .B1(new_n488), .B2(new_n349), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n486), .B1(KEYINPUT85), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(KEYINPUT85), .B2(new_n489), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n362), .B1(new_n486), .B2(new_n487), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n491), .A2(KEYINPUT40), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT40), .B1(new_n491), .B2(new_n492), .ZN(new_n494));
  INV_X1    g293(.A(new_n363), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n447), .A2(new_n452), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n465), .B1(new_n484), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT88), .B1(new_n456), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n469), .B1(new_n368), .B2(new_n369), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n468), .B1(new_n375), .B2(new_n295), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT38), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n466), .ZN(new_n503));
  INV_X1    g302(.A(new_n479), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n478), .A2(KEYINPUT86), .B1(new_n286), .B2(new_n372), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n468), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT38), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n507), .B1(new_n449), .B2(new_n469), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n502), .B(new_n503), .C1(new_n506), .C2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n497), .A2(new_n509), .A3(new_n440), .ZN(new_n510));
  INV_X1    g309(.A(new_n465), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n439), .B1(new_n403), .B2(new_n410), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n451), .B1(new_n450), .B2(new_n308), .ZN(new_n514));
  AND4_X1   g313(.A1(new_n451), .A2(new_n308), .A3(new_n370), .A4(new_n377), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n513), .B(new_n455), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n445), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n450), .A2(new_n513), .A3(new_n367), .A4(new_n308), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT87), .B1(new_n518), .B2(KEYINPUT35), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n516), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT88), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n512), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(G36gat), .ZN(new_n523));
  AND2_X1   g322(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(G29gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n527), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n529), .A2(KEYINPUT15), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(KEYINPUT15), .ZN(new_n531));
  XNOR2_X1  g330(.A(G43gat), .B(G50gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n531), .A2(new_n532), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT17), .ZN(new_n536));
  XNOR2_X1  g335(.A(G15gat), .B(G22gat), .ZN(new_n537));
  INV_X1    g336(.A(G1gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT16), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(G1gat), .B2(new_n537), .ZN(new_n541));
  INV_X1    g340(.A(G8gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n536), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G229gat), .A2(G233gat), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n543), .A2(KEYINPUT90), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n543), .A2(KEYINPUT90), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n535), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT18), .ZN(new_n550));
  OR3_X1    g349(.A1(new_n546), .A2(new_n547), .A3(new_n535), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n548), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n545), .B(KEYINPUT13), .Z(new_n553));
  AOI22_X1  g352(.A1(new_n549), .A2(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n544), .A2(KEYINPUT18), .A3(new_n545), .A4(new_n548), .ZN(new_n555));
  XNOR2_X1  g354(.A(G113gat), .B(G141gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G169gat), .B(G197gat), .Z(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT12), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n554), .A2(new_n555), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n561), .B1(new_n554), .B2(new_n555), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G71gat), .A2(G78gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(G71gat), .A2(G78gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT91), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n570), .B1(new_n569), .B2(new_n568), .ZN(new_n571));
  INV_X1    g370(.A(G57gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(G64gat), .ZN(new_n573));
  INV_X1    g372(.A(G64gat), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n574), .A2(G57gat), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT9), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n567), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT92), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n580), .A2(KEYINPUT93), .A3(G57gat), .A4(G64gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT93), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n574), .B1(new_n582), .B2(new_n572), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n572), .A2(KEYINPUT92), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n579), .A2(new_n581), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n577), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT21), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(new_n329), .ZN(new_n591));
  INV_X1    g390(.A(new_n586), .ZN(new_n592));
  AOI211_X1 g391(.A(new_n547), .B(new_n546), .C1(KEYINPUT21), .C2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n591), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G183gat), .B(G211gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT94), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(new_n334), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n596), .B(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n594), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(G85gat), .ZN(new_n604));
  INV_X1    g403(.A(G92gat), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT96), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT96), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n607), .A2(G85gat), .A3(G92gat), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(KEYINPUT7), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT7), .ZN(new_n610));
  OAI211_X1 g409(.A(KEYINPUT96), .B(new_n610), .C1(new_n604), .C2(new_n605), .ZN(new_n611));
  NAND2_X1  g410(.A1(G99gat), .A2(G106gat), .ZN(new_n612));
  AOI22_X1  g411(.A1(KEYINPUT8), .A2(new_n612), .B1(new_n604), .B2(new_n605), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n609), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G99gat), .B(G106gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n536), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g417(.A1(G232gat), .A2(G233gat), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n535), .A2(new_n616), .B1(KEYINPUT41), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G190gat), .B(G218gat), .Z(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n619), .A2(KEYINPUT41), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT95), .ZN(new_n625));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n622), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n618), .A2(new_n628), .A3(new_n620), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n623), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n627), .B1(new_n623), .B2(new_n629), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n603), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n592), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  OR3_X1    g434(.A1(new_n634), .A2(KEYINPUT97), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n617), .A2(new_n586), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n637), .A2(new_n635), .A3(new_n634), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT97), .B1(new_n634), .B2(new_n635), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT98), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n637), .A2(new_n634), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n642), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G120gat), .B(G148gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(G176gat), .B(G204gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n647), .B(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n633), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n499), .A2(new_n522), .A3(new_n566), .A4(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(new_n367), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(new_n538), .ZN(G1324gat));
  NAND2_X1  g454(.A1(new_n447), .A2(new_n452), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT16), .B(G8gat), .Z(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(new_n542), .B2(new_n657), .ZN(new_n660));
  MUX2_X1   g459(.A(new_n659), .B(new_n660), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g460(.A(G15gat), .B1(new_n653), .B2(new_n463), .ZN(new_n662));
  INV_X1    g461(.A(new_n411), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n663), .A2(G15gat), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n662), .B1(new_n653), .B2(new_n664), .ZN(G1326gat));
  NOR2_X1   g464(.A1(new_n653), .A2(new_n440), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT43), .B(G22gat), .Z(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1327gat));
  NOR3_X1   g467(.A1(new_n603), .A2(new_n632), .A3(new_n651), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n499), .A2(new_n522), .A3(new_n566), .A4(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n671), .A2(new_n527), .A3(new_n454), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT45), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n603), .B(KEYINPUT99), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n651), .B(KEYINPUT100), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(new_n566), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT101), .ZN(new_n677));
  INV_X1    g476(.A(new_n632), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n499), .A2(new_n522), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT44), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n516), .B(new_n681), .C1(new_n517), .C2(new_n519), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n444), .A2(new_n445), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n681), .B1(new_n684), .B2(new_n516), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n512), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(new_n678), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n677), .B1(new_n680), .B2(new_n688), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n689), .A2(new_n454), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n673), .B1(new_n690), .B2(new_n527), .ZN(G1328gat));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n693));
  INV_X1    g492(.A(new_n656), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n523), .ZN(new_n695));
  OR3_X1    g494(.A1(new_n670), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n693), .B1(new_n670), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n692), .B1(new_n698), .B2(KEYINPUT46), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n696), .A2(KEYINPUT105), .A3(new_n700), .A4(new_n697), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n523), .B1(new_n689), .B2(new_n694), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n703), .B1(KEYINPUT46), .B2(new_n698), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(G1329gat));
  INV_X1    g504(.A(KEYINPUT47), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n680), .A2(new_n688), .ZN(new_n707));
  INV_X1    g506(.A(new_n677), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(new_n462), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G43gat), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n670), .A2(G43gat), .A3(new_n663), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n706), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  AOI211_X1 g512(.A(KEYINPUT47), .B(new_n711), .C1(new_n709), .C2(G43gat), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(G1330gat));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT48), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n707), .A2(new_n439), .A3(new_n708), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(G50gat), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n440), .A2(G50gat), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n670), .B2(KEYINPUT106), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n670), .A2(KEYINPUT106), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n724), .A2(new_n725), .B1(new_n716), .B2(new_n717), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n719), .B1(new_n721), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(G50gat), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(new_n689), .B2(new_n439), .ZN(new_n729));
  INV_X1    g528(.A(new_n725), .ZN(new_n730));
  OAI22_X1  g529(.A1(new_n730), .A2(new_n723), .B1(KEYINPUT107), .B2(KEYINPUT48), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n729), .A2(new_n731), .A3(new_n718), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n727), .A2(new_n732), .ZN(G1331gat));
  NOR3_X1   g532(.A1(new_n675), .A2(new_n633), .A3(new_n566), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT108), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n686), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n454), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n580), .A2(G57gat), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n584), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n738), .B(new_n740), .ZN(G1332gat));
  AOI21_X1  g540(.A(new_n656), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n736), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT109), .ZN(new_n745));
  OR2_X1    g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1333gat));
  OAI21_X1  g546(.A(G71gat), .B1(new_n736), .B2(new_n463), .ZN(new_n748));
  INV_X1    g547(.A(G71gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n411), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n748), .B1(new_n736), .B2(new_n750), .ZN(new_n751));
  XOR2_X1   g550(.A(new_n751), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n440), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT110), .B(G78gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1335gat));
  NOR2_X1   g554(.A1(new_n566), .A2(new_n603), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n651), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n757), .B1(new_n680), .B2(new_n688), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759), .B2(new_n367), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n686), .A2(new_n678), .A3(new_n756), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n520), .A2(KEYINPUT102), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n682), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n632), .B1(new_n765), .B2(new_n512), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n766), .A2(KEYINPUT51), .A3(new_n756), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n651), .A2(new_n604), .A3(new_n454), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n760), .B1(new_n769), .B2(new_n770), .ZN(G1336gat));
  NOR3_X1   g570(.A1(new_n675), .A2(new_n656), .A3(G92gat), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT51), .B1(new_n766), .B2(new_n756), .ZN(new_n773));
  AND4_X1   g572(.A1(KEYINPUT51), .A2(new_n686), .A3(new_n678), .A4(new_n756), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n605), .B1(new_n758), .B2(new_n694), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT52), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n758), .A2(new_n694), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G92gat), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT111), .B1(new_n768), .B2(new_n772), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n779), .A2(new_n784), .ZN(G1337gat));
  OAI21_X1  g584(.A(G99gat), .B1(new_n759), .B2(new_n463), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n647), .B(new_n650), .Z(new_n787));
  NOR3_X1   g586(.A1(new_n787), .A2(G99gat), .A3(new_n663), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT112), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n786), .B1(new_n769), .B2(new_n789), .ZN(G1338gat));
  INV_X1    g589(.A(G106gat), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n791), .B1(new_n758), .B2(new_n439), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n675), .A2(G106gat), .A3(new_n440), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(new_n763), .B2(new_n767), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n793), .A2(new_n794), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT53), .B1(new_n792), .B2(new_n797), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(G1339gat));
  NAND4_X1  g600(.A1(new_n603), .A2(new_n565), .A3(new_n632), .A4(new_n787), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n636), .A2(new_n638), .A3(new_n642), .A4(new_n639), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n644), .A2(KEYINPUT54), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n640), .A2(new_n806), .A3(new_n643), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n650), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n803), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n647), .A2(new_n650), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n644), .A2(KEYINPUT54), .A3(new_n804), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n650), .A4(new_n807), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n809), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n552), .A2(new_n553), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n545), .B1(new_n544), .B2(new_n548), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n560), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n562), .B(new_n816), .C1(new_n630), .C2(new_n631), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n562), .A2(new_n816), .ZN(new_n819));
  OAI22_X1  g618(.A1(new_n565), .A2(new_n813), .B1(new_n787), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n818), .B1(new_n820), .B2(new_n632), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT99), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n603), .B(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n802), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(new_n367), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n826), .A2(new_n453), .ZN(new_n827));
  AOI21_X1  g626(.A(G113gat), .B1(new_n827), .B2(new_n566), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n656), .A2(new_n454), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n825), .A2(new_n441), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n565), .A2(new_n324), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(G1340gat));
  INV_X1    g631(.A(new_n830), .ZN(new_n833));
  OAI21_X1  g632(.A(G120gat), .B1(new_n833), .B2(new_n675), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n651), .A2(new_n326), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT113), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n827), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n834), .A2(new_n837), .ZN(G1341gat));
  NAND3_X1  g637(.A1(new_n827), .A2(new_n329), .A3(new_n603), .ZN(new_n839));
  OAI21_X1  g638(.A(G127gat), .B1(new_n833), .B2(new_n674), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(G1342gat));
  INV_X1    g640(.A(G134gat), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n842), .A3(new_n678), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n844));
  OAI21_X1  g643(.A(G134gat), .B1(new_n833), .B2(new_n632), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(G1343gat));
  INV_X1    g646(.A(G141gat), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n656), .A2(new_n454), .A3(new_n463), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n824), .A2(new_n439), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n850), .B1(new_n851), .B2(KEYINPUT57), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT114), .B1(new_n787), .B2(new_n819), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n651), .A2(new_n854), .A3(new_n562), .A4(new_n816), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n812), .A2(new_n810), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n811), .A2(new_n650), .A3(new_n807), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n859), .A2(KEYINPUT115), .A3(new_n803), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT115), .B1(new_n859), .B2(new_n803), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n857), .B(new_n858), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n566), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n809), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n859), .A2(KEYINPUT115), .A3(new_n803), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n857), .B1(new_n867), .B2(new_n858), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n856), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n632), .ZN(new_n870));
  INV_X1    g669(.A(new_n818), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n603), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n802), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n439), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n852), .B1(new_n874), .B2(KEYINPUT57), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n848), .B1(new_n875), .B2(new_n566), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n694), .A2(new_n440), .A3(new_n462), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n565), .A2(G141gat), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n826), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT117), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT58), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n882));
  INV_X1    g681(.A(new_n852), .ZN(new_n883));
  INV_X1    g682(.A(new_n603), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT116), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n566), .A3(new_n862), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n678), .B1(new_n887), .B2(new_n856), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n884), .B1(new_n888), .B2(new_n818), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n440), .B1(new_n889), .B2(new_n802), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n883), .B(new_n566), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(G141gat), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT58), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n882), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  AOI211_X1 g696(.A(KEYINPUT118), .B(new_n895), .C1(new_n892), .C2(G141gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n881), .B1(new_n897), .B2(new_n898), .ZN(G1344gat));
  AND2_X1   g698(.A1(new_n826), .A2(new_n877), .ZN(new_n900));
  INV_X1    g699(.A(G148gat), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(new_n901), .A3(new_n651), .ZN(new_n902));
  AOI211_X1 g701(.A(KEYINPUT59), .B(new_n901), .C1(new_n875), .C2(new_n651), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n891), .B(new_n439), .C1(new_n872), .C2(new_n873), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n851), .A2(KEYINPUT57), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n905), .A2(new_n651), .A3(new_n850), .A4(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n904), .B1(new_n907), .B2(G148gat), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n902), .B1(new_n903), .B2(new_n908), .ZN(G1345gat));
  AOI21_X1  g708(.A(G155gat), .B1(new_n900), .B2(new_n603), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n823), .A2(G155gat), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT119), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n910), .B1(new_n875), .B2(new_n912), .ZN(G1346gat));
  AOI21_X1  g712(.A(G162gat), .B1(new_n900), .B2(new_n678), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n632), .A2(new_n335), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n914), .B1(new_n875), .B2(new_n915), .ZN(G1347gat));
  NAND3_X1  g715(.A1(new_n694), .A2(new_n367), .A3(new_n513), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n825), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n566), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(G169gat), .ZN(G1348gat));
  NAND3_X1  g719(.A1(new_n918), .A2(new_n224), .A3(new_n651), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n825), .A2(new_n675), .A3(new_n917), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n224), .ZN(G1349gat));
  AOI21_X1  g722(.A(new_n208), .B1(new_n918), .B2(new_n823), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n603), .A2(new_n209), .A3(new_n211), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n918), .B2(new_n925), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT60), .Z(G1350gat));
  NAND2_X1  g726(.A1(new_n918), .A2(new_n678), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n928), .B(G190gat), .C1(KEYINPUT120), .C2(new_n929), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n929), .A2(KEYINPUT120), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  INV_X1    g732(.A(new_n215), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n932), .B(new_n933), .C1(new_n934), .C2(new_n928), .ZN(G1351gat));
  NOR3_X1   g734(.A1(new_n656), .A2(new_n454), .A3(new_n462), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n905), .A2(new_n566), .A3(new_n906), .A4(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(G197gat), .ZN(new_n938));
  INV_X1    g737(.A(new_n936), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT121), .B1(new_n851), .B2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT121), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n824), .A2(new_n941), .A3(new_n439), .A4(new_n936), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n565), .A2(G197gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n940), .A2(KEYINPUT122), .A3(new_n942), .A4(new_n943), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n938), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT123), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n938), .A2(new_n948), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1352gat));
  INV_X1    g752(.A(G204gat), .ZN(new_n954));
  INV_X1    g753(.A(new_n675), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n905), .A2(new_n955), .A3(new_n906), .A4(new_n936), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT124), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n958), .B1(new_n957), .B2(new_n956), .ZN(new_n959));
  NOR4_X1   g758(.A1(new_n851), .A2(G204gat), .A3(new_n787), .A4(new_n939), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT62), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(G1353gat));
  NAND4_X1  g761(.A1(new_n905), .A2(new_n603), .A3(new_n906), .A4(new_n936), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(G211gat), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n964), .A2(KEYINPUT63), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(KEYINPUT63), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n940), .A2(new_n277), .A3(new_n603), .A4(new_n942), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n967), .B(KEYINPUT125), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n965), .A2(new_n966), .A3(new_n968), .ZN(G1354gat));
  NAND3_X1  g768(.A1(new_n905), .A2(new_n906), .A3(new_n936), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n970), .A2(new_n278), .A3(new_n632), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n940), .A2(new_n678), .A3(new_n942), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(new_n278), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT126), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT126), .B1(new_n972), .B2(new_n278), .ZN(new_n976));
  NOR3_X1   g775(.A1(new_n971), .A2(new_n975), .A3(new_n976), .ZN(G1355gat));
endmodule


