//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  OR3_X1    g0023(.A1(new_n209), .A2(KEYINPUT64), .A3(G13), .ZN(new_n224));
  OAI21_X1  g0024(.A(KEYINPUT64), .B1(new_n209), .B2(G13), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT0), .Z(new_n228));
  INV_X1    g0028(.A(KEYINPUT65), .ZN(new_n229));
  INV_X1    g0029(.A(G13), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n229), .B1(new_n206), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g0031(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n234), .A2(new_n207), .ZN(new_n235));
  OAI21_X1  g0035(.A(G50), .B1(G58), .B2(G68), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT66), .Z(new_n237));
  AOI211_X1 g0037(.A(new_n223), .B(new_n228), .C1(new_n235), .C2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT67), .ZN(new_n248));
  XOR2_X1   g0048(.A(G50), .B(G58), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  AOI21_X1  g0055(.A(G20), .B1(new_n255), .B2(G97), .ZN(new_n256));
  INV_X1    g0056(.A(G283), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n256), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n231), .A2(new_n232), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G116), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G20), .ZN(new_n263));
  AND3_X1   g0063(.A1(new_n261), .A2(KEYINPUT83), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(KEYINPUT83), .B1(new_n261), .B2(new_n263), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n258), .B(new_n259), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G116), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n231), .A2(new_n232), .A3(new_n260), .A4(new_n267), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n269), .B1(new_n206), .B2(G33), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n268), .B1(new_n270), .B2(G116), .ZN(new_n271));
  INV_X1    g0071(.A(new_n258), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n261), .A2(new_n263), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT83), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n261), .A2(KEYINPUT83), .A3(new_n263), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n272), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT84), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT20), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n266), .B(new_n271), .C1(new_n277), .C2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT85), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n258), .B1(new_n264), .B2(new_n265), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(new_n278), .A3(KEYINPUT20), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT85), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n283), .A2(new_n284), .A3(new_n266), .A4(new_n271), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n233), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT68), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT68), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G1698), .ZN(new_n292));
  AND2_X1   g0092(.A1(KEYINPUT3), .A2(G33), .ZN(new_n293));
  NOR2_X1   g0093(.A1(KEYINPUT3), .A2(G33), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n290), .B(new_n292), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT82), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(new_n297), .A3(G257), .ZN(new_n298));
  INV_X1    g0098(.A(G257), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT82), .B1(new_n295), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT3), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n255), .ZN(new_n303));
  NAND2_X1  g0103(.A1(KEYINPUT3), .A2(G33), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G1698), .ZN(new_n306));
  INV_X1    g0106(.A(G303), .ZN(new_n307));
  OAI22_X1  g0107(.A1(new_n306), .A2(new_n220), .B1(new_n307), .B2(new_n305), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n288), .B1(new_n301), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT5), .B(G41), .ZN(new_n311));
  INV_X1    g0111(.A(G45), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n312), .A2(G1), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n287), .A2(G1), .A3(G13), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G274), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n314), .A2(new_n315), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(G270), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  OAI211_X1 g0120(.A(KEYINPUT21), .B(G169), .C1(new_n310), .C2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n308), .B1(new_n298), .B2(new_n300), .ZN(new_n322));
  OAI211_X1 g0122(.A(G179), .B(new_n319), .C1(new_n322), .C2(new_n288), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n286), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n319), .B1(new_n322), .B2(new_n288), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G169), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(new_n281), .B2(new_n285), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n325), .B1(KEYINPUT21), .B2(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(KEYINPUT78), .A2(G190), .ZN(new_n330));
  NOR2_X1   g0130(.A1(KEYINPUT78), .A2(G190), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n326), .A2(G200), .ZN(new_n334));
  AND4_X1   g0134(.A1(new_n285), .A2(new_n333), .A3(new_n281), .A4(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n337));
  INV_X1    g0137(.A(G150), .ZN(new_n338));
  NOR2_X1   g0138(.A1(G20), .A2(G33), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n207), .A2(G33), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT8), .B(G58), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n337), .B1(new_n338), .B2(new_n340), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n267), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n343), .A2(new_n261), .B1(new_n201), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n269), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n206), .A2(G20), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(G50), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n349), .B(KEYINPUT9), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n233), .A2(new_n287), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n290), .A2(new_n292), .A3(G222), .ZN(new_n352));
  INV_X1    g0152(.A(G223), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n352), .B(new_n305), .C1(new_n353), .C2(new_n289), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n351), .B(new_n354), .C1(G77), .C2(new_n305), .ZN(new_n355));
  INV_X1    g0155(.A(G41), .ZN(new_n356));
  AOI21_X1  g0156(.A(G1), .B1(new_n356), .B2(new_n312), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n357), .A2(new_n315), .A3(G274), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n315), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n359), .B1(G226), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n355), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G190), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(G200), .B2(new_n364), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n350), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT71), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT10), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n370), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n368), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n350), .A2(new_n367), .A3(KEYINPUT71), .A4(KEYINPUT10), .ZN(new_n375));
  INV_X1    g0175(.A(G169), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n364), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G179), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n355), .A2(new_n378), .A3(new_n363), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(new_n349), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n374), .A2(new_n375), .A3(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n293), .A2(new_n294), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT69), .B(G107), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n296), .A2(G232), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(new_n212), .B2(new_n306), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n351), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n359), .B1(G244), .B2(new_n362), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n389), .A2(new_n365), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(G200), .B2(new_n389), .ZN(new_n391));
  XOR2_X1   g0191(.A(KEYINPUT15), .B(G87), .Z(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n393), .A2(new_n341), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n342), .A2(new_n340), .B1(new_n207), .B2(new_n217), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n261), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n346), .A2(G77), .A3(new_n347), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n396), .B(new_n397), .C1(G77), .C2(new_n267), .ZN(new_n398));
  OR2_X1    g0198(.A1(new_n398), .A2(KEYINPUT70), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(KEYINPUT70), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n391), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n389), .A2(G179), .ZN(new_n404));
  AOI21_X1  g0204(.A(G169), .B1(new_n387), .B2(new_n388), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n401), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  XOR2_X1   g0208(.A(KEYINPUT8), .B(G58), .Z(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n347), .ZN(new_n410));
  OAI22_X1  g0210(.A1(new_n410), .A2(new_n269), .B1(new_n267), .B2(new_n409), .ZN(new_n411));
  INV_X1    g0211(.A(new_n261), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT7), .B1(new_n382), .B2(new_n207), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n303), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n304), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(G68), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n202), .A2(new_n211), .ZN(new_n417));
  NOR2_X1   g0217(.A1(G58), .A2(G68), .ZN(new_n418));
  OAI21_X1  g0218(.A(G20), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n339), .A2(G159), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(KEYINPUT16), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n412), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT16), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n303), .A2(new_n207), .A3(new_n304), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT7), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n211), .B1(new_n427), .B2(new_n414), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n419), .A2(new_n420), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n424), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n411), .B1(new_n423), .B2(new_n430), .ZN(new_n431));
  OAI211_X1 g0231(.A(G226), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n432));
  NAND2_X1  g0232(.A1(G33), .A2(G87), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n432), .B(new_n433), .C1(new_n295), .C2(new_n353), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n351), .ZN(new_n435));
  INV_X1    g0235(.A(G232), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n358), .B1(new_n436), .B2(new_n361), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n435), .A2(new_n438), .A3(new_n378), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n437), .B1(new_n351), .B2(new_n434), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n439), .B1(G169), .B2(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n431), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT18), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n411), .ZN(new_n445));
  INV_X1    g0245(.A(new_n429), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT16), .B1(new_n416), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n261), .B1(new_n428), .B2(new_n421), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n445), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n332), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n435), .A2(new_n438), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G200), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n451), .B1(new_n452), .B2(new_n440), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT17), .ZN(new_n455));
  INV_X1    g0255(.A(new_n440), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n376), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n449), .A2(new_n457), .A3(new_n439), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT18), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n456), .A2(G200), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n431), .A2(new_n460), .A3(new_n451), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT17), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n444), .A2(new_n455), .A3(new_n459), .A4(new_n463), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n381), .A2(new_n408), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G226), .ZN(new_n466));
  INV_X1    g0266(.A(G97), .ZN(new_n467));
  OAI22_X1  g0267(.A1(new_n295), .A2(new_n466), .B1(new_n255), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(G232), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT72), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n305), .A2(KEYINPUT72), .A3(G232), .A4(G1698), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n288), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n359), .B1(G238), .B2(new_n362), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT13), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT73), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT13), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n468), .B1(new_n472), .B2(new_n473), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n480), .B(new_n476), .C1(new_n481), .C2(new_n288), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n478), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n475), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n484), .A2(KEYINPUT73), .A3(new_n480), .A4(new_n476), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(G200), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n478), .A2(G190), .A3(new_n482), .ZN(new_n487));
  OR3_X1    g0287(.A1(new_n267), .A2(KEYINPUT12), .A3(G68), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT12), .B1(new_n267), .B2(G68), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n347), .A2(G68), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n490), .B1(new_n269), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT75), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n207), .A2(G33), .A3(G77), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n211), .A2(G20), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT74), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(KEYINPUT74), .A3(new_n495), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n339), .A2(G50), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n493), .B1(new_n501), .B2(new_n261), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n493), .A3(new_n261), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n492), .B1(new_n505), .B2(KEYINPUT11), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT11), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n503), .A2(new_n507), .A3(new_n504), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT76), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n504), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT11), .B1(new_n510), .B2(new_n502), .ZN(new_n511));
  INV_X1    g0311(.A(new_n492), .ZN(new_n512));
  AND4_X1   g0312(.A1(KEYINPUT76), .A2(new_n511), .A3(new_n508), .A4(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n486), .B(new_n487), .C1(new_n509), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT77), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n506), .A2(KEYINPUT76), .A3(new_n508), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n511), .A2(new_n508), .A3(new_n512), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT76), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT77), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n520), .A2(new_n521), .A3(new_n486), .A4(new_n487), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n515), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n465), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n483), .A2(G169), .A3(new_n485), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT14), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n483), .A2(KEYINPUT14), .A3(G169), .A4(new_n485), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n478), .A2(G179), .A3(new_n482), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n520), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n524), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(G257), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n535));
  INV_X1    g0335(.A(G294), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n535), .B1(new_n255), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n295), .A2(new_n214), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n351), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n318), .A2(G264), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n315), .A2(G274), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(new_n313), .A3(new_n311), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT88), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n539), .A2(new_n540), .A3(KEYINPUT88), .A4(new_n542), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(G169), .A3(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n539), .A2(new_n540), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n548), .A2(G179), .A3(new_n542), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n270), .A2(G107), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n344), .A2(new_n219), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT25), .ZN(new_n553));
  XNOR2_X1  g0353(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT23), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n556), .A2(new_n219), .A3(G20), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n262), .B2(new_n341), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n383), .A2(G20), .ZN(new_n559));
  XNOR2_X1  g0359(.A(KEYINPUT87), .B(KEYINPUT23), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n305), .A2(new_n207), .A3(G87), .ZN(new_n562));
  XNOR2_X1  g0362(.A(KEYINPUT86), .B(KEYINPUT22), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n305), .A2(new_n563), .A3(new_n207), .A4(G87), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n561), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT24), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT24), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n561), .A2(new_n565), .A3(new_n569), .A4(new_n566), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n555), .B1(new_n571), .B2(new_n261), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n550), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n314), .A2(new_n315), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n542), .B1(new_n299), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n382), .A2(new_n289), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT4), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT79), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n296), .A2(G244), .A3(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(KEYINPUT79), .B(new_n579), .C1(new_n295), .C2(new_n218), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n578), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n576), .B1(new_n583), .B2(new_n351), .ZN(new_n584));
  OR3_X1    g0384(.A1(new_n584), .A2(KEYINPUT80), .A3(new_n452), .ZN(new_n585));
  OAI21_X1  g0385(.A(KEYINPUT80), .B1(new_n584), .B2(new_n452), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n270), .A2(G97), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(G97), .B2(new_n267), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n219), .A2(KEYINPUT6), .A3(G97), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n467), .A2(new_n219), .ZN(new_n590));
  NOR2_X1   g0390(.A1(G97), .A2(G107), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n589), .B1(new_n592), .B2(KEYINPUT6), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n593), .A2(G20), .B1(G77), .B2(new_n339), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n384), .B1(new_n413), .B2(new_n415), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n412), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n588), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n584), .A2(G190), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n585), .A2(new_n586), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n383), .A2(new_n213), .A3(new_n467), .ZN(new_n600));
  NAND3_X1  g0400(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n207), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n305), .A2(new_n207), .A3(G68), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT19), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n341), .B2(new_n467), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n607), .A2(new_n261), .B1(new_n344), .B2(new_n393), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n270), .A2(G87), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n541), .A2(new_n313), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n315), .B(G250), .C1(G1), .C2(new_n312), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(G244), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n614));
  OAI221_X1 g0414(.A(new_n614), .B1(new_n255), .B2(new_n262), .C1(new_n295), .C2(new_n212), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n613), .B1(new_n615), .B2(new_n351), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n616), .A2(new_n452), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n610), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n615), .A2(new_n351), .ZN(new_n619));
  INV_X1    g0419(.A(new_n613), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(KEYINPUT81), .B1(new_n621), .B2(new_n365), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT81), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n616), .A2(new_n623), .A3(G190), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n270), .A2(new_n392), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n608), .A2(new_n626), .B1(new_n621), .B2(new_n376), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n616), .A2(new_n378), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n618), .A2(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(G190), .B1(new_n545), .B2(new_n546), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n543), .A2(new_n452), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n572), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n584), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n376), .ZN(new_n634));
  INV_X1    g0434(.A(new_n597), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n584), .A2(new_n378), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n599), .A2(new_n629), .A3(new_n632), .A4(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  AND4_X1   g0439(.A1(new_n336), .A2(new_n534), .A3(new_n574), .A4(new_n639), .ZN(G372));
  INV_X1    g0440(.A(new_n380), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n455), .A2(new_n463), .ZN(new_n642));
  INV_X1    g0442(.A(new_n407), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n514), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n642), .B1(new_n533), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n444), .A2(new_n459), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n374), .A2(new_n375), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n641), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n534), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n574), .B(new_n325), .C1(KEYINPUT21), .C2(new_n328), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT89), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n327), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n286), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT21), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n657), .A2(KEYINPUT89), .A3(new_n325), .A4(new_n574), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n653), .A2(new_n639), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n618), .A2(new_n625), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n627), .A2(new_n628), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n660), .B1(new_n663), .B2(new_n637), .ZN(new_n664));
  INV_X1    g0464(.A(new_n637), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(KEYINPUT26), .A3(new_n629), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n664), .A2(new_n666), .B1(new_n628), .B2(new_n627), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n659), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n649), .B1(new_n650), .B2(new_n668), .ZN(G369));
  NAND3_X1  g0469(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n286), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n336), .A2(new_n676), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n655), .A2(new_n656), .B1(new_n286), .B2(new_n324), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n677), .B(KEYINPUT90), .C1(new_n678), .C2(new_n676), .ZN(new_n679));
  OR3_X1    g0479(.A1(new_n678), .A2(KEYINPUT90), .A3(new_n676), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G330), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n550), .A2(new_n573), .A3(new_n675), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n573), .B1(new_n550), .B2(new_n675), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT91), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(new_n685), .A3(new_n632), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n685), .B1(new_n684), .B2(new_n632), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n683), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n682), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n574), .A2(new_n675), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT92), .B1(new_n678), .B2(new_n675), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT92), .ZN(new_n693));
  INV_X1    g0493(.A(new_n675), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n329), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n691), .B1(new_n696), .B2(new_n689), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n690), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT93), .Z(G399));
  INV_X1    g0499(.A(new_n226), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  OR4_X1    g0501(.A1(new_n206), .A2(new_n701), .A3(G116), .A4(new_n600), .ZN(new_n702));
  INV_X1    g0502(.A(new_n237), .ZN(new_n703));
  INV_X1    g0503(.A(new_n701), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  XOR2_X1   g0505(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n706));
  XNOR2_X1  g0506(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n336), .A2(new_n639), .A3(new_n574), .A4(new_n694), .ZN(new_n708));
  INV_X1    g0508(.A(new_n323), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n548), .A2(new_n616), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n709), .A2(new_n710), .A3(KEYINPUT30), .A4(new_n584), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n584), .A2(new_n548), .A3(new_n616), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n323), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n616), .A2(G179), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n633), .A2(new_n326), .A3(new_n715), .A4(new_n543), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n711), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n717), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n718));
  AOI21_X1  g0518(.A(KEYINPUT31), .B1(new_n717), .B2(new_n675), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n708), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(G330), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n675), .B1(new_n659), .B2(new_n667), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n725), .A2(KEYINPUT29), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n639), .A2(new_n651), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n675), .B1(new_n667), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT29), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n724), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n707), .B1(new_n730), .B2(G1), .ZN(G364));
  NOR2_X1   g0531(.A1(new_n230), .A2(G20), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n206), .B1(new_n732), .B2(G45), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n701), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n682), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n679), .A2(new_n680), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G330), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G13), .A2(G33), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n234), .B1(G20), .B2(new_n376), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n743), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n700), .A2(new_n305), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(G45), .B2(new_n703), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n749), .B1(new_n250), .B2(G45), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n226), .A2(G355), .A3(new_n305), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(G116), .B2(new_n226), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n747), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n735), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n207), .A2(G179), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(G190), .A3(G200), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n307), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n755), .A2(new_n365), .A3(new_n452), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n305), .B(new_n757), .C1(G329), .C2(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n207), .A2(new_n378), .A3(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n365), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n755), .A2(new_n365), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n763), .A2(G311), .B1(new_n765), .B2(G283), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n450), .A2(new_n761), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n378), .A2(new_n452), .A3(G190), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n768), .A2(G322), .B1(G294), .B2(new_n770), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n207), .A2(new_n378), .A3(new_n452), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n332), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(G190), .ZN(new_n775));
  XNOR2_X1  g0575(.A(KEYINPUT33), .B(G317), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G326), .A2(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n760), .A2(new_n766), .A3(new_n771), .A4(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G159), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n758), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT32), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n768), .A2(G58), .B1(new_n775), .B2(G68), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n764), .A2(new_n219), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(new_n774), .B2(G50), .ZN(new_n784));
  INV_X1    g0584(.A(new_n756), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n382), .B1(new_n785), .B2(G87), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n781), .A2(new_n782), .A3(new_n784), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n770), .B(KEYINPUT96), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G97), .ZN(new_n789));
  AND2_X1   g0589(.A1(new_n762), .A2(KEYINPUT95), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n762), .A2(KEYINPUT95), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n789), .B1(new_n792), .B2(new_n217), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n778), .B1(new_n787), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n754), .B1(new_n794), .B2(new_n746), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n753), .A2(new_n795), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n737), .A2(new_n740), .B1(new_n745), .B2(new_n796), .ZN(G396));
  NAND3_X1  g0597(.A1(new_n406), .A2(new_n401), .A3(new_n694), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n694), .B1(new_n399), .B2(new_n400), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(new_n391), .B2(new_n402), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n798), .B1(new_n800), .B2(new_n643), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n725), .B(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n724), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n735), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(new_n804), .B2(new_n803), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n746), .A2(new_n741), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n754), .B1(new_n807), .B2(new_n217), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n765), .A2(G68), .ZN(new_n809));
  INV_X1    g0609(.A(G132), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n809), .B(new_n305), .C1(new_n810), .C2(new_n758), .ZN(new_n811));
  INV_X1    g0611(.A(new_n770), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n812), .A2(new_n202), .B1(new_n756), .B2(new_n201), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G137), .A2(new_n774), .B1(new_n775), .B2(G150), .ZN(new_n814));
  INV_X1    g0614(.A(G143), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n814), .B1(new_n815), .B2(new_n767), .C1(new_n792), .C2(new_n779), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT97), .Z(new_n817));
  INV_X1    g0617(.A(KEYINPUT34), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n811), .B(new_n813), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n818), .B2(new_n817), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n764), .A2(new_n213), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n767), .A2(new_n536), .B1(new_n219), .B2(new_n756), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n821), .B(new_n822), .C1(G283), .C2(new_n775), .ZN(new_n823));
  INV_X1    g0623(.A(G311), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n382), .B1(new_n758), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(new_n774), .B2(G303), .ZN(new_n826));
  INV_X1    g0626(.A(new_n792), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(G116), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n823), .A2(new_n826), .A3(new_n789), .A4(new_n828), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n820), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n746), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n808), .B1(new_n802), .B2(new_n742), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n806), .A2(new_n832), .ZN(G384));
  NOR2_X1   g0633(.A1(new_n732), .A2(new_n206), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT101), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT37), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n442), .A2(new_n454), .ZN(new_n837));
  OAI21_X1  g0637(.A(KEYINPUT100), .B1(new_n431), .B2(new_n673), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT100), .ZN(new_n839));
  INV_X1    g0639(.A(new_n673), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n449), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n836), .B1(new_n837), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n449), .A2(new_n840), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n458), .A2(new_n461), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n845), .A2(KEYINPUT37), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n835), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  NOR3_X1   g0647(.A1(new_n431), .A2(KEYINPUT100), .A3(new_n673), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n839), .B1(new_n449), .B2(new_n840), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n458), .A2(new_n461), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT37), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n837), .A2(new_n836), .A3(new_n844), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n852), .A2(KEYINPUT101), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n464), .A2(new_n850), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n847), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT38), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n847), .A2(new_n854), .A3(KEYINPUT38), .A4(new_n855), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(KEYINPUT102), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n532), .A2(new_n675), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT99), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT99), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n516), .A2(new_n519), .A3(new_n863), .A4(new_n675), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n514), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n533), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n531), .B1(new_n515), .B2(new_n522), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n866), .B1(new_n861), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT102), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n856), .A2(new_n869), .A3(new_n857), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n801), .B1(new_n708), .B2(new_n720), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n860), .A2(new_n868), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT40), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT106), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT106), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n872), .A2(new_n876), .A3(new_n873), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n868), .A2(new_n871), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n464), .A2(new_n449), .A3(new_n840), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n845), .A2(KEYINPUT37), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n853), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n857), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n859), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n885), .A2(new_n873), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n879), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n878), .A2(new_n887), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n888), .B(KEYINPUT107), .Z(new_n889));
  NOR2_X1   g0689(.A1(new_n650), .A2(new_n722), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n723), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n889), .B2(new_n890), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n534), .A2(new_n726), .A3(new_n729), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n649), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT105), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n675), .B(new_n801), .C1(new_n659), .C2(new_n667), .ZN(new_n896));
  INV_X1    g0696(.A(new_n798), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n868), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n860), .A2(new_n870), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n899), .A2(new_n900), .B1(new_n646), .B2(new_n673), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n860), .A2(KEYINPUT39), .A3(new_n870), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT104), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT39), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n903), .B1(new_n885), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n533), .A2(new_n675), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT103), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n907), .B(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n860), .A2(new_n903), .A3(KEYINPUT39), .A4(new_n870), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n906), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n901), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n895), .B(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n834), .B1(new_n892), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n914), .B2(new_n892), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n593), .A2(KEYINPUT35), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n593), .A2(KEYINPUT35), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n917), .A2(G116), .A3(new_n235), .A4(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT36), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n703), .A2(new_n217), .A3(new_n417), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n201), .B2(G68), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n922), .A2(new_n206), .A3(G13), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT98), .Z(new_n924));
  NAND3_X1  g0724(.A1(new_n916), .A2(new_n920), .A3(new_n924), .ZN(G367));
  INV_X1    g0725(.A(new_n748), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n926), .A2(new_n245), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n747), .B1(new_n226), .B2(new_n393), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n735), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(G137), .ZN(new_n930));
  INV_X1    g0730(.A(new_n775), .ZN(new_n931));
  OAI221_X1 g0731(.A(new_n305), .B1(new_n930), .B2(new_n758), .C1(new_n931), .C2(new_n779), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n202), .A2(new_n756), .B1(new_n764), .B2(new_n217), .ZN(new_n933));
  INV_X1    g0733(.A(new_n774), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n934), .A2(new_n815), .B1(new_n338), .B2(new_n767), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n788), .A2(G68), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n936), .B(new_n937), .C1(new_n201), .C2(new_n792), .ZN(new_n938));
  INV_X1    g0738(.A(G317), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n382), .B1(new_n939), .B2(new_n758), .C1(new_n934), .C2(new_n824), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT46), .B1(new_n785), .B2(G116), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n785), .A2(KEYINPUT46), .A3(G116), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n931), .A2(new_n536), .B1(new_n307), .B2(new_n767), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(G97), .B2(new_n765), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n827), .A2(G283), .B1(new_n384), .B2(new_n770), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT115), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n943), .B(new_n945), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n946), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n949), .A2(KEYINPUT115), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n938), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT47), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n929), .B1(new_n952), .B2(new_n746), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n610), .A2(new_n675), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n662), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n629), .B2(new_n954), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n743), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n689), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n681), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n681), .A2(new_n959), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n695), .B(new_n692), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n690), .A2(new_n696), .A3(new_n960), .ZN(new_n964));
  AND3_X1   g0764(.A1(new_n963), .A2(new_n964), .A3(new_n730), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n599), .B(new_n637), .C1(new_n597), .C2(new_n694), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n665), .A2(new_n675), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(KEYINPUT113), .B1(new_n697), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT113), .ZN(new_n970));
  INV_X1    g0770(.A(new_n968), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n684), .A2(new_n632), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(KEYINPUT91), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n686), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n974), .A2(new_n683), .B1(new_n692), .B2(new_n695), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n970), .B(new_n971), .C1(new_n975), .C2(new_n691), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n969), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT44), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n980));
  NOR4_X1   g0780(.A1(new_n975), .A2(new_n691), .A3(new_n971), .A4(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n980), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(new_n697), .B2(new_n968), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n969), .A2(KEYINPUT44), .A3(new_n976), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n979), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n986), .A2(KEYINPUT114), .A3(new_n962), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n965), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n962), .B1(new_n986), .B2(KEYINPUT114), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n730), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n701), .B(KEYINPUT41), .Z(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n734), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n962), .A2(new_n968), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT111), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n975), .A2(new_n968), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(KEYINPUT42), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n966), .A2(new_n574), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n675), .B1(new_n999), .B2(new_n637), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT109), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT42), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n975), .A2(new_n1005), .A3(new_n968), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT110), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n998), .A2(KEYINPUT109), .A3(new_n1001), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT43), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1009), .A2(KEYINPUT108), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(KEYINPUT108), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n956), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1004), .A2(new_n1007), .A3(new_n1008), .A4(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n995), .B2(new_n994), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1004), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1012), .B1(new_n1009), .B2(new_n956), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n996), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1019), .A2(new_n995), .A3(new_n994), .A4(new_n1013), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n958), .B1(new_n993), .B2(new_n1021), .ZN(G387));
  INV_X1    g0822(.A(new_n730), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n964), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n696), .B1(new_n690), .B2(new_n960), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n963), .A2(new_n964), .A3(new_n730), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1026), .A2(new_n701), .A3(new_n1027), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n242), .A2(new_n312), .A3(new_n305), .ZN(new_n1029));
  OR3_X1    g0829(.A1(new_n342), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1030));
  OAI21_X1  g0830(.A(KEYINPUT50), .B1(new_n342), .B2(G50), .ZN(new_n1031));
  AOI21_X1  g0831(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  AOI211_X1 g0833(.A(G116), .B(new_n600), .C1(new_n1033), .C2(new_n382), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1029), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1035), .A2(new_n700), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n747), .B1(new_n219), .B2(new_n226), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n774), .A2(G159), .B1(new_n763), .B2(G68), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n201), .B2(new_n767), .C1(new_n342), .C2(new_n931), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n382), .B1(new_n759), .B2(G150), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n217), .B2(new_n756), .C1(new_n467), .C2(new_n764), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT116), .Z(new_n1042));
  AOI211_X1 g0842(.A(new_n1039), .B(new_n1042), .C1(new_n392), .C2(new_n788), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n764), .A2(new_n262), .ZN(new_n1044));
  INV_X1    g0844(.A(G326), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n382), .B1(new_n758), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n774), .A2(G322), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n768), .A2(G317), .B1(new_n775), .B2(G311), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(new_n792), .C2(new_n307), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT48), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n785), .A2(G294), .B1(new_n770), .B2(G283), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1044), .B(new_n1046), .C1(new_n1055), .C2(KEYINPUT49), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1055), .A2(KEYINPUT49), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1043), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n735), .B1(new_n1036), .B2(new_n1037), .C1(new_n1058), .C2(new_n831), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n959), .B2(new_n743), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1060), .B1(new_n1061), .B2(new_n734), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1028), .A2(new_n1062), .ZN(G393));
  NAND2_X1  g0863(.A1(new_n986), .A2(new_n962), .ZN(new_n1064));
  AOI21_X1  g0864(.A(KEYINPUT44), .B1(new_n969), .B2(new_n976), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n981), .A2(new_n983), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1067), .A2(new_n690), .A3(new_n985), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1064), .A2(new_n1068), .A3(new_n734), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n926), .A2(new_n253), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n747), .B1(new_n467), .B2(new_n226), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n735), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n934), .A2(new_n939), .B1(new_n824), .B2(new_n767), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT52), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n305), .B(new_n783), .C1(G322), .C2(new_n759), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n812), .A2(new_n262), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n762), .A2(new_n536), .B1(new_n756), .B2(new_n257), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(G303), .C2(new_n775), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1074), .A2(new_n1075), .A3(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n934), .A2(new_n338), .B1(new_n779), .B2(new_n767), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT51), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n342), .B2(new_n792), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n382), .B(new_n821), .C1(G143), .C2(new_n759), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n788), .A2(G77), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n775), .A2(G50), .B1(G68), .B2(new_n785), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1079), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1072), .B1(new_n1087), .B2(new_n746), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n968), .B2(new_n744), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1069), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n986), .A2(new_n962), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n690), .B1(new_n1067), .B2(new_n985), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1027), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n701), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n988), .A2(new_n989), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1091), .B1(new_n1095), .B2(new_n1096), .ZN(G390));
  NAND2_X1  g0897(.A1(new_n906), .A2(new_n911), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n898), .A2(new_n909), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n868), .A2(new_n871), .A3(G330), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n885), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n909), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n800), .A2(new_n643), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n897), .B1(new_n728), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n531), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n861), .B1(new_n523), .B2(new_n1107), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n862), .A2(new_n865), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1108), .B1(new_n533), .B2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1106), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1103), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1100), .A2(new_n1101), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1101), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n906), .A2(new_n911), .B1(new_n909), .B2(new_n898), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n1112), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1114), .A2(new_n1117), .A3(new_n734), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1098), .A2(new_n741), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n807), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n735), .B1(new_n409), .B2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT119), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n827), .A2(G97), .B1(new_n384), .B2(new_n775), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1123), .A2(KEYINPUT120), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(KEYINPUT120), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n382), .B1(new_n758), .B2(new_n536), .C1(new_n213), .C2(new_n756), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n809), .B1(new_n767), .B2(new_n262), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1126), .B(new_n1127), .C1(G283), .C2(new_n774), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1124), .A2(new_n1084), .A3(new_n1125), .A4(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n931), .A2(new_n930), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n382), .B(new_n1130), .C1(G125), .C2(new_n759), .ZN(new_n1131));
  INV_X1    g0931(.A(G128), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n934), .A2(new_n1132), .B1(new_n201), .B2(new_n764), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G132), .B2(new_n768), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n788), .A2(G159), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT54), .B(G143), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT53), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n756), .B2(new_n338), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n785), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n827), .A2(new_n1137), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1131), .A2(new_n1134), .A3(new_n1135), .A4(new_n1141), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1129), .A2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1119), .B(new_n1122), .C1(new_n831), .C2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT117), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n721), .A2(new_n1146), .A3(G330), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n802), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1146), .B1(new_n721), .B2(G330), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1110), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n721), .A2(new_n802), .A3(G330), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1110), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n1101), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n896), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n798), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1150), .A2(new_n1151), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n893), .B(new_n649), .C1(new_n650), .C2(new_n804), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1145), .A2(new_n1160), .A3(KEYINPUT118), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT118), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1117), .B(new_n1114), .C1(new_n1159), .C2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n701), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1118), .B(new_n1144), .C1(new_n1162), .C2(new_n1165), .ZN(G378));
  AOI21_X1  g0966(.A(new_n723), .B1(new_n879), .B2(new_n886), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n872), .A2(new_n876), .A3(new_n873), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n876), .B1(new_n872), .B2(new_n873), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n349), .A2(new_n840), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n381), .B(new_n1171), .Z(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1172), .B(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1170), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1174), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1167), .B(new_n1176), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1175), .A2(new_n913), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n913), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n734), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1174), .A2(new_n741), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n735), .B1(G50), .B2(new_n1120), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT123), .Z(new_n1183));
  OAI22_X1  g0983(.A1(new_n762), .A2(new_n930), .B1(new_n756), .B2(new_n1136), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n768), .A2(G128), .B1(new_n774), .B2(G125), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n810), .B2(new_n931), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1184), .B(new_n1186), .C1(G150), .C2(new_n788), .ZN(new_n1187));
  XOR2_X1   g0987(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1188));
  OR2_X1    g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n765), .A2(G159), .ZN(new_n1191));
  AOI211_X1 g0991(.A(G33), .B(G41), .C1(new_n759), .C2(G124), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n774), .A2(G116), .B1(G58), .B2(new_n765), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1194), .B1(new_n467), .B2(new_n931), .C1(new_n393), .C2(new_n762), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n767), .A2(new_n219), .B1(new_n257), .B2(new_n758), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n382), .A2(new_n356), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n785), .B2(G77), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1198), .A2(KEYINPUT121), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(KEYINPUT121), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n937), .A2(new_n1200), .ZN(new_n1201));
  NOR4_X1   g1001(.A1(new_n1195), .A2(new_n1196), .A3(new_n1199), .A4(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(KEYINPUT58), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1197), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1202), .A2(KEYINPUT58), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1193), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1183), .B1(new_n1206), .B2(new_n746), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1181), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1180), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n913), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1176), .B1(new_n878), .B2(new_n1167), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1177), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1210), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1175), .A2(new_n913), .A3(new_n1177), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1158), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1157), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1114), .A2(new_n1117), .A3(new_n1216), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1213), .A2(new_n1214), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n704), .B1(new_n1218), .B2(KEYINPUT57), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1217), .A2(new_n1215), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT57), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1209), .B1(new_n1219), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(G375));
  NAND2_X1  g1026(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1160), .A2(new_n992), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n754), .B1(new_n807), .B2(new_n211), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n931), .A2(new_n1136), .B1(new_n779), .B2(new_n756), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n934), .A2(new_n810), .B1(new_n930), .B2(new_n767), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n762), .A2(new_n338), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n305), .B1(new_n758), .B2(new_n1132), .C1(new_n202), .C2(new_n764), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n788), .A2(G50), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n827), .A2(new_n384), .B1(new_n392), .B2(new_n788), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n934), .A2(new_n536), .B1(new_n467), .B2(new_n756), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n931), .A2(new_n262), .B1(new_n257), .B2(new_n767), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n382), .B1(new_n758), .B2(new_n307), .C1(new_n217), .C2(new_n764), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1234), .A2(new_n1235), .B1(new_n1236), .B2(new_n1240), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1229), .B1(new_n831), .B2(new_n1241), .C1(new_n868), .C2(new_n742), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1216), .B2(new_n734), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1228), .A2(new_n1244), .ZN(G381));
  INV_X1    g1045(.A(G396), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1028), .A2(new_n1062), .A3(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(G384), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1248), .A2(new_n1249), .A3(new_n1244), .A4(new_n1228), .ZN(new_n1250));
  NOR4_X1   g1050(.A1(G387), .A2(G378), .A3(new_n1250), .A4(G390), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1225), .ZN(G407));
  NAND2_X1  g1052(.A1(new_n1118), .A2(new_n1144), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1165), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1253), .B1(new_n1254), .B2(new_n1161), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n674), .A2(G213), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1225), .A2(new_n1255), .A3(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(G407), .A2(G213), .A3(new_n1258), .ZN(new_n1259));
  XOR2_X1   g1059(.A(new_n1259), .B(KEYINPUT124), .Z(G409));
  AOI22_X1  g1060(.A1(new_n1220), .A2(new_n734), .B1(new_n1181), .B2(new_n1207), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1221), .B(KEYINPUT57), .C1(new_n1178), .C2(new_n1179), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n701), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT57), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1264));
  OAI211_X1 g1064(.A(G378), .B(new_n1261), .C1(new_n1263), .C2(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1221), .B(new_n992), .C1(new_n1178), .C2(new_n1179), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1266), .A2(new_n1180), .A3(new_n1208), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1255), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1257), .B1(new_n1265), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT62), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT60), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1227), .B1(new_n1159), .B2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1157), .A2(KEYINPUT60), .A3(new_n1158), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(new_n701), .A3(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(G384), .A3(new_n1244), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(G384), .B1(new_n1274), .B2(new_n1244), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1269), .A2(new_n1270), .A3(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT61), .ZN(new_n1280));
  OAI211_X1 g1080(.A(G2897), .B(new_n1257), .C1(new_n1276), .C2(new_n1277), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1277), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1257), .A2(G2897), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1282), .A2(new_n1275), .A3(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1281), .A2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1280), .B1(new_n1269), .B2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1270), .B1(new_n1269), .B2(new_n1278), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1279), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n958), .B(G390), .C1(new_n993), .C2(new_n1021), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(KEYINPUT126), .ZN(new_n1290));
  INV_X1    g1090(.A(G390), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(G387), .A2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1246), .B1(new_n1028), .B2(new_n1062), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1247), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n986), .A2(KEYINPUT114), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n690), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1298), .A2(new_n965), .A3(new_n987), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n991), .B1(new_n1299), .B2(new_n730), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1296), .B1(new_n1300), .B2(new_n734), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT126), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1301), .A2(new_n1302), .A3(new_n958), .A4(G390), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1290), .A2(new_n1292), .A3(new_n1295), .A4(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1294), .A2(KEYINPUT125), .A3(new_n1247), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT125), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1306), .B1(new_n1248), .B2(new_n1293), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1289), .ZN(new_n1309));
  AOI21_X1  g1109(.A(G390), .B1(new_n1301), .B2(new_n958), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1308), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1304), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1265), .A2(new_n1268), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1256), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1285), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT61), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1313), .A2(new_n1256), .A3(new_n1278), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT63), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1316), .A2(new_n1312), .A3(new_n1319), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1313), .A2(KEYINPUT63), .A3(new_n1278), .A4(new_n1256), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(KEYINPUT127), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT127), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1269), .A2(new_n1323), .A3(KEYINPUT63), .A4(new_n1278), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  OAI22_X1  g1125(.A1(new_n1288), .A2(new_n1312), .B1(new_n1320), .B2(new_n1325), .ZN(G405));
  NOR2_X1   g1126(.A1(new_n1225), .A2(G378), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1265), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1312), .A2(new_n1329), .ZN(new_n1330));
  OAI211_X1 g1130(.A(new_n1304), .B(new_n1311), .C1(new_n1327), .C2(new_n1328), .ZN(new_n1331));
  AND3_X1   g1131(.A1(new_n1330), .A2(new_n1278), .A3(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1278), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1332), .A2(new_n1333), .ZN(G402));
endmodule


