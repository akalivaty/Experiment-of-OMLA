//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n548, new_n549, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n561, new_n565, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n593, new_n594, new_n597,
    new_n598, new_n600, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT67), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(G125), .ZN(new_n457));
  INV_X1    g032(.A(KEYINPUT68), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n458), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n459), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT68), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n457), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(G2105), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n464), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT69), .B(KEYINPUT3), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n473), .B1(new_n474), .B2(new_n461), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(KEYINPUT3), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n459), .A2(KEYINPUT69), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n472), .B(G2104), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G2105), .ZN(new_n480));
  NAND4_X1  g055(.A1(new_n475), .A2(G137), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n461), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G101), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT71), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n471), .A2(new_n485), .ZN(G160));
  AND2_X1   g061(.A1(new_n475), .A2(new_n479), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT72), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n489), .B(new_n490), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n487), .A2(new_n480), .ZN(new_n492));
  MUX2_X1   g067(.A(G100), .B(G112), .S(G2105), .Z(new_n493));
  AOI22_X1  g068(.A1(new_n492), .A2(G136), .B1(G2104), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  AND2_X1   g071(.A1(new_n480), .A2(G138), .ZN(new_n497));
  AND2_X1   g072(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n498));
  NOR2_X1   g073(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n500), .B1(new_n466), .B2(new_n463), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n475), .A2(G138), .A3(new_n479), .A4(new_n480), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n475), .A2(G126), .A3(new_n479), .A4(G2105), .ZN(new_n504));
  MUX2_X1   g079(.A(G102), .B(G114), .S(G2105), .Z(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G2104), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n503), .A2(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G50), .ZN(new_n511));
  XNOR2_X1  g086(.A(new_n511), .B(KEYINPUT74), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G88), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n512), .A2(new_n518), .ZN(G166));
  NAND2_X1  g094(.A1(new_n509), .A2(G543), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT75), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n521), .A2(G51), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT76), .B(G89), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n509), .A2(new_n525), .B1(G63), .B2(G651), .ZN(new_n526));
  XOR2_X1   g101(.A(KEYINPUT5), .B(G543), .Z(new_n527));
  OAI21_X1  g102(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n522), .A2(new_n528), .ZN(G168));
  NAND2_X1  g104(.A1(G77), .A2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G651), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  INV_X1    g109(.A(new_n514), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n536), .B1(new_n521), .B2(G52), .ZN(G171));
  NAND2_X1  g112(.A1(new_n521), .A2(G43), .ZN(new_n538));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G56), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n527), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n541), .A2(G651), .B1(new_n514), .B2(G81), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  AND3_X1   g120(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G36), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n546), .A2(new_n549), .ZN(G188));
  XNOR2_X1  g125(.A(new_n513), .B(KEYINPUT77), .ZN(new_n551));
  INV_X1    g126(.A(G65), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g128(.A1(G78), .A2(G543), .ZN(new_n554));
  OAI21_X1  g129(.A(G651), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OR3_X1    g131(.A1(new_n520), .A2(KEYINPUT9), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT9), .B1(new_n520), .B2(new_n556), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n557), .A2(new_n558), .B1(G91), .B2(new_n514), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n555), .A2(new_n559), .ZN(G299));
  NAND2_X1  g135(.A1(new_n521), .A2(G52), .ZN(new_n561));
  OAI211_X1 g136(.A(new_n561), .B(new_n533), .C1(new_n534), .C2(new_n535), .ZN(G301));
  INV_X1    g137(.A(G168), .ZN(G286));
  INV_X1    g138(.A(G166), .ZN(G303));
  NAND2_X1  g139(.A1(new_n514), .A2(G87), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n510), .A2(G49), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n567));
  AND3_X1   g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT78), .ZN(G288));
  NAND2_X1  g144(.A1(new_n514), .A2(G86), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n510), .A2(G48), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n573), .A2(new_n516), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G305));
  AOI22_X1  g151(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(new_n516), .ZN(new_n578));
  XOR2_X1   g153(.A(new_n578), .B(KEYINPUT79), .Z(new_n579));
  AOI22_X1  g154(.A1(new_n521), .A2(G47), .B1(G85), .B2(new_n514), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G290));
  NAND2_X1  g156(.A1(new_n514), .A2(G92), .ZN(new_n582));
  XOR2_X1   g157(.A(new_n582), .B(KEYINPUT10), .Z(new_n583));
  INV_X1    g158(.A(G66), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n551), .A2(new_n584), .ZN(new_n585));
  AND2_X1   g160(.A1(G79), .A2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n521), .A2(G54), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n583), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(G868), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g166(.A(new_n590), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g167(.A1(G286), .A2(G868), .ZN(new_n593));
  XOR2_X1   g168(.A(G299), .B(KEYINPUT80), .Z(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(G868), .ZN(G297));
  OAI21_X1  g170(.A(new_n593), .B1(new_n594), .B2(G868), .ZN(G280));
  AND3_X1   g171(.A1(new_n583), .A2(new_n587), .A3(new_n588), .ZN(new_n597));
  INV_X1    g172(.A(G559), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(G860), .ZN(G148));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n598), .ZN(new_n600));
  MUX2_X1   g175(.A(new_n543), .B(new_n600), .S(G868), .Z(G323));
  XNOR2_X1  g176(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g177(.A1(new_n463), .A2(new_n466), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(new_n482), .ZN(new_n604));
  XOR2_X1   g179(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n605));
  XOR2_X1   g180(.A(new_n604), .B(new_n605), .Z(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT13), .ZN(new_n607));
  INV_X1    g182(.A(G2100), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n492), .A2(G135), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n488), .A2(G123), .ZN(new_n611));
  OAI21_X1  g186(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT82), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n614), .B(new_n615), .C1(G111), .C2(new_n480), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n610), .A2(new_n611), .A3(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G2096), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n609), .A2(new_n619), .ZN(G156));
  XNOR2_X1  g195(.A(KEYINPUT15), .B(G2435), .ZN(new_n621));
  INV_X1    g196(.A(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2427), .ZN(new_n624));
  INV_X1    g199(.A(G2430), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n626), .A2(KEYINPUT14), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT83), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  AND2_X1   g206(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n629), .A2(new_n631), .ZN(new_n633));
  XOR2_X1   g208(.A(G2443), .B(G2446), .Z(new_n634));
  OR3_X1    g209(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n632), .B2(new_n633), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G14), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n638), .B1(new_n635), .B2(new_n636), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n640), .A2(new_n641), .ZN(G401));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  NOR3_X1   g222(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT18), .ZN(new_n649));
  INV_X1    g224(.A(new_n645), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n650), .A2(KEYINPUT17), .A3(new_n643), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n643), .B1(new_n650), .B2(KEYINPUT17), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n651), .B1(new_n652), .B2(new_n647), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n644), .A2(new_n647), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n650), .B1(new_n654), .B2(KEYINPUT17), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n649), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(new_n618), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(new_n608), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G227));
  XOR2_X1   g234(.A(G1971), .B(G1976), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1956), .B(G2474), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1961), .B(G1966), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  NOR3_X1   g240(.A1(new_n661), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n661), .A2(new_n664), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT20), .Z(new_n668));
  AOI211_X1 g243(.A(new_n666), .B(new_n668), .C1(new_n661), .C2(new_n665), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1981), .B(G1986), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT84), .ZN(new_n673));
  XOR2_X1   g248(.A(G1991), .B(G1996), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n671), .B(new_n675), .ZN(G229));
  NOR2_X1   g251(.A1(G16), .A2(G24), .ZN(new_n677));
  INV_X1    g252(.A(G290), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n677), .B1(new_n678), .B2(G16), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G1986), .ZN(new_n680));
  MUX2_X1   g255(.A(G95), .B(G107), .S(G2105), .Z(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G2104), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT86), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(new_n488), .B2(G119), .ZN(new_n684));
  AND3_X1   g259(.A1(new_n492), .A2(KEYINPUT85), .A3(G131), .ZN(new_n685));
  AOI21_X1  g260(.A(KEYINPUT85), .B1(new_n492), .B2(G131), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  MUX2_X1   g262(.A(G25), .B(new_n687), .S(G29), .Z(new_n688));
  XOR2_X1   g263(.A(KEYINPUT35), .B(G1991), .Z(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n688), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT34), .ZN(new_n692));
  NOR2_X1   g267(.A1(G16), .A2(G22), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(G166), .B2(G16), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1971), .ZN(new_n695));
  NOR2_X1   g270(.A1(G6), .A2(G16), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n575), .B2(G16), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT32), .B(G1981), .Z(new_n698));
  XOR2_X1   g273(.A(new_n697), .B(new_n698), .Z(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G23), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n568), .B2(new_n700), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT33), .B(G1976), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n702), .B(new_n703), .Z(new_n704));
  NOR3_X1   g279(.A1(new_n695), .A2(new_n699), .A3(new_n704), .ZN(new_n705));
  AOI211_X1 g280(.A(new_n680), .B(new_n691), .C1(new_n692), .C2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT87), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n705), .A2(new_n692), .ZN(new_n708));
  OR3_X1    g283(.A1(new_n707), .A2(KEYINPUT36), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(KEYINPUT36), .B1(new_n707), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(G4), .A2(G16), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT88), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n589), .B2(new_n700), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT90), .B(G1348), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT89), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n714), .B(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(KEYINPUT30), .A2(G28), .ZN(new_n718));
  NAND2_X1  g293(.A1(KEYINPUT30), .A2(G28), .ZN(new_n719));
  AOI21_X1  g294(.A(G29), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT31), .B(G11), .Z(new_n721));
  NOR2_X1   g296(.A1(G168), .A2(new_n700), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n700), .B2(G21), .ZN(new_n723));
  INV_X1    g298(.A(G1966), .ZN(new_n724));
  AOI211_X1 g299(.A(new_n720), .B(new_n721), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n617), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n723), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(G1966), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n700), .A2(G19), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT91), .Z(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n544), .B2(new_n700), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(G1341), .Z(new_n733));
  NAND3_X1  g308(.A1(new_n725), .A2(new_n729), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G2084), .ZN(new_n735));
  NAND2_X1  g310(.A1(G160), .A2(G29), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT24), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n726), .B1(new_n737), .B2(G34), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(KEYINPUT95), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(KEYINPUT95), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n737), .A2(G34), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n736), .A2(new_n742), .ZN(new_n743));
  AOI211_X1 g318(.A(new_n717), .B(new_n734), .C1(new_n735), .C2(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(G29), .A2(G35), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G162), .B2(G29), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT97), .B(KEYINPUT29), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G2090), .ZN(new_n749));
  NOR2_X1   g324(.A1(G27), .A2(G29), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G164), .B2(G29), .ZN(new_n751));
  INV_X1    g326(.A(G2078), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n744), .A2(new_n749), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n743), .A2(new_n735), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n492), .A2(G141), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n488), .A2(G129), .ZN(new_n757));
  NAND3_X1  g332(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT26), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n760), .A2(new_n761), .B1(G105), .B2(new_n482), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n756), .A2(new_n757), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(new_n726), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n726), .B2(G32), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT27), .B(G1996), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n726), .A2(G26), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT28), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n488), .A2(G128), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n492), .A2(G140), .ZN(new_n771));
  MUX2_X1   g346(.A(G104), .B(G116), .S(G2105), .Z(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G2104), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT92), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n770), .A2(new_n771), .A3(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n769), .B1(new_n776), .B2(new_n726), .ZN(new_n777));
  OAI22_X1  g352(.A1(new_n766), .A2(new_n767), .B1(G2067), .B2(new_n777), .ZN(new_n778));
  AOI211_X1 g353(.A(new_n755), .B(new_n778), .C1(new_n766), .C2(new_n767), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n726), .A2(G33), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n492), .A2(G139), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT94), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT93), .B(KEYINPUT25), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n482), .A2(G103), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n603), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(new_n480), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n780), .B1(new_n788), .B2(new_n726), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(G2072), .Z(new_n790));
  NAND2_X1  g365(.A1(new_n700), .A2(G20), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT23), .Z(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G299), .B2(G16), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(G1956), .Z(new_n794));
  NAND2_X1  g369(.A1(G171), .A2(G16), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G5), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT96), .ZN(new_n797));
  INV_X1    g372(.A(G1961), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n797), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n800), .A2(G1961), .B1(G2067), .B2(new_n777), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n779), .A2(new_n790), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n748), .A2(G2090), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n754), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n711), .A2(new_n804), .ZN(G311));
  NAND2_X1  g380(.A1(new_n711), .A2(new_n804), .ZN(G150));
  AOI22_X1  g381(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(new_n516), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT98), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n521), .A2(G55), .B1(G93), .B2(new_n514), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(G860), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT37), .Z(new_n814));
  INV_X1    g389(.A(new_n812), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(new_n544), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n812), .A2(new_n543), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT38), .Z(new_n819));
  NOR2_X1   g394(.A1(new_n589), .A2(new_n598), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n822), .A2(KEYINPUT39), .ZN(new_n823));
  INV_X1    g398(.A(G860), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n822), .B2(KEYINPUT39), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n814), .B1(new_n823), .B2(new_n825), .ZN(G145));
  NAND2_X1  g401(.A1(new_n788), .A2(new_n764), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n763), .B1(new_n782), .B2(new_n787), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n830));
  INV_X1    g405(.A(new_n501), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT99), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n507), .B1(new_n503), .B2(KEYINPUT99), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n775), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n829), .B(new_n837), .ZN(new_n838));
  MUX2_X1   g413(.A(G106), .B(G118), .S(G2105), .Z(new_n839));
  AOI22_X1  g414(.A1(new_n488), .A2(G130), .B1(G2104), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n492), .A2(G142), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n687), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n606), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n838), .A2(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n829), .A2(new_n837), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n829), .A2(new_n837), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n847), .A2(new_n844), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n617), .B(G160), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n495), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n846), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n846), .A2(new_n849), .A3(KEYINPUT101), .A4(new_n851), .ZN(new_n855));
  AOI21_X1  g430(.A(G37), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n851), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n846), .A2(KEYINPUT100), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(new_n849), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n846), .A2(KEYINPUT100), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g438(.A(new_n568), .ZN(new_n864));
  XNOR2_X1  g439(.A(G290), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(G166), .B(new_n575), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(KEYINPUT102), .B1(new_n865), .B2(new_n866), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n869), .A2(new_n870), .B1(new_n865), .B2(new_n866), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT42), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n597), .B(G299), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT41), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n589), .B(G299), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT41), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n818), .B(new_n600), .ZN(new_n879));
  MUX2_X1   g454(.A(new_n878), .B(new_n873), .S(new_n879), .Z(new_n880));
  AND2_X1   g455(.A1(new_n872), .A2(new_n880), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n881), .A2(KEYINPUT103), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(KEYINPUT103), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n882), .B(new_n883), .C1(new_n880), .C2(new_n872), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(G868), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(G868), .B2(new_n815), .ZN(G295));
  OAI21_X1  g461(.A(new_n885), .B1(G868), .B2(new_n815), .ZN(G331));
  NAND2_X1  g462(.A1(G301), .A2(KEYINPUT104), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n889));
  NAND2_X1  g464(.A1(G171), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n890), .A3(G168), .ZN(new_n891));
  NAND3_X1  g466(.A1(G286), .A2(KEYINPUT104), .A3(G301), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n818), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT105), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n893), .A2(new_n818), .ZN(new_n896));
  AOI22_X1  g471(.A1(new_n891), .A2(new_n892), .B1(new_n816), .B2(new_n817), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n895), .A2(new_n896), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n874), .A2(new_n877), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n893), .A2(new_n818), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n902), .A2(new_n897), .ZN(new_n903));
  OAI22_X1  g478(.A1(new_n900), .A2(new_n875), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n871), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT106), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n904), .A2(new_n907), .A3(new_n871), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n902), .A2(new_n875), .A3(new_n897), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n909), .B1(new_n900), .B2(new_n878), .ZN(new_n910));
  INV_X1    g485(.A(new_n871), .ZN(new_n911));
  AOI21_X1  g486(.A(G37), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n906), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n902), .B1(KEYINPUT105), .B2(new_n894), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n901), .B1(new_n916), .B2(new_n899), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n871), .B1(new_n917), .B2(new_n909), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n912), .A2(KEYINPUT43), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n915), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n912), .A2(new_n914), .A3(new_n918), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n922), .A2(KEYINPUT44), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n912), .A2(new_n908), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n907), .B1(new_n904), .B2(new_n871), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n924), .B(KEYINPUT43), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n924), .B1(new_n913), .B2(KEYINPUT43), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n921), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n921), .B(KEYINPUT108), .C1(new_n928), .C2(new_n929), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(G397));
  INV_X1    g509(.A(G1384), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n830), .A2(KEYINPUT99), .A3(new_n831), .ZN(new_n936));
  INV_X1    g511(.A(new_n507), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n503), .A2(KEYINPUT99), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n470), .A2(G40), .A3(new_n481), .A4(new_n484), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(G290), .A2(G1986), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n947), .A2(KEYINPUT48), .ZN(new_n948));
  INV_X1    g523(.A(G2067), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n775), .B(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G1996), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n763), .B(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n687), .B(new_n690), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n944), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n947), .A2(KEYINPUT48), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n948), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n944), .A2(new_n951), .ZN(new_n958));
  XOR2_X1   g533(.A(new_n958), .B(KEYINPUT46), .Z(new_n959));
  NAND2_X1  g534(.A1(new_n950), .A2(new_n764), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n959), .B1(new_n944), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT47), .ZN(new_n962));
  OR2_X1    g537(.A1(new_n687), .A2(new_n690), .ZN(new_n963));
  OAI22_X1  g538(.A1(new_n953), .A2(new_n963), .B1(G2067), .B2(new_n775), .ZN(new_n964));
  AOI211_X1 g539(.A(new_n957), .B(new_n962), .C1(new_n944), .C2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n935), .B1(new_n503), .B2(new_n507), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT50), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n943), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n940), .A2(KEYINPUT110), .A3(KEYINPUT50), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n973));
  AOI21_X1  g548(.A(G1384), .B1(new_n834), .B2(new_n835), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n735), .B(new_n971), .C1(new_n972), .C2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n943), .ZN(new_n980));
  OAI211_X1 g555(.A(KEYINPUT115), .B(new_n980), .C1(new_n974), .C2(KEYINPUT45), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT116), .ZN(new_n982));
  OR3_X1    g557(.A1(new_n966), .A2(new_n982), .A3(new_n941), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n982), .B1(new_n966), .B2(new_n941), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT115), .B1(new_n942), .B2(new_n980), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n724), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT110), .B1(new_n940), .B2(KEYINPUT50), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n974), .A2(new_n973), .A3(new_n975), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n991), .A2(KEYINPUT117), .A3(new_n735), .A4(new_n971), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n979), .A2(new_n988), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G2090), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n994), .B(new_n971), .C1(new_n972), .C2(new_n976), .ZN(new_n995));
  OAI211_X1 g570(.A(KEYINPUT45), .B(new_n935), .C1(new_n938), .C2(new_n939), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n943), .B1(new_n966), .B2(new_n941), .ZN(new_n997));
  AOI21_X1  g572(.A(G1971), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(G8), .B1(KEYINPUT112), .B2(KEYINPUT55), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(KEYINPUT112), .A2(KEYINPUT55), .ZN(new_n1003));
  AND3_X1   g578(.A1(G303), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1003), .B1(G303), .B2(new_n1002), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1000), .A2(G8), .A3(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n935), .B(new_n980), .C1(new_n938), .C2(new_n939), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n568), .A2(G1976), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(G8), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT52), .ZN(new_n1011));
  OAI21_X1  g586(.A(G1981), .B1(new_n572), .B2(new_n574), .ZN(new_n1012));
  INV_X1    g587(.A(new_n574), .ZN(new_n1013));
  INV_X1    g588(.A(G1981), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1013), .A2(new_n1014), .A3(new_n570), .A4(new_n571), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT49), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1017), .A2(G8), .A3(new_n1008), .ZN(new_n1018));
  INV_X1    g593(.A(G1976), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT52), .B1(G288), .B2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1020), .A2(new_n1008), .A3(G8), .A4(new_n1009), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1011), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  OAI211_X1 g597(.A(KEYINPUT50), .B(new_n935), .C1(new_n938), .C2(new_n939), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n966), .A2(new_n975), .ZN(new_n1024));
  AOI211_X1 g599(.A(G2090), .B(new_n943), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(G8), .B1(new_n1025), .B2(new_n998), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1006), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1022), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G8), .ZN(new_n1029));
  NOR2_X1   g604(.A1(G286), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n993), .A2(new_n1007), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT63), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT118), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1031), .A2(new_n1035), .A3(new_n1032), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n993), .A2(new_n1030), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1007), .A2(KEYINPUT63), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1000), .A2(G8), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n1027), .ZN(new_n1040));
  XOR2_X1   g615(.A(new_n1022), .B(KEYINPUT113), .Z(new_n1041));
  NAND4_X1  g616(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1034), .A2(new_n1036), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1007), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1008), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1045), .A2(new_n1029), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1015), .B(KEYINPUT114), .ZN(new_n1047));
  OR2_X1    g622(.A1(G288), .A2(G1976), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1047), .B1(new_n1048), .B2(new_n1017), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n1041), .A2(new_n1044), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n979), .A2(new_n988), .A3(G168), .A4(new_n992), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(G8), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT51), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT62), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n993), .B2(G286), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1053), .B(new_n1054), .C1(new_n1052), .C2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT123), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n996), .A2(new_n752), .A3(new_n997), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1059), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n966), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT111), .B1(new_n966), .B2(KEYINPUT50), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n980), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(new_n989), .B2(new_n990), .ZN(new_n1066));
  OAI22_X1  g641(.A1(new_n1061), .A2(new_n1062), .B1(new_n1066), .B2(G1961), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1060), .A2(G2078), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n986), .A2(new_n987), .A3(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(G171), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1007), .A2(new_n1028), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1057), .A2(new_n1073), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1051), .A2(G8), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n993), .A2(G286), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1075), .B1(new_n1076), .B2(new_n1055), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1054), .B1(new_n1077), .B2(new_n1053), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1043), .B(new_n1050), .C1(new_n1074), .C2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(G301), .ZN(new_n1082));
  AND4_X1   g657(.A1(new_n980), .A2(new_n942), .A3(new_n996), .A4(new_n1068), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT123), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1059), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n1066), .B2(G1961), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n991), .A2(new_n971), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1090), .A2(KEYINPUT124), .A3(new_n798), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1087), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT125), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1092), .A2(new_n1093), .A3(G171), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1093), .B1(new_n1092), .B2(G171), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1082), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1053), .B1(new_n1052), .B2(new_n1056), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1087), .A2(new_n1089), .A3(new_n1091), .A4(G301), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1071), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1072), .B1(new_n1099), .B2(new_n1080), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1096), .A2(new_n1097), .A3(new_n1100), .A4(KEYINPUT126), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1090), .A2(new_n715), .B1(new_n949), .B2(new_n1045), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1102), .A2(new_n589), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n943), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(G1956), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT56), .B(G2072), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n996), .A2(new_n997), .A3(new_n1107), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n1108), .A2(KEYINPUT120), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n1110));
  NOR3_X1   g685(.A1(G299), .A2(new_n1110), .A3(KEYINPUT57), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1111), .B1(G299), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1108), .A2(KEYINPUT120), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1106), .A2(new_n1109), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1103), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1113), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1109), .A2(new_n1114), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1117), .B1(new_n1118), .B2(new_n1105), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1102), .A2(new_n589), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT60), .B1(new_n1121), .B2(new_n1103), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n996), .A2(new_n951), .A3(new_n997), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT58), .B(G1341), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1123), .B1(new_n1045), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1125), .A2(KEYINPUT122), .A3(new_n544), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1128), .A2(KEYINPUT121), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT122), .B1(new_n1125), .B2(new_n544), .ZN(new_n1130));
  OR3_X1    g705(.A1(new_n1127), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1129), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1119), .A2(KEYINPUT61), .A3(new_n1115), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1122), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT60), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1102), .A2(new_n1136), .A3(new_n597), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1119), .A2(new_n1115), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1137), .B1(new_n1138), .B2(KEYINPUT61), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1120), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1101), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1096), .A2(new_n1097), .A3(new_n1100), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT126), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1079), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  AND2_X1   g720(.A1(G290), .A2(G1986), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n944), .B1(new_n945), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT109), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1149), .A2(new_n1150), .A3(new_n955), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n965), .B1(new_n1145), .B2(new_n1151), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g727(.A1(new_n658), .A2(G319), .ZN(new_n1154));
  NOR2_X1   g728(.A1(G229), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g729(.A(new_n1155), .B1(new_n640), .B2(new_n641), .ZN(new_n1156));
  AOI21_X1  g730(.A(new_n1156), .B1(new_n856), .B2(new_n861), .ZN(new_n1157));
  INV_X1    g731(.A(new_n919), .ZN(new_n1158));
  AOI21_X1  g732(.A(new_n1158), .B1(new_n914), .B2(new_n913), .ZN(new_n1159));
  AND3_X1   g733(.A1(new_n1157), .A2(new_n1159), .A3(KEYINPUT127), .ZN(new_n1160));
  AOI21_X1  g734(.A(KEYINPUT127), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1161));
  NOR2_X1   g735(.A1(new_n1160), .A2(new_n1161), .ZN(G308));
  NAND2_X1  g736(.A1(new_n1157), .A2(new_n1159), .ZN(G225));
endmodule


