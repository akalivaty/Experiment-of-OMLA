//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(KEYINPUT87), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(KEYINPUT87), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(KEYINPUT15), .A3(new_n204), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n206));
  XNOR2_X1  g005(.A(KEYINPUT89), .B(G29gat), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NOR3_X1   g010(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n205), .B(new_n206), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n212), .A2(KEYINPUT88), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n210), .B1(new_n212), .B2(KEYINPUT88), .ZN(new_n215));
  OAI22_X1  g014(.A1(new_n214), .A2(new_n215), .B1(new_n208), .B2(new_n207), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n216), .A2(KEYINPUT15), .A3(new_n203), .A4(new_n204), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT17), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G15gat), .B(G22gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT16), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n221), .B1(new_n222), .B2(G1gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n223), .B(new_n224), .C1(G1gat), .C2(new_n221), .ZN(new_n225));
  NOR2_X1   g024(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n213), .A2(new_n217), .A3(KEYINPUT17), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n220), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n227), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n218), .ZN(new_n231));
  NAND2_X1  g030(.A1(G229gat), .A2(G233gat), .ZN(new_n232));
  XOR2_X1   g031(.A(new_n232), .B(KEYINPUT91), .Z(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n229), .A2(KEYINPUT18), .A3(new_n231), .A4(new_n234), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n233), .B(KEYINPUT13), .Z(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n230), .A2(new_n218), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n227), .B1(new_n217), .B2(new_n213), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n229), .A2(new_n231), .A3(new_n234), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT18), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT92), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n235), .A2(new_n240), .A3(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G113gat), .B(G141gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(G197gat), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT11), .B(G169gat), .Z(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT12), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n245), .A2(new_n247), .A3(new_n253), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n241), .B(new_n244), .C1(new_n246), .C2(new_n252), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(G57gat), .B(G64gat), .Z(new_n257));
  INV_X1    g056(.A(KEYINPUT9), .ZN(new_n258));
  INV_X1    g057(.A(G71gat), .ZN(new_n259));
  INV_X1    g058(.A(G78gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G71gat), .B(G78gat), .Z(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT21), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G231gat), .A2(G233gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G127gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n227), .B1(new_n265), .B2(new_n264), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT93), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(G155gat), .ZN(new_n275));
  XOR2_X1   g074(.A(G183gat), .B(G211gat), .Z(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n272), .B(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G134gat), .B(G162gat), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G99gat), .A2(G106gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT8), .ZN(new_n283));
  OR2_X1    g082(.A1(G85gat), .A2(G92gat), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n283), .A2(KEYINPUT94), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT94), .B1(new_n283), .B2(new_n284), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT95), .ZN(new_n288));
  XOR2_X1   g087(.A(G99gat), .B(G106gat), .Z(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G85gat), .A2(G92gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT7), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n287), .A2(new_n288), .A3(new_n290), .A4(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n292), .B1(new_n285), .B2(new_n286), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(new_n289), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n290), .B(new_n292), .C1(new_n285), .C2(new_n286), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(KEYINPUT95), .A3(new_n296), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n220), .A2(new_n228), .A3(new_n293), .A4(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G190gat), .B(G218gat), .ZN(new_n299));
  XOR2_X1   g098(.A(new_n299), .B(KEYINPUT96), .Z(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(new_n293), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n218), .ZN(new_n303));
  NAND3_X1  g102(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n298), .A2(new_n301), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n281), .B1(new_n306), .B2(KEYINPUT97), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n298), .A2(new_n303), .A3(new_n304), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n300), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT97), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(new_n310), .A3(new_n305), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n309), .A2(new_n281), .A3(new_n305), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT98), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n309), .A2(KEYINPUT98), .A3(new_n281), .A4(new_n305), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n312), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n278), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G120gat), .B(G148gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(G176gat), .B(G204gat), .ZN(new_n321));
  XOR2_X1   g120(.A(new_n320), .B(new_n321), .Z(new_n322));
  XNOR2_X1  g121(.A(new_n322), .B(KEYINPUT100), .ZN(new_n323));
  NAND2_X1  g122(.A1(G230gat), .A2(G233gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n297), .A2(new_n264), .A3(new_n293), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT99), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n297), .A2(KEYINPUT99), .A3(new_n264), .A4(new_n293), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT10), .ZN(new_n331));
  INV_X1    g130(.A(new_n264), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n332), .A2(new_n296), .A3(new_n295), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n330), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n302), .A2(KEYINPUT10), .A3(new_n332), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n325), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n333), .B1(new_n328), .B2(new_n329), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n338), .A2(new_n324), .ZN(new_n339));
  OAI211_X1 g138(.A(KEYINPUT101), .B(new_n323), .C1(new_n337), .C2(new_n339), .ZN(new_n340));
  AOI211_X1 g139(.A(KEYINPUT10), .B(new_n333), .C1(new_n328), .C2(new_n329), .ZN(new_n341));
  INV_X1    g140(.A(new_n336), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n324), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OR2_X1    g142(.A1(new_n338), .A2(new_n324), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(new_n344), .A3(new_n322), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n342), .B1(new_n338), .B2(new_n331), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n344), .B1(new_n347), .B2(new_n325), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT101), .B1(new_n348), .B2(new_n323), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n319), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT36), .ZN(new_n353));
  XNOR2_X1  g152(.A(G15gat), .B(G43gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT68), .ZN(new_n355));
  XNOR2_X1  g154(.A(G71gat), .B(G99gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G183gat), .A2(G190gat), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G169gat), .ZN(new_n360));
  INV_X1    g159(.A(G176gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(G169gat), .A2(G176gat), .ZN(new_n363));
  NOR3_X1   g162(.A1(new_n362), .A2(KEYINPUT26), .A3(new_n363), .ZN(new_n364));
  AOI211_X1 g163(.A(new_n359), .B(new_n364), .C1(KEYINPUT26), .C2(new_n363), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT28), .ZN(new_n366));
  NOR2_X1   g165(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT64), .B(G183gat), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n367), .B1(new_n368), .B2(KEYINPUT27), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n366), .B1(new_n369), .B2(G190gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT27), .B(G183gat), .ZN(new_n371));
  INV_X1    g170(.A(G190gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(KEYINPUT28), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n365), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT25), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n363), .A2(KEYINPUT23), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT23), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n378), .B1(G169gat), .B2(G176gat), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n377), .B(new_n379), .C1(new_n360), .C2(new_n361), .ZN(new_n380));
  NOR2_X1   g179(.A1(G183gat), .A2(G190gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n358), .A2(KEYINPUT24), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT24), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(G183gat), .A3(G190gat), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n381), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n376), .B1(new_n380), .B2(new_n385), .ZN(new_n386));
  OR2_X1    g185(.A1(new_n380), .A2(new_n376), .ZN(new_n387));
  INV_X1    g186(.A(new_n368), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n388), .A2(new_n372), .B1(new_n384), .B2(new_n382), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n386), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(G113gat), .ZN(new_n392));
  INV_X1    g191(.A(G120gat), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT1), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n394), .B1(new_n392), .B2(new_n393), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT65), .ZN(new_n396));
  XNOR2_X1  g195(.A(G127gat), .B(G134gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n391), .B(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(G227gat), .A3(G233gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT32), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n357), .B1(new_n401), .B2(KEYINPUT67), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n402), .B1(KEYINPUT67), .B2(new_n401), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT33), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT66), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n357), .A2(new_n404), .ZN(new_n408));
  OAI22_X1  g207(.A1(new_n403), .A2(new_n407), .B1(new_n401), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n399), .B1(G227gat), .B2(G233gat), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n409), .B(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n413));
  AND2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n412), .A2(new_n413), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n353), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT83), .ZN(new_n417));
  XNOR2_X1  g216(.A(G1gat), .B(G29gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(KEYINPUT0), .ZN(new_n419));
  XNOR2_X1  g218(.A(G57gat), .B(G85gat), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n419), .B(new_n420), .Z(new_n421));
  XOR2_X1   g220(.A(G141gat), .B(G148gat), .Z(new_n422));
  INV_X1    g221(.A(KEYINPUT2), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G155gat), .B(G162gat), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT74), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT74), .B1(G155gat), .B2(G162gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT75), .B(G162gat), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n423), .B1(new_n430), .B2(G155gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n422), .A2(new_n425), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n429), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n398), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(KEYINPUT4), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT78), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n434), .A2(new_n436), .A3(KEYINPUT4), .ZN(new_n438));
  OR2_X1    g237(.A1(new_n433), .A2(KEYINPUT3), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n433), .A2(KEYINPUT3), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(new_n398), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  OR2_X1    g241(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(G225gat), .A2(G233gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n444), .B(KEYINPUT76), .Z(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n421), .B1(new_n446), .B2(KEYINPUT39), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n398), .B(new_n433), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT39), .B1(new_n448), .B2(new_n445), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n443), .B2(new_n445), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n417), .B1(new_n451), .B2(KEYINPUT40), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT40), .ZN(new_n453));
  OAI211_X1 g252(.A(KEYINPUT83), .B(new_n453), .C1(new_n447), .C2(new_n450), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT79), .ZN(new_n456));
  INV_X1    g255(.A(new_n445), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT5), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n456), .B1(new_n443), .B2(new_n459), .ZN(new_n460));
  OR4_X1    g259(.A1(new_n456), .A2(new_n437), .A3(new_n442), .A4(new_n459), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n435), .A2(new_n457), .A3(new_n441), .ZN(new_n463));
  XOR2_X1   g262(.A(new_n463), .B(KEYINPUT77), .Z(new_n464));
  AOI21_X1  g263(.A(new_n458), .B1(new_n448), .B2(new_n445), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n421), .ZN(new_n468));
  AOI22_X1  g267(.A1(KEYINPUT40), .A2(new_n451), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT29), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n391), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(G226gat), .A2(G233gat), .ZN(new_n472));
  MUX2_X1   g271(.A(new_n391), .B(new_n471), .S(new_n472), .Z(new_n473));
  XNOR2_X1  g272(.A(G197gat), .B(G204gat), .ZN(new_n474));
  INV_X1    g273(.A(G211gat), .ZN(new_n475));
  INV_X1    g274(.A(G218gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n474), .B1(KEYINPUT22), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(G211gat), .B(G218gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  XOR2_X1   g279(.A(new_n480), .B(KEYINPUT70), .Z(new_n481));
  OR2_X1    g280(.A1(new_n473), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n473), .A2(new_n481), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G8gat), .B(G36gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(KEYINPUT71), .ZN(new_n486));
  XOR2_X1   g285(.A(G64gat), .B(G92gat), .Z(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n484), .A2(KEYINPUT30), .A3(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n489), .A2(KEYINPUT73), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n489), .A2(KEYINPUT73), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n488), .B(KEYINPUT72), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT30), .B1(new_n484), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n484), .A2(new_n488), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n490), .B1(new_n491), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n455), .A2(new_n469), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT82), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n439), .A2(new_n470), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT3), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(new_n480), .B2(KEYINPUT29), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n481), .A2(new_n500), .B1(new_n433), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT81), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n499), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n505), .B(G22gat), .Z(new_n506));
  OAI211_X1 g305(.A(G228gat), .B(G233gat), .C1(new_n503), .C2(new_n499), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n507), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G78gat), .B(G106gat), .ZN(new_n511));
  INV_X1    g310(.A(G50gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n508), .A2(new_n515), .A3(new_n509), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n467), .A2(new_n468), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT6), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n462), .A2(new_n466), .A3(new_n421), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n467), .A2(KEYINPUT6), .A3(new_n468), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n482), .A2(new_n483), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n525), .A2(KEYINPUT37), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT85), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT38), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n492), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT84), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n482), .A2(new_n530), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n531), .A2(KEYINPUT37), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n484), .A2(new_n530), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n529), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n527), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n523), .A2(new_n524), .A3(new_n495), .A4(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n488), .B1(new_n525), .B2(KEYINPUT37), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n528), .B1(new_n527), .B2(new_n537), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n498), .B(new_n519), .C1(new_n536), .C2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n497), .B1(new_n523), .B2(new_n524), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n540), .A2(new_n519), .ZN(new_n541));
  INV_X1    g340(.A(new_n413), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n409), .A2(new_n410), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n409), .A2(new_n410), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n412), .A2(new_n413), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(KEYINPUT36), .A3(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n416), .A2(new_n539), .A3(new_n541), .A4(new_n548), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n519), .B(new_n540), .C1(new_n414), .C2(new_n415), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n550), .A2(KEYINPUT35), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT35), .ZN(new_n552));
  INV_X1    g351(.A(new_n519), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n553), .B1(new_n546), .B2(new_n547), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n552), .B1(new_n554), .B2(new_n540), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n549), .B(KEYINPUT86), .C1(new_n551), .C2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n550), .A2(KEYINPUT35), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n554), .A2(new_n552), .A3(new_n540), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT86), .B1(new_n560), .B2(new_n549), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n256), .B(new_n352), .C1(new_n557), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n523), .A2(new_n524), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n564), .B(G1gat), .Z(G1324gat));
  INV_X1    g364(.A(new_n497), .ZN(new_n566));
  XOR2_X1   g365(.A(KEYINPUT16), .B(G8gat), .Z(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n562), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n569), .A2(KEYINPUT104), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT104), .ZN(new_n571));
  INV_X1    g370(.A(new_n256), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n549), .B1(new_n551), .B2(new_n555), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT86), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n572), .B1(new_n575), .B2(new_n556), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n576), .A2(new_n497), .A3(new_n352), .A4(new_n567), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n571), .B1(new_n577), .B2(KEYINPUT102), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT42), .B1(new_n570), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT102), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT104), .B1(new_n569), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT42), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(G8gat), .B1(new_n562), .B2(new_n566), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT103), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n579), .A2(new_n583), .A3(new_n585), .ZN(G1325gat));
  NAND2_X1  g385(.A1(new_n416), .A2(new_n548), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(G15gat), .B1(new_n562), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n546), .A2(new_n547), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n591), .A2(G15gat), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n589), .B1(new_n562), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT105), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(G1326gat));
  OR3_X1    g394(.A1(new_n562), .A2(KEYINPUT106), .A3(new_n519), .ZN(new_n596));
  OAI21_X1  g395(.A(KEYINPUT106), .B1(new_n562), .B2(new_n519), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT43), .B(G22gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(G1327gat));
  NOR3_X1   g402(.A1(new_n351), .A2(new_n278), .A3(new_n318), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT107), .ZN(new_n605));
  AOI211_X1 g404(.A(new_n572), .B(new_n605), .C1(new_n575), .C2(new_n556), .ZN(new_n606));
  INV_X1    g405(.A(new_n563), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n606), .A2(new_n607), .A3(new_n207), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT45), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT44), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n318), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n557), .B2(new_n561), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n573), .A2(new_n317), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n610), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n350), .B(KEYINPUT108), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n617), .A2(new_n572), .A3(new_n278), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n615), .A2(new_n607), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n609), .B1(new_n207), .B2(new_n619), .ZN(G1328gat));
  NAND4_X1  g419(.A1(new_n612), .A2(new_n497), .A3(new_n614), .A4(new_n618), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(G36gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n605), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n576), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n566), .A2(G36gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(KEYINPUT46), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT46), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n606), .A2(new_n628), .A3(new_n625), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n622), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT109), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n622), .A2(new_n627), .A3(KEYINPUT109), .A4(new_n629), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(G1329gat));
  NAND4_X1  g433(.A1(new_n612), .A2(new_n587), .A3(new_n614), .A4(new_n618), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(G43gat), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT47), .ZN(new_n637));
  INV_X1    g436(.A(G43gat), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n606), .A2(new_n638), .A3(new_n590), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n637), .B1(new_n636), .B2(new_n639), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(G1330gat));
  NAND4_X1  g441(.A1(new_n612), .A2(new_n553), .A3(new_n614), .A4(new_n618), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(G50gat), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT110), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT48), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n606), .A2(new_n512), .A3(new_n553), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n644), .B(new_n647), .C1(new_n645), .C2(KEYINPUT48), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(G1331gat));
  NOR2_X1   g450(.A1(new_n319), .A2(new_n256), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n617), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT111), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n573), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n607), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G57gat), .ZN(G1332gat));
  INV_X1    g456(.A(new_n655), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n658), .A2(new_n566), .ZN(new_n659));
  NOR2_X1   g458(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n660));
  AND2_X1   g459(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n659), .B2(new_n660), .ZN(G1333gat));
  NAND3_X1  g462(.A1(new_n655), .A2(G71gat), .A3(new_n587), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT112), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n259), .B1(new_n658), .B2(new_n591), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(G1334gat));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n553), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g473(.A1(new_n278), .A2(new_n256), .A3(new_n350), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n612), .A2(new_n607), .A3(new_n614), .A4(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(G85gat), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n563), .A2(G85gat), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n318), .B1(new_n560), .B2(new_n549), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n278), .A2(new_n256), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n679), .A2(KEYINPUT51), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT51), .B1(new_n679), .B2(new_n680), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n351), .B(new_n678), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT114), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n677), .A2(KEYINPUT114), .A3(new_n683), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(G1336gat));
  NAND4_X1  g487(.A1(new_n612), .A2(new_n497), .A3(new_n614), .A4(new_n675), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(G92gat), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n681), .A2(new_n682), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n566), .A2(new_n616), .A3(G92gat), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n690), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT52), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT52), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n690), .B(new_n696), .C1(new_n691), .C2(new_n693), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(G1337gat));
  OR4_X1    g497(.A1(G99gat), .A2(new_n691), .A3(new_n591), .A4(new_n350), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n615), .A2(new_n587), .A3(new_n675), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(G99gat), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(G1338gat));
  NAND4_X1  g501(.A1(new_n612), .A2(new_n553), .A3(new_n614), .A4(new_n675), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(G106gat), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT53), .ZN(new_n705));
  OR3_X1    g504(.A1(new_n519), .A2(G106gat), .A3(new_n616), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n704), .B(new_n705), .C1(new_n691), .C2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n691), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n706), .B(KEYINPUT115), .ZN(new_n709));
  AOI22_X1  g508(.A1(new_n708), .A2(new_n709), .B1(new_n703), .B2(G106gat), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n707), .B1(new_n705), .B2(new_n710), .ZN(G1339gat));
  INV_X1    g510(.A(new_n278), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT54), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n322), .B1(new_n337), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n335), .A2(new_n325), .A3(new_n336), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n343), .A2(new_n715), .A3(KEYINPUT54), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT55), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n241), .A2(new_n244), .A3(new_n252), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n234), .B1(new_n229), .B2(new_n231), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n238), .A2(new_n239), .A3(new_n237), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n251), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n719), .A2(new_n317), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n714), .A2(new_n716), .A3(KEYINPUT55), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n345), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT116), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n719), .A2(new_n256), .A3(new_n345), .A4(new_n726), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n724), .B1(new_n346), .B2(new_n349), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n317), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n712), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n652), .A2(new_n350), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n519), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n563), .A2(new_n497), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n590), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n392), .B1(new_n739), .B2(new_n256), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(KEYINPUT117), .Z(new_n741));
  INV_X1    g540(.A(new_n735), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n563), .ZN(new_n743));
  INV_X1    g542(.A(new_n554), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n497), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(new_n392), .A3(new_n256), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n741), .A2(new_n748), .ZN(G1340gat));
  AOI21_X1  g548(.A(G120gat), .B1(new_n747), .B2(new_n351), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n616), .A2(new_n393), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n739), .B2(new_n751), .ZN(G1341gat));
  INV_X1    g551(.A(new_n739), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n753), .A2(new_n269), .A3(new_n712), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n746), .A2(new_n712), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n755), .A2(KEYINPUT118), .ZN(new_n756));
  AOI21_X1  g555(.A(G127gat), .B1(new_n755), .B2(KEYINPUT118), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n754), .B1(new_n756), .B2(new_n757), .ZN(G1342gat));
  NOR3_X1   g557(.A1(new_n746), .A2(G134gat), .A3(new_n318), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n760), .A2(KEYINPUT56), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(KEYINPUT56), .ZN(new_n762));
  OAI21_X1  g561(.A(G134gat), .B1(new_n753), .B2(new_n318), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(G1343gat));
  NOR3_X1   g563(.A1(new_n587), .A2(new_n497), .A3(new_n519), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n743), .A2(new_n765), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n766), .A2(G141gat), .A3(new_n572), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n588), .A2(new_n737), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT57), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n742), .B2(new_n519), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n519), .A2(new_n769), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n731), .A2(KEYINPUT119), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT119), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n724), .B(new_n773), .C1(new_n346), .C2(new_n349), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n772), .A2(new_n730), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n318), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n729), .B1(KEYINPUT120), .B2(new_n776), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n776), .A2(KEYINPUT120), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n278), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n734), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n771), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n768), .B1(new_n770), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n256), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n767), .B1(new_n783), .B2(G141gat), .ZN(new_n784));
  XNOR2_X1  g583(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n784), .B(new_n785), .ZN(G1344gat));
  INV_X1    g585(.A(new_n766), .ZN(new_n787));
  INV_X1    g586(.A(G148gat), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(new_n788), .A3(new_n351), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT59), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n735), .A2(new_n771), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n728), .B1(new_n775), .B2(new_n318), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n734), .B1(new_n792), .B2(new_n278), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT122), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n519), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n734), .B(KEYINPUT122), .C1(new_n792), .C2(new_n278), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT57), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n791), .B1(new_n797), .B2(KEYINPUT123), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT123), .ZN(new_n799));
  AOI211_X1 g598(.A(new_n799), .B(KEYINPUT57), .C1(new_n795), .C2(new_n796), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n801), .A2(new_n588), .A3(new_n351), .A4(new_n737), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n790), .B1(new_n802), .B2(G148gat), .ZN(new_n803));
  AOI211_X1 g602(.A(KEYINPUT59), .B(new_n788), .C1(new_n782), .C2(new_n351), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n789), .B1(new_n803), .B2(new_n804), .ZN(G1345gat));
  INV_X1    g604(.A(G155gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n787), .A2(new_n806), .A3(new_n278), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n782), .A2(new_n278), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n807), .B1(new_n808), .B2(new_n806), .ZN(G1346gat));
  INV_X1    g608(.A(new_n430), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n787), .A2(new_n810), .A3(new_n317), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n782), .A2(new_n317), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n811), .B1(new_n812), .B2(new_n810), .ZN(G1347gat));
  NOR2_X1   g612(.A1(new_n742), .A2(new_n607), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n744), .A2(new_n566), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(G169gat), .B1(new_n817), .B2(new_n256), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n590), .A2(new_n563), .A3(new_n497), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n736), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n572), .A2(new_n360), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n818), .B1(new_n820), .B2(new_n821), .ZN(G1348gat));
  INV_X1    g621(.A(new_n820), .ZN(new_n823));
  OAI21_X1  g622(.A(G176gat), .B1(new_n823), .B2(new_n616), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n351), .A2(new_n361), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n816), .B2(new_n825), .ZN(G1349gat));
  NAND3_X1  g625(.A1(new_n817), .A2(new_n371), .A3(new_n278), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n368), .B1(new_n823), .B2(new_n712), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT60), .ZN(G1350gat));
  NOR3_X1   g629(.A1(new_n816), .A2(G190gat), .A3(new_n318), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(KEYINPUT124), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n372), .B1(new_n820), .B2(new_n317), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT61), .Z(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(G1351gat));
  NAND3_X1  g634(.A1(new_n588), .A2(new_n497), .A3(new_n553), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT125), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n814), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(G197gat), .B1(new_n839), .B2(new_n256), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n587), .A2(new_n607), .A3(new_n566), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n801), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n256), .A2(G197gat), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n840), .B1(new_n842), .B2(new_n843), .ZN(G1352gat));
  INV_X1    g643(.A(G204gat), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n837), .A2(new_n845), .A3(new_n351), .A4(new_n814), .ZN(new_n846));
  XOR2_X1   g645(.A(new_n846), .B(KEYINPUT62), .Z(new_n847));
  NAND2_X1  g646(.A1(new_n842), .A2(new_n617), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n847), .B1(new_n849), .B2(new_n845), .ZN(G1353gat));
  INV_X1    g649(.A(KEYINPUT127), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n278), .B(new_n841), .C1(new_n798), .C2(new_n800), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT126), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT63), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n852), .A2(G211gat), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n852), .B2(G211gat), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n853), .A2(new_n854), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n838), .A2(G211gat), .A3(new_n712), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n851), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n857), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n852), .A2(G211gat), .A3(new_n855), .ZN(new_n863));
  INV_X1    g662(.A(new_n858), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n839), .A2(new_n475), .A3(new_n278), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(KEYINPUT127), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n861), .A2(new_n867), .ZN(G1354gat));
  AOI21_X1  g667(.A(new_n476), .B1(new_n842), .B2(new_n317), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n838), .A2(G218gat), .A3(new_n318), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n869), .A2(new_n870), .ZN(G1355gat));
endmodule


