//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1285, new_n1286, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(KEYINPUT64), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT64), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n216), .A2(G1), .A3(G13), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n208), .ZN(new_n219));
  OAI21_X1  g0019(.A(G50), .B1(G58), .B2(G68), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(KEYINPUT66), .B(G244), .Z(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G77), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G97), .A2(G257), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT65), .Z(new_n231));
  OAI21_X1  g0031(.A(new_n210), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n213), .B(new_n222), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G226), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XOR2_X1   g0044(.A(G50), .B(G58), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  NAND2_X1  g0050(.A1(new_n204), .A2(G20), .ZN(new_n251));
  INV_X1    g0051(.A(G150), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT8), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G58), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI221_X1 g0061(.A(new_n251), .B1(new_n252), .B2(new_n254), .C1(new_n258), .C2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n218), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n262), .A2(new_n264), .B1(new_n201), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n264), .A2(new_n266), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n207), .A2(G20), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(G50), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n271), .B(KEYINPUT9), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G1), .A3(G13), .ZN(new_n277));
  AND3_X1   g0077(.A1(new_n275), .A2(new_n277), .A3(G274), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT67), .B(G226), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n278), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n215), .A2(new_n217), .A3(new_n276), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT3), .B(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G222), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G223), .A2(G1698), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n285), .B(new_n290), .C1(G77), .C2(new_n286), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n283), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G200), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(G190), .B2(new_n292), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n272), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(KEYINPUT10), .B1(new_n294), .B2(KEYINPUT70), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n296), .B(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n292), .A2(G169), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n292), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(new_n271), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n255), .A2(new_n257), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n269), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n268), .A2(new_n307), .B1(new_n266), .B2(new_n258), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  AOI22_X1  g0109(.A1(G33), .A2(new_n209), .B1(new_n215), .B2(new_n217), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n202), .A2(new_n203), .ZN(new_n311));
  NOR2_X1   g0111(.A1(G58), .A2(G68), .ZN(new_n312));
  OAI21_X1  g0112(.A(G20), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n253), .A2(G159), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT74), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT3), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n316), .B1(new_n317), .B2(G33), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(G33), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n259), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n208), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n203), .B1(new_n322), .B2(KEYINPUT7), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT7), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n321), .A2(new_n324), .A3(new_n208), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n315), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n310), .B1(new_n326), .B2(KEYINPUT16), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT16), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n324), .B1(new_n286), .B2(G20), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n319), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n203), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n328), .B1(new_n333), .B2(new_n315), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n309), .B1(new_n327), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(G223), .A2(G1698), .ZN(new_n336));
  INV_X1    g0136(.A(G226), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(G1698), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n338), .A2(new_n319), .A3(new_n318), .A4(new_n320), .ZN(new_n339));
  NAND2_X1  g0139(.A1(G33), .A2(G87), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n284), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n275), .A2(new_n277), .A3(G274), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n277), .A2(G232), .A3(new_n279), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(G169), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n337), .A2(G1698), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(G223), .B2(G1698), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n340), .B1(new_n321), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n344), .B1(new_n348), .B2(new_n285), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G179), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(KEYINPUT18), .B1(new_n335), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n322), .A2(KEYINPUT7), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(G68), .A3(new_n325), .ZN(new_n354));
  INV_X1    g0154(.A(new_n315), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(KEYINPUT16), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n356), .A2(new_n334), .A3(new_n264), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n351), .B1(new_n357), .B2(new_n308), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT18), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT17), .ZN(new_n361));
  INV_X1    g0161(.A(G190), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n349), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(G200), .B2(new_n349), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n361), .B1(new_n335), .B2(new_n364), .ZN(new_n365));
  AND4_X1   g0165(.A1(new_n361), .A2(new_n357), .A3(new_n308), .A4(new_n364), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n352), .B(new_n360), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT72), .B1(new_n265), .B2(G68), .ZN(new_n369));
  XOR2_X1   g0169(.A(new_n369), .B(KEYINPUT12), .Z(new_n370));
  NAND3_X1  g0170(.A1(new_n268), .A2(G68), .A3(new_n269), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n253), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n372));
  INV_X1    g0172(.A(G77), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n372), .B1(new_n261), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n264), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT11), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n374), .A2(KEYINPUT11), .A3(new_n264), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n370), .A2(new_n371), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT14), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G97), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n238), .A2(G1698), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(G226), .B2(G1698), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n381), .B1(new_n383), .B2(new_n331), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n278), .B1(new_n384), .B2(new_n285), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT13), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT71), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n280), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n277), .A2(KEYINPUT71), .A3(new_n279), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(G238), .A3(new_n389), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n385), .A2(new_n386), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n386), .B1(new_n385), .B2(new_n390), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n380), .B(G169), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(G226), .A2(G1698), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n394), .B1(new_n238), .B2(G1698), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n395), .A2(new_n286), .B1(G33), .B2(G97), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n342), .B1(new_n396), .B2(new_n284), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n388), .A2(G238), .A3(new_n389), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT13), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n385), .A2(new_n386), .A3(new_n390), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(G179), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n393), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n399), .A2(new_n400), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n380), .B1(new_n403), .B2(G169), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n379), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n379), .B1(new_n403), .B2(G200), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n399), .A2(G190), .A3(new_n400), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT73), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(G200), .B1(new_n391), .B2(new_n392), .ZN(new_n409));
  INV_X1    g0209(.A(new_n379), .ZN(new_n410));
  AND4_X1   g0210(.A1(KEYINPUT73), .A2(new_n409), .A3(new_n407), .A4(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n405), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G169), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G238), .A2(G1698), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n286), .B(new_n415), .C1(new_n238), .C2(G1698), .ZN(new_n416));
  INV_X1    g0216(.A(G107), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n331), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(new_n285), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n342), .B1(new_n223), .B2(new_n280), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n414), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n421), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n423), .A2(new_n419), .A3(new_n300), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n305), .A2(new_n253), .B1(G20), .B2(G77), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n425), .A2(KEYINPUT68), .ZN(new_n426));
  XNOR2_X1  g0226(.A(KEYINPUT15), .B(G87), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n425), .A2(KEYINPUT68), .B1(new_n260), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n310), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n373), .B1(new_n207), .B2(G20), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n268), .A2(new_n431), .B1(new_n373), .B2(new_n266), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n422), .B(new_n424), .C1(new_n430), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n426), .A2(new_n429), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n264), .ZN(new_n436));
  OAI21_X1  g0236(.A(G200), .B1(new_n420), .B2(new_n421), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n423), .A2(new_n419), .A3(G190), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n436), .A2(new_n437), .A3(new_n432), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  XOR2_X1   g0240(.A(new_n440), .B(KEYINPUT69), .Z(new_n441));
  NAND4_X1  g0241(.A1(new_n304), .A2(new_n368), .A3(new_n413), .A4(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  XNOR2_X1  g0243(.A(KEYINPUT81), .B(KEYINPUT21), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT80), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n207), .A2(G33), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n310), .A2(G116), .A3(new_n265), .A4(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G116), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n266), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(G20), .B1(G33), .B2(G283), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n259), .A2(G97), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n449), .A2(G20), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT20), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n310), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n451), .A2(new_n452), .B1(G20), .B2(new_n449), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT20), .B1(new_n264), .B2(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n448), .B(new_n450), .C1(new_n457), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G169), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT5), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n207), .B(G45), .C1(new_n462), .C2(G41), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n273), .A2(KEYINPUT5), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G274), .ZN(new_n466));
  INV_X1    g0266(.A(new_n214), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n466), .B1(new_n467), .B2(new_n276), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(G270), .B(new_n277), .C1(new_n463), .C2(new_n464), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G264), .A2(G1698), .ZN(new_n472));
  INV_X1    g0272(.A(G257), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(G1698), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n474), .A2(new_n318), .A3(new_n319), .A4(new_n320), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n331), .A2(G303), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n285), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT79), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT79), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n477), .A2(new_n480), .A3(new_n285), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n471), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n446), .B1(new_n461), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n471), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n480), .B1(new_n477), .B2(new_n285), .ZN(new_n485));
  AOI211_X1 g0285(.A(KEYINPUT79), .B(new_n284), .C1(new_n475), .C2(new_n476), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n487), .A2(KEYINPUT80), .A3(G169), .A4(new_n460), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n445), .B1(new_n483), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n460), .B1(new_n487), .B2(G200), .ZN(new_n490));
  OAI211_X1 g0290(.A(G190), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n456), .B1(new_n310), .B2(new_n455), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n264), .A2(KEYINPUT20), .A3(new_n458), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n493), .A2(new_n494), .B1(new_n449), .B2(new_n266), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n414), .B1(new_n495), .B2(new_n448), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(KEYINPUT21), .A3(new_n487), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n482), .A2(G179), .A3(new_n460), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n489), .A2(new_n492), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n265), .A2(G97), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n310), .A2(new_n265), .A3(new_n447), .ZN(new_n503));
  INV_X1    g0303(.A(G97), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT75), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n254), .A2(new_n373), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  XNOR2_X1  g0308(.A(G97), .B(G107), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT6), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(new_n504), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n509), .A2(new_n510), .B1(new_n417), .B2(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n506), .B(new_n508), .C1(new_n512), .C2(new_n208), .ZN(new_n513));
  AND2_X1   g0313(.A1(G97), .A2(G107), .ZN(new_n514));
  NOR2_X1   g0314(.A1(G97), .A2(G107), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n510), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n417), .A2(KEYINPUT6), .A3(G97), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n208), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(KEYINPUT75), .B1(new_n518), .B2(new_n507), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT7), .B1(new_n331), .B2(new_n208), .ZN(new_n520));
  AOI211_X1 g0320(.A(new_n324), .B(G20), .C1(new_n319), .C2(new_n330), .ZN(new_n521));
  OAI21_X1  g0321(.A(G107), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n513), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n505), .B1(new_n523), .B2(new_n264), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n319), .A2(new_n330), .A3(G250), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n287), .B1(new_n525), .B2(KEYINPUT4), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n287), .A2(KEYINPUT4), .A3(G244), .ZN(new_n527));
  INV_X1    g0327(.A(G283), .ZN(new_n528));
  OAI22_X1  g0328(.A1(new_n331), .A2(new_n527), .B1(new_n259), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n318), .A2(new_n320), .A3(G244), .A4(new_n319), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT4), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n284), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(G257), .B(new_n277), .C1(new_n463), .C2(new_n464), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n469), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(G200), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n527), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n286), .A2(new_n538), .B1(G33), .B2(G283), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n532), .B1(new_n286), .B2(G250), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n533), .B(new_n539), .C1(new_n287), .C2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n536), .B1(new_n541), .B2(new_n285), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G190), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n524), .A2(new_n537), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n541), .A2(new_n285), .ZN(new_n545));
  INV_X1    g0345(.A(new_n536), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n414), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI211_X1 g0347(.A(new_n300), .B(new_n536), .C1(new_n541), .C2(new_n285), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n544), .B1(new_n549), .B2(new_n524), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT84), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n320), .A2(new_n319), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n552), .A2(new_n208), .A3(G87), .A4(new_n318), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT83), .ZN(new_n554));
  INV_X1    g0354(.A(G87), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(G20), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n556), .A2(new_n319), .A3(new_n330), .ZN(new_n557));
  XNOR2_X1  g0357(.A(KEYINPUT82), .B(KEYINPUT22), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT22), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT82), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT82), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT22), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n564), .A2(new_n286), .A3(KEYINPUT83), .A4(new_n556), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n553), .A2(KEYINPUT22), .B1(new_n559), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT23), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n208), .B2(G107), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n417), .A2(KEYINPUT23), .A3(G20), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n568), .A2(new_n569), .B1(new_n260), .B2(G116), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT24), .B1(new_n566), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n559), .A2(new_n565), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n318), .A2(new_n320), .A3(new_n208), .A4(new_n319), .ZN(new_n574));
  OAI21_X1  g0374(.A(KEYINPUT22), .B1(new_n574), .B2(new_n555), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT24), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(new_n577), .A3(new_n570), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n310), .B1(new_n572), .B2(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n207), .A2(new_n417), .A3(G13), .A4(G20), .ZN(new_n580));
  XNOR2_X1  g0380(.A(new_n580), .B(KEYINPUT25), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n310), .A2(new_n265), .A3(new_n447), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n581), .B1(new_n582), .B2(G107), .ZN(new_n583));
  NAND2_X1  g0383(.A1(G257), .A2(G1698), .ZN(new_n584));
  INV_X1    g0384(.A(G250), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n584), .B1(new_n585), .B2(G1698), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n586), .A2(new_n318), .A3(new_n319), .A4(new_n320), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G33), .A2(G294), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n285), .ZN(new_n590));
  OAI211_X1 g0390(.A(G264), .B(new_n277), .C1(new_n463), .C2(new_n464), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n590), .A2(G190), .A3(new_n469), .A4(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n284), .B1(new_n587), .B2(new_n588), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n465), .A2(new_n468), .ZN(new_n594));
  INV_X1    g0394(.A(new_n591), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n583), .B(new_n592), .C1(new_n596), .C2(new_n293), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n551), .B1(new_n579), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n597), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n577), .B1(new_n576), .B2(new_n570), .ZN(new_n600));
  AOI211_X1 g0400(.A(KEYINPUT24), .B(new_n571), .C1(new_n573), .C2(new_n575), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n264), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n602), .A3(KEYINPUT84), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n550), .B1(new_n598), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n582), .A2(new_n428), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT77), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT19), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n381), .B2(new_n208), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n555), .A2(new_n504), .A3(new_n417), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n208), .A2(G33), .A3(G97), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n608), .A2(new_n609), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n203), .B2(new_n574), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n264), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n428), .A2(new_n265), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n606), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  AOI211_X1 g0416(.A(KEYINPUT77), .B(new_n614), .C1(new_n612), .C2(new_n264), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n605), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT76), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n585), .B1(new_n274), .B2(G1), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n207), .A2(new_n466), .A3(G45), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n277), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  OR2_X1    g0423(.A1(G238), .A2(G1698), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(G244), .B2(new_n287), .ZN(new_n625));
  OAI22_X1  g0425(.A1(new_n321), .A2(new_n625), .B1(new_n259), .B2(new_n449), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n623), .B1(new_n626), .B2(new_n285), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n627), .A2(new_n414), .ZN(new_n628));
  AOI211_X1 g0428(.A(new_n300), .B(new_n623), .C1(new_n626), .C2(new_n285), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n619), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(G179), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n631), .B(KEYINPUT76), .C1(new_n414), .C2(new_n627), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n618), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT78), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n626), .A2(new_n285), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n293), .B1(new_n635), .B2(new_n622), .ZN(new_n636));
  AOI211_X1 g0436(.A(new_n362), .B(new_n623), .C1(new_n626), .C2(new_n285), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n552), .A2(new_n208), .A3(G68), .A4(new_n318), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n310), .B1(new_n639), .B2(new_n611), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT77), .B1(new_n640), .B2(new_n614), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n613), .A2(new_n606), .A3(new_n615), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n503), .A2(new_n555), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n627), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT78), .B1(new_n646), .B2(new_n362), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n638), .A2(new_n643), .A3(new_n645), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n633), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n596), .A2(new_n300), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(G169), .B2(new_n596), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n602), .B2(new_n583), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  AND4_X1   g0453(.A1(new_n443), .A2(new_n500), .A3(new_n604), .A4(new_n653), .ZN(G372));
  NAND2_X1  g0454(.A1(new_n598), .A2(new_n603), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n524), .A2(new_n537), .A3(new_n543), .ZN(new_n656));
  OAI21_X1  g0456(.A(G169), .B1(new_n534), .B2(new_n536), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n542), .A2(G179), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n523), .A2(new_n264), .ZN(new_n659));
  INV_X1    g0459(.A(new_n505), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n657), .A2(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n628), .A2(new_n629), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n643), .B2(new_n605), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n645), .B1(new_n616), .B2(new_n617), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT85), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n636), .A2(new_n637), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n643), .A2(KEYINPUT85), .A3(new_n645), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n655), .A2(new_n662), .A3(new_n665), .A4(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT86), .ZN(new_n673));
  AOI21_X1  g0473(.A(KEYINPUT85), .B1(new_n643), .B2(new_n645), .ZN(new_n674));
  AOI211_X1 g0474(.A(new_n667), .B(new_n644), .C1(new_n641), .C2(new_n642), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n664), .B1(new_n676), .B2(new_n669), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT86), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n604), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n488), .ZN(new_n680));
  AOI21_X1  g0480(.A(KEYINPUT80), .B1(new_n496), .B2(new_n487), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n444), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n499), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT87), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT87), .B1(new_n489), .B2(new_n499), .ZN(new_n686));
  INV_X1    g0486(.A(new_n652), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n673), .A2(new_n679), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(KEYINPUT88), .B1(new_n547), .B2(new_n548), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT88), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n657), .A2(new_n658), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n524), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(new_n671), .A3(new_n665), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(KEYINPUT26), .ZN(new_n695));
  INV_X1    g0495(.A(new_n661), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT26), .B1(new_n649), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n665), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n689), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n443), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n360), .A2(new_n352), .ZN(new_n702));
  INV_X1    g0502(.A(new_n434), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n408), .B2(new_n411), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n704), .A2(new_n405), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n365), .A2(new_n366), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n702), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n296), .B(new_n297), .Z(new_n708));
  AOI21_X1  g0508(.A(new_n303), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n701), .A2(new_n709), .ZN(G369));
  NAND2_X1  g0510(.A1(new_n685), .A2(new_n686), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n712), .A2(KEYINPUT27), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(KEYINPUT27), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(G213), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(G343), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n718), .B1(new_n495), .B2(new_n448), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n711), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g0520(.A(new_n500), .B(KEYINPUT89), .Z(new_n721));
  OAI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n719), .ZN(new_n722));
  INV_X1    g0522(.A(new_n583), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n717), .B1(new_n579), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n652), .B1(new_n655), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n652), .B2(new_n718), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n722), .A2(G330), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n652), .A2(new_n718), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n717), .B1(new_n682), .B2(new_n683), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(G399));
  NAND2_X1  g0531(.A1(new_n211), .A2(new_n273), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n609), .A2(G116), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n732), .A2(G1), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(new_n220), .B2(new_n732), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT28), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n694), .A2(KEYINPUT26), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT26), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n633), .A2(new_n648), .A3(new_n661), .A4(new_n738), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n739), .A2(new_n665), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n489), .A2(new_n652), .A3(new_n499), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n737), .B(new_n740), .C1(new_n672), .C2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT91), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n718), .A2(KEYINPUT29), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n743), .B1(new_n742), .B2(new_n744), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n717), .B1(new_n689), .B2(new_n699), .ZN(new_n747));
  XNOR2_X1  g0547(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n745), .A2(new_n746), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G330), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n604), .A2(new_n500), .A3(new_n653), .A4(new_n718), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT30), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n593), .A2(new_n595), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n542), .A2(new_n755), .A3(new_n629), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n754), .B1(new_n756), .B2(new_n487), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n755), .A2(new_n627), .A3(G179), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n758), .A2(new_n482), .A3(KEYINPUT30), .A4(new_n542), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n596), .A2(G179), .A3(new_n627), .ZN(new_n760));
  INV_X1    g0560(.A(new_n542), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n760), .A2(new_n487), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n757), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  AND3_X1   g0563(.A1(new_n763), .A2(KEYINPUT31), .A3(new_n717), .ZN(new_n764));
  AOI21_X1  g0564(.A(KEYINPUT31), .B1(new_n763), .B2(new_n717), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n752), .B1(new_n753), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n751), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n736), .B1(new_n768), .B2(G1), .ZN(G364));
  INV_X1    g0569(.A(G13), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G45), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n732), .A2(G1), .A3(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n211), .A2(new_n286), .ZN(new_n775));
  INV_X1    g0575(.A(G355), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n775), .A2(new_n776), .B1(G116), .B2(new_n211), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n246), .A2(G45), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n211), .A2(new_n321), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n274), .B2(new_n221), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n777), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n218), .B1(G20), .B2(new_n414), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G13), .A2(G33), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n774), .B1(new_n781), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G179), .A2(G200), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n208), .B1(new_n789), .B2(G190), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n504), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n208), .A2(new_n300), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(G190), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT95), .B(G159), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n789), .A2(G20), .A3(new_n362), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n795), .A2(new_n203), .B1(KEYINPUT32), .B2(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n791), .B(new_n799), .C1(KEYINPUT32), .C2(new_n798), .ZN(new_n800));
  NOR4_X1   g0600(.A1(new_n208), .A2(new_n293), .A3(G179), .A4(G190), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT96), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G107), .ZN(new_n803));
  NOR4_X1   g0603(.A1(new_n208), .A2(new_n362), .A3(new_n293), .A4(G179), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n286), .B1(new_n805), .B2(new_n555), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n793), .A2(new_n362), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(G50), .B2(new_n807), .ZN(new_n808));
  AND3_X1   g0608(.A1(new_n800), .A2(new_n803), .A3(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n792), .B(KEYINPUT92), .Z(new_n810));
  NAND3_X1  g0610(.A1(new_n810), .A2(G190), .A3(new_n293), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT93), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n810), .A2(new_n362), .A3(new_n293), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n816), .A2(KEYINPUT94), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(KEYINPUT94), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n809), .B1(new_n202), .B2(new_n815), .C1(new_n373), .C2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n790), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n807), .A2(G326), .B1(G294), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(G311), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n819), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT97), .ZN(new_n825));
  INV_X1    g0625(.A(G303), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n331), .B1(new_n805), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n797), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n827), .B1(G329), .B2(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(KEYINPUT33), .B(G317), .Z(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n795), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(G283), .B2(new_n802), .ZN(new_n832));
  INV_X1    g0632(.A(G322), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(new_n815), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n820), .B1(new_n825), .B2(new_n834), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n835), .A2(KEYINPUT98), .ZN(new_n836));
  INV_X1    g0636(.A(new_n782), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n835), .B2(KEYINPUT98), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n788), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n785), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n722), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n722), .A2(G330), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n773), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n722), .A2(G330), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n841), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT99), .Z(G396));
  NOR2_X1   g0646(.A1(new_n782), .A2(new_n783), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n807), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n849), .A2(new_n826), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n791), .B(new_n850), .C1(G283), .C2(new_n794), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n331), .B1(new_n797), .B2(new_n823), .C1(new_n805), .C2(new_n417), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(G87), .B2(new_n802), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(G294), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n854), .B1(new_n449), .B2(new_n819), .C1(new_n855), .C2(new_n815), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n794), .A2(G150), .B1(new_n807), .B2(G137), .ZN(new_n858));
  INV_X1    g0658(.A(G143), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n858), .B1(new_n819), .B2(new_n796), .C1(new_n859), .C2(new_n815), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT34), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n790), .A2(new_n202), .ZN(new_n862));
  INV_X1    g0662(.A(new_n321), .ZN(new_n863));
  INV_X1    g0663(.A(G132), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n863), .B1(new_n864), .B2(new_n797), .C1(new_n805), .C2(new_n201), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n862), .B(new_n865), .C1(G68), .C2(new_n802), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n857), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n774), .B1(G77), .B2(new_n848), .C1(new_n867), .C2(new_n837), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n868), .A2(KEYINPUT100), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(KEYINPUT100), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n717), .B1(new_n430), .B2(new_n433), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n434), .A2(new_n439), .A3(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT101), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n434), .A2(new_n439), .A3(KEYINPUT101), .A4(new_n871), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n703), .A2(new_n717), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n869), .B(new_n870), .C1(new_n784), .C2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n747), .A2(new_n877), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n879), .A2(KEYINPUT102), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(KEYINPUT102), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n717), .B1(new_n874), .B2(new_n875), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n689), .B2(new_n699), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n880), .A2(new_n881), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n767), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n773), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n886), .A2(new_n887), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n878), .B1(new_n889), .B2(new_n890), .ZN(G384));
  NOR2_X1   g0691(.A1(new_n771), .A2(new_n207), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n753), .A2(new_n766), .ZN(new_n893));
  INV_X1    g0693(.A(new_n877), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n379), .A2(new_n717), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n412), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n405), .B(new_n895), .C1(new_n408), .C2(new_n411), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n893), .A2(new_n899), .A3(KEYINPUT40), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n715), .B1(new_n357), .B2(new_n308), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n357), .A2(new_n308), .ZN(new_n902));
  INV_X1    g0702(.A(new_n351), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n715), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n357), .A2(new_n308), .A3(new_n364), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT37), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n904), .A2(new_n906), .A3(new_n910), .A4(new_n907), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n367), .A2(new_n901), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT106), .B1(new_n912), .B2(KEYINPUT38), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n367), .A2(new_n901), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n357), .A2(new_n308), .A3(new_n364), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n915), .A2(new_n358), .A3(new_n901), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n911), .B1(new_n916), .B2(new_n910), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT106), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT38), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n913), .A2(new_n921), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n345), .A2(new_n350), .A3(new_n715), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n321), .A2(new_n324), .A3(new_n208), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n324), .B1(new_n321), .B2(new_n208), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n924), .A2(new_n925), .A3(new_n203), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n328), .B1(new_n926), .B2(new_n315), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(new_n264), .A3(new_n356), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n923), .B1(new_n928), .B2(new_n308), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT37), .B1(new_n929), .B2(new_n915), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n911), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT104), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n911), .A2(new_n930), .A3(KEYINPUT104), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n715), .B1(new_n928), .B2(new_n308), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n920), .B1(new_n367), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n900), .B1(new_n922), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n367), .A2(new_n936), .ZN(new_n940));
  AND3_X1   g0740(.A1(new_n911), .A2(new_n930), .A3(KEYINPUT104), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT104), .B1(new_n911), .B2(new_n930), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n920), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT105), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n937), .B(new_n945), .C1(new_n942), .C2(new_n941), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n945), .B1(new_n935), .B2(new_n937), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n893), .A2(new_n899), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT40), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n939), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AND3_X1   g0754(.A1(new_n954), .A2(new_n443), .A3(new_n893), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n954), .B1(new_n443), .B2(new_n893), .ZN(new_n956));
  OR3_X1    g0756(.A1(new_n955), .A2(new_n956), .A3(new_n752), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n702), .A2(new_n905), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n897), .A2(new_n898), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n434), .A2(new_n717), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n959), .B1(new_n884), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n958), .B1(new_n962), .B2(new_n949), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n919), .B1(new_n918), .B2(new_n920), .ZN(new_n964));
  AOI211_X1 g0764(.A(KEYINPUT106), .B(KEYINPUT38), .C1(new_n914), .C2(new_n917), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n938), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT39), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n405), .ZN(new_n969));
  OAI211_X1 g0769(.A(KEYINPUT39), .B(new_n944), .C1(new_n947), .C2(new_n948), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n968), .A2(new_n969), .A3(new_n718), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n963), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n709), .B1(new_n750), .B2(new_n442), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n972), .B(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n892), .B1(new_n957), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n974), .B2(new_n957), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n311), .A2(new_n220), .A3(new_n373), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n203), .A2(G50), .ZN(new_n978));
  OAI211_X1 g0778(.A(G1), .B(new_n770), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n512), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n980), .A2(KEYINPUT35), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(KEYINPUT35), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n981), .A2(new_n982), .A3(G116), .A4(new_n219), .ZN(new_n983));
  XNOR2_X1  g0783(.A(KEYINPUT103), .B(KEYINPUT36), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n983), .B(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n976), .A2(new_n979), .A3(new_n985), .ZN(G367));
  OAI21_X1  g0786(.A(new_n662), .B1(new_n524), .B2(new_n718), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n693), .A2(new_n717), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n726), .A2(new_n729), .A3(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n989), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n696), .B1(new_n991), .B2(new_n687), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n990), .A2(KEYINPUT42), .B1(new_n992), .B2(new_n718), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(KEYINPUT42), .B2(new_n990), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n676), .A2(new_n718), .ZN(new_n995));
  MUX2_X1   g0795(.A(new_n677), .B(new_n664), .S(new_n995), .Z(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(KEYINPUT43), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n996), .A2(KEYINPUT43), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n998), .B(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n727), .A2(new_n991), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n772), .A2(G1), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n730), .A2(new_n728), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(KEYINPUT44), .B1(new_n1006), .B2(new_n989), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT44), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1005), .A2(new_n1008), .A3(new_n991), .ZN(new_n1009));
  XOR2_X1   g0809(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n1010));
  NAND4_X1  g0810(.A1(new_n730), .A2(new_n728), .A3(new_n989), .A4(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1010), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n1005), .B2(new_n991), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1007), .A2(new_n1009), .A3(new_n1011), .A4(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n727), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1013), .A2(new_n1011), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1017), .A2(new_n727), .A3(new_n1007), .A4(new_n1009), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT108), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n730), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n726), .A2(KEYINPUT108), .A3(new_n729), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(new_n726), .C2(new_n729), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(new_n842), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n768), .B1(new_n1019), .B2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n732), .B(KEYINPUT41), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT109), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1004), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1025), .A2(KEYINPUT109), .A3(new_n1027), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1003), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n996), .A2(new_n840), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n242), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n786), .B1(new_n211), .B2(new_n427), .C1(new_n1034), .C2(new_n779), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n774), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n805), .A2(new_n449), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(KEYINPUT46), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n417), .B2(new_n790), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n1037), .A2(KEYINPUT46), .B1(new_n855), .B2(new_n795), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n849), .A2(new_n823), .ZN(new_n1041));
  INV_X1    g0841(.A(G317), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n801), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n321), .B1(new_n797), .B2(new_n1042), .C1(new_n1043), .C2(new_n504), .ZN(new_n1044));
  NOR4_X1   g0844(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .A4(new_n1044), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n819), .B2(new_n528), .C1(new_n826), .C2(new_n815), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n821), .A2(G68), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n849), .B2(new_n859), .C1(new_n795), .C2(new_n796), .ZN(new_n1048));
  INV_X1    g0848(.A(G137), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n286), .B1(new_n797), .B2(new_n1049), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n805), .A2(new_n202), .B1(new_n1043), .B2(new_n373), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n1048), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n819), .B2(new_n201), .C1(new_n252), .C2(new_n815), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1046), .A2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT47), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1036), .B1(new_n1055), .B2(new_n782), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1033), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1032), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(G387));
  NOR2_X1   g0860(.A1(new_n726), .A2(new_n840), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n775), .A2(new_n733), .B1(G107), .B2(new_n211), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n239), .A2(G45), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n733), .ZN(new_n1064));
  AOI211_X1 g0864(.A(G45), .B(new_n1064), .C1(G68), .C2(G77), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n305), .A2(new_n201), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT50), .Z(new_n1067));
  AOI21_X1  g0867(.A(new_n779), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1062), .B1(new_n1063), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n774), .B1(new_n1069), .B2(new_n787), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n863), .B1(new_n252), .B2(new_n797), .C1(new_n805), .C2(new_n373), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n821), .A2(new_n428), .ZN(new_n1072));
  INV_X1    g0872(.A(G159), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1072), .B1(new_n849), .B2(new_n1073), .C1(new_n258), .C2(new_n795), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1071), .B(new_n1074), .C1(G97), .C2(new_n802), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n201), .B2(new_n815), .C1(new_n203), .C2(new_n819), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n804), .A2(G294), .B1(new_n821), .B2(G283), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n794), .A2(G311), .B1(new_n807), .B2(G322), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1078), .B1(new_n819), .B2(new_n826), .C1(new_n1042), .C2(new_n815), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT48), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1077), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT110), .Z(new_n1082));
  NAND2_X1  g0882(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1082), .A2(KEYINPUT49), .A3(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G326), .A2(new_n828), .B1(new_n801), .B2(G116), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1084), .A2(new_n321), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT49), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1076), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1061), .B(new_n1070), .C1(new_n1088), .C2(new_n782), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1024), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1089), .B1(new_n1090), .B2(new_n1004), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1024), .A2(new_n767), .A3(new_n751), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n1092), .A2(new_n732), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1090), .A2(new_n768), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(G393));
  INV_X1    g0895(.A(new_n1019), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n732), .B1(new_n1096), .B2(new_n1092), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1004), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n786), .B1(new_n504), .B2(new_n211), .C1(new_n249), .C2(new_n779), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n1100), .A2(new_n774), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n815), .A2(new_n823), .B1(new_n1042), .B2(new_n849), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT52), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n795), .A2(new_n826), .B1(new_n790), .B2(new_n449), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n331), .B1(new_n797), .B2(new_n833), .C1(new_n805), .C2(new_n528), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1104), .B(new_n1105), .C1(G107), .C2(new_n802), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1103), .B(new_n1106), .C1(new_n855), .C2(new_n819), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n815), .A2(new_n1073), .B1(new_n252), .B2(new_n849), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT51), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n790), .A2(new_n373), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n794), .B2(G50), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n804), .A2(G68), .B1(new_n828), .B2(G143), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1111), .A2(new_n863), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(G87), .B2(new_n802), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1109), .B(new_n1114), .C1(new_n258), .C2(new_n819), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n1107), .A2(new_n1115), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1101), .B1(new_n840), .B2(new_n989), .C1(new_n1116), .C2(new_n837), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1098), .A2(new_n1099), .A3(new_n1117), .ZN(G390));
  NAND2_X1  g0918(.A1(new_n443), .A2(new_n767), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n709), .B(new_n1119), .C1(new_n750), .C2(new_n442), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT112), .ZN(new_n1121));
  AND4_X1   g0921(.A1(new_n1121), .A2(new_n893), .A3(new_n899), .A4(G330), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1121), .B1(new_n767), .B2(new_n899), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n960), .B1(new_n742), .B2(new_n882), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n752), .B(new_n894), .C1(new_n753), .C2(new_n766), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1125), .B1(new_n1126), .B2(new_n959), .ZN(new_n1127));
  OAI21_X1  g0927(.A(KEYINPUT113), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n893), .A2(new_n899), .A3(G330), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(KEYINPUT112), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n767), .A2(new_n1121), .A3(new_n899), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n959), .B1(new_n767), .B2(new_n877), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n740), .B1(new_n672), .B2(new_n741), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n737), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n882), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n960), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT113), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1132), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1128), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1129), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1143), .A2(new_n1133), .B1(new_n884), .B2(new_n960), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1120), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT115), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n969), .A2(new_n718), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n968), .A2(new_n970), .B1(new_n1147), .B2(new_n961), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n913), .A2(new_n921), .B1(new_n935), .B2(new_n937), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n959), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1125), .A2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1147), .B(KEYINPUT111), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1149), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1143), .B1(new_n1148), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n961), .A2(new_n1147), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n941), .A2(new_n942), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n940), .A2(KEYINPUT38), .ZN(new_n1157));
  OAI21_X1  g0957(.A(KEYINPUT105), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AOI221_X4 g0958(.A(new_n967), .B1(new_n920), .B2(new_n943), .C1(new_n1158), .C2(new_n946), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT39), .B1(new_n922), .B2(new_n938), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1155), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  OR3_X1    g0961(.A1(new_n1149), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1161), .A2(new_n1132), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1154), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1146), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n732), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT114), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n1124), .A2(KEYINPUT113), .A3(new_n1127), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1140), .B1(new_n1132), .B2(new_n1139), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1144), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1120), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1167), .B1(new_n1164), .B2(new_n1172), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1145), .A2(KEYINPUT114), .A3(new_n1163), .A4(new_n1154), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1165), .A2(new_n1166), .A3(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1154), .A2(new_n1163), .A3(new_n1004), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n783), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n331), .B1(new_n797), .B2(new_n855), .C1(new_n805), .C2(new_n555), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1110), .B1(new_n794), .B2(G107), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n528), .B2(new_n849), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1179), .B(new_n1181), .C1(G68), .C2(new_n802), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1182), .B1(new_n819), .B2(new_n504), .C1(new_n449), .C2(new_n815), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n804), .A2(G150), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1184), .B(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(G128), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n795), .A2(new_n1049), .B1(new_n849), .B2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n790), .A2(new_n1073), .ZN(new_n1189));
  INV_X1    g0989(.A(G125), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n286), .B1(new_n797), .B2(new_n1190), .C1(new_n1043), .C2(new_n201), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(new_n1186), .A2(new_n1188), .A3(new_n1189), .A4(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT54), .B(G143), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1192), .B1(new_n819), .B2(new_n1193), .C1(new_n864), .C2(new_n815), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n837), .B1(new_n1183), .B2(new_n1194), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n773), .B(new_n1195), .C1(new_n258), .C2(new_n847), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1178), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1176), .A2(new_n1177), .A3(new_n1197), .ZN(G378));
  INV_X1    g0998(.A(KEYINPUT57), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1120), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n708), .A2(new_n302), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n271), .A2(new_n905), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT55), .Z(new_n1205));
  NOR2_X1   g1005(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1205), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n304), .A2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1202), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n304), .A2(new_n1207), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1210), .A2(new_n1201), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1209), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n954), .B2(G330), .ZN(new_n1215));
  AOI21_X1  g1015(.A(KEYINPUT40), .B1(new_n949), .B2(new_n951), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1216), .A2(new_n939), .A3(new_n1213), .A4(new_n752), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n972), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n963), .A2(new_n971), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n954), .A2(G330), .A3(new_n1214), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n966), .A2(KEYINPUT40), .A3(new_n951), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1158), .A2(new_n946), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n950), .B1(new_n1222), .B2(new_n944), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1221), .B(G330), .C1(new_n1223), .C2(KEYINPUT40), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n1213), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1219), .A2(new_n1220), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1218), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1199), .B1(new_n1200), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT121), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT121), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1231), .B(new_n1199), .C1(new_n1200), .C2(new_n1228), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1218), .A2(KEYINPUT120), .A3(new_n1226), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT120), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1219), .A2(new_n1220), .A3(new_n1234), .A4(new_n1225), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1233), .A2(KEYINPUT57), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1175), .A2(new_n1171), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n732), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1230), .A2(new_n1232), .A3(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n774), .B1(new_n848), .B2(G50), .ZN(new_n1240));
  AOI211_X1 g1040(.A(G33), .B(G41), .C1(new_n828), .C2(G124), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1043), .B2(new_n796), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n795), .A2(new_n864), .B1(new_n805), .B2(new_n1193), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n815), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1243), .B1(new_n1244), .B2(G128), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n807), .A2(G125), .B1(G150), .B2(new_n821), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT117), .Z(new_n1247));
  OAI211_X1 g1047(.A(new_n1245), .B(new_n1247), .C1(new_n1049), .C2(new_n819), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1242), .B1(new_n1248), .B2(KEYINPUT59), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(KEYINPUT59), .B2(new_n1248), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1043), .A2(new_n202), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(G77), .B2(new_n804), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n528), .B2(new_n797), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1047), .B1(new_n849), .B2(new_n449), .C1(new_n504), .C2(new_n795), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n321), .A2(new_n273), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n1256), .B1(new_n819), .B2(new_n427), .C1(new_n417), .C2(new_n815), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT58), .ZN(new_n1258));
  AOI21_X1  g1058(.A(G50), .B1(new_n259), .B2(new_n273), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1257), .A2(new_n1258), .B1(new_n1255), .B2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1250), .B(new_n1260), .C1(new_n1258), .C2(new_n1257), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1240), .B1(new_n1261), .B2(new_n782), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n1214), .B2(new_n784), .ZN(new_n1263));
  XOR2_X1   g1063(.A(new_n1263), .B(KEYINPUT119), .Z(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n1227), .B2(new_n1004), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1239), .A2(new_n1265), .ZN(G375));
  NAND3_X1  g1066(.A1(new_n1142), .A2(new_n1120), .A3(new_n1144), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1146), .A2(new_n1027), .A3(new_n1267), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n795), .A2(new_n1193), .B1(new_n201), .B2(new_n790), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n321), .B(new_n1269), .C1(G132), .C2(new_n807), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n797), .A2(new_n1187), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n1271), .B(new_n1251), .C1(G159), .C2(new_n804), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1273));
  OAI221_X1 g1073(.A(new_n1273), .B1(new_n1049), .B2(new_n815), .C1(new_n252), .C2(new_n819), .ZN(new_n1274));
  OAI221_X1 g1074(.A(new_n331), .B1(new_n797), .B2(new_n826), .C1(new_n805), .C2(new_n504), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n1072), .B1(new_n849), .B2(new_n855), .C1(new_n449), .C2(new_n795), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n1275), .B(new_n1276), .C1(G77), .C2(new_n802), .ZN(new_n1277));
  OAI221_X1 g1077(.A(new_n1277), .B1(new_n417), .B2(new_n819), .C1(new_n528), .C2(new_n815), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n837), .B1(new_n1274), .B2(new_n1278), .ZN(new_n1279));
  AOI211_X1 g1079(.A(new_n773), .B(new_n1279), .C1(new_n203), .C2(new_n847), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1280), .B(KEYINPUT122), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(new_n783), .B2(new_n1150), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(new_n1170), .B2(new_n1004), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1268), .A2(new_n1283), .ZN(G381));
  NOR4_X1   g1084(.A1(G390), .A2(G396), .A3(G393), .A4(G384), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1285), .A2(new_n1059), .A3(new_n1283), .A4(new_n1268), .ZN(new_n1286));
  OR3_X1    g1086(.A1(new_n1286), .A2(G375), .A3(G378), .ZN(G407));
  INV_X1    g1087(.A(G378), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n716), .A2(G213), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(G407), .B(G213), .C1(G375), .C2(new_n1291), .ZN(G409));
  INV_X1    g1092(.A(KEYINPUT60), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1267), .A2(new_n1293), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1142), .A2(KEYINPUT60), .A3(new_n1120), .A4(new_n1144), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1294), .A2(new_n1166), .A3(new_n1172), .A4(new_n1295), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1296), .A2(G384), .A3(new_n1283), .ZN(new_n1297));
  AOI21_X1  g1097(.A(G384), .B1(new_n1296), .B2(new_n1283), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT125), .B1(new_n1299), .B2(KEYINPUT124), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT124), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT125), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1301), .B(new_n1302), .C1(new_n1297), .C2(new_n1298), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1300), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1290), .A2(G2897), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1305), .B1(new_n1299), .B2(KEYINPUT124), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1305), .ZN(new_n1308));
  OR2_X1    g1108(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1308), .B1(new_n1309), .B2(new_n1301), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1310), .A2(new_n1300), .A3(new_n1303), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1307), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1239), .A2(G378), .A3(new_n1265), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1237), .A2(KEYINPUT123), .A3(new_n1027), .A4(new_n1227), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1233), .A2(new_n1004), .A3(new_n1235), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1315), .A2(new_n1263), .A3(new_n1316), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1200), .A2(new_n1228), .ZN(new_n1318));
  AOI21_X1  g1118(.A(KEYINPUT123), .B1(new_n1318), .B2(new_n1027), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1288), .B1(new_n1317), .B2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1314), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1289), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT61), .B1(new_n1313), .B2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1324), .B1(new_n1322), .B2(new_n1309), .ZN(new_n1325));
  INV_X1    g1125(.A(G390), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1326), .B1(new_n1032), .B2(new_n1058), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1031), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT109), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1329));
  NOR3_X1   g1129(.A1(new_n1328), .A2(new_n1329), .A3(new_n1004), .ZN(new_n1330));
  OAI211_X1 g1130(.A(G390), .B(new_n1057), .C1(new_n1330), .C2(new_n1003), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1327), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT126), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1333), .B1(new_n1059), .B2(G390), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(G393), .B(G396), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1332), .B1(new_n1334), .B2(new_n1336), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1327), .A2(new_n1331), .A3(new_n1333), .A4(new_n1335), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1290), .B1(new_n1314), .B2(new_n1320), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1340), .A2(KEYINPUT63), .A3(new_n1299), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1323), .A2(new_n1325), .A3(new_n1339), .A4(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT62), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1340), .A2(new_n1343), .A3(new_n1299), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT61), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1345), .B1(new_n1340), .B2(new_n1312), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1343), .B1(new_n1340), .B2(new_n1299), .ZN(new_n1347));
  NOR3_X1   g1147(.A1(new_n1344), .A2(new_n1346), .A3(new_n1347), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1342), .B1(new_n1348), .B2(new_n1339), .ZN(G405));
  NAND3_X1  g1149(.A1(G375), .A2(new_n1288), .A3(new_n1299), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1299), .B1(G375), .B2(new_n1288), .ZN(new_n1352));
  OAI211_X1 g1152(.A(new_n1338), .B(new_n1337), .C1(new_n1351), .C2(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1352), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1339), .A2(new_n1354), .A3(new_n1350), .ZN(new_n1355));
  AND2_X1   g1155(.A1(new_n1314), .A2(KEYINPUT127), .ZN(new_n1356));
  AND3_X1   g1156(.A1(new_n1353), .A2(new_n1355), .A3(new_n1356), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1356), .B1(new_n1353), .B2(new_n1355), .ZN(new_n1358));
  NOR2_X1   g1158(.A1(new_n1357), .A2(new_n1358), .ZN(G402));
endmodule


