

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582;

  XOR2_X1 U324 ( .A(n419), .B(n418), .Z(n560) );
  XNOR2_X1 U325 ( .A(n330), .B(n329), .ZN(n519) );
  XNOR2_X1 U326 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n292) );
  INV_X1 U327 ( .A(KEYINPUT95), .ZN(n312) );
  XNOR2_X1 U328 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n471) );
  XNOR2_X1 U329 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U330 ( .A(n472), .B(n471), .ZN(n526) );
  XNOR2_X1 U331 ( .A(n440), .B(n314), .ZN(n315) );
  NOR2_X1 U332 ( .A1(n420), .A2(n579), .ZN(n421) );
  NOR2_X1 U333 ( .A1(n530), .A2(n478), .ZN(n561) );
  XNOR2_X1 U334 ( .A(n479), .B(KEYINPUT121), .ZN(n480) );
  XNOR2_X1 U335 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U336 ( .A(n481), .B(n480), .ZN(G1348GAT) );
  XNOR2_X1 U337 ( .A(n458), .B(n457), .ZN(G1330GAT) );
  XOR2_X1 U338 ( .A(G155GAT), .B(G211GAT), .Z(n294) );
  XNOR2_X1 U339 ( .A(G127GAT), .B(G71GAT), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n308) );
  XOR2_X1 U341 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n296) );
  XNOR2_X1 U342 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n301) );
  XNOR2_X1 U344 ( .A(G8GAT), .B(G183GAT), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n297), .B(KEYINPUT76), .ZN(n323) );
  XOR2_X1 U346 ( .A(n323), .B(KEYINPUT12), .Z(n299) );
  NAND2_X1 U347 ( .A1(G231GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U348 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n306) );
  XOR2_X1 U350 ( .A(G57GAT), .B(KEYINPUT13), .Z(n439) );
  XOR2_X1 U351 ( .A(n439), .B(G78GAT), .Z(n304) );
  XNOR2_X1 U352 ( .A(G15GAT), .B(G1GAT), .ZN(n302) );
  XNOR2_X1 U353 ( .A(n302), .B(KEYINPUT68), .ZN(n423) );
  XNOR2_X1 U354 ( .A(G22GAT), .B(n423), .ZN(n303) );
  XNOR2_X1 U355 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U356 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U357 ( .A(n308), .B(n307), .Z(n574) );
  INV_X1 U358 ( .A(n574), .ZN(n482) );
  XOR2_X1 U359 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n310) );
  XNOR2_X1 U360 ( .A(KEYINPUT97), .B(KEYINPUT96), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n310), .B(n309), .ZN(n316) );
  XNOR2_X1 U362 ( .A(G176GAT), .B(G92GAT), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n311), .B(G64GAT), .ZN(n440) );
  NAND2_X1 U364 ( .A1(G226GAT), .A2(G233GAT), .ZN(n313) );
  XOR2_X1 U365 ( .A(n316), .B(n315), .Z(n322) );
  XOR2_X1 U366 ( .A(KEYINPUT21), .B(G204GAT), .Z(n318) );
  XNOR2_X1 U367 ( .A(G197GAT), .B(G211GAT), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n320) );
  XOR2_X1 U369 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n319) );
  XOR2_X1 U370 ( .A(n320), .B(n319), .Z(n370) );
  XNOR2_X1 U371 ( .A(n370), .B(G218GAT), .ZN(n321) );
  XOR2_X1 U372 ( .A(n322), .B(n321), .Z(n324) );
  XNOR2_X1 U373 ( .A(n324), .B(n323), .ZN(n330) );
  XOR2_X1 U374 ( .A(KEYINPUT79), .B(KEYINPUT17), .Z(n326) );
  XNOR2_X1 U375 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n325) );
  XNOR2_X1 U376 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U377 ( .A(G169GAT), .B(n327), .Z(n387) );
  XNOR2_X1 U378 ( .A(G36GAT), .B(G190GAT), .ZN(n328) );
  XNOR2_X1 U379 ( .A(n328), .B(KEYINPUT75), .ZN(n415) );
  XNOR2_X1 U380 ( .A(n387), .B(n415), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n519), .B(KEYINPUT27), .ZN(n391) );
  XOR2_X1 U382 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n332) );
  XNOR2_X1 U383 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U385 ( .A(KEYINPUT91), .B(KEYINPUT5), .Z(n334) );
  XNOR2_X1 U386 ( .A(G57GAT), .B(KEYINPUT92), .ZN(n333) );
  XNOR2_X1 U387 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U388 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U389 ( .A(G85GAT), .B(G148GAT), .Z(n338) );
  XNOR2_X1 U390 ( .A(G141GAT), .B(G120GAT), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U392 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U393 ( .A(n341), .B(KEYINPUT89), .Z(n345) );
  XOR2_X1 U394 ( .A(G155GAT), .B(KEYINPUT85), .Z(n343) );
  XNOR2_X1 U395 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n343), .B(n342), .ZN(n367) );
  XNOR2_X1 U397 ( .A(n367), .B(KEYINPUT90), .ZN(n344) );
  XNOR2_X1 U398 ( .A(n345), .B(n344), .ZN(n352) );
  XOR2_X1 U399 ( .A(G127GAT), .B(KEYINPUT0), .Z(n347) );
  XNOR2_X1 U400 ( .A(G113GAT), .B(G134GAT), .ZN(n346) );
  XNOR2_X1 U401 ( .A(n347), .B(n346), .ZN(n381) );
  XOR2_X1 U402 ( .A(G162GAT), .B(n381), .Z(n349) );
  NAND2_X1 U403 ( .A1(G225GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U404 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U405 ( .A(G29GAT), .B(n350), .Z(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n517) );
  NOR2_X1 U407 ( .A1(n391), .A2(n517), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n353), .B(KEYINPUT98), .ZN(n525) );
  XOR2_X1 U409 ( .A(KEYINPUT22), .B(KEYINPUT86), .Z(n355) );
  XNOR2_X1 U410 ( .A(KEYINPUT82), .B(KEYINPUT23), .ZN(n354) );
  XNOR2_X1 U411 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U412 ( .A(n356), .B(KEYINPUT24), .Z(n358) );
  XOR2_X1 U413 ( .A(G141GAT), .B(G22GAT), .Z(n422) );
  XNOR2_X1 U414 ( .A(n422), .B(KEYINPUT88), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n358), .B(n357), .ZN(n364) );
  XOR2_X1 U416 ( .A(G162GAT), .B(KEYINPUT71), .Z(n360) );
  XNOR2_X1 U417 ( .A(G50GAT), .B(G218GAT), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n360), .B(n359), .ZN(n410) );
  XOR2_X1 U419 ( .A(n410), .B(KEYINPUT87), .Z(n362) );
  NAND2_X1 U420 ( .A1(G228GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U421 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U422 ( .A(n364), .B(n363), .Z(n369) );
  XOR2_X1 U423 ( .A(G78GAT), .B(G148GAT), .Z(n366) );
  XNOR2_X1 U424 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n441) );
  XNOR2_X1 U426 ( .A(n441), .B(n367), .ZN(n368) );
  XNOR2_X1 U427 ( .A(n369), .B(n368), .ZN(n371) );
  XOR2_X1 U428 ( .A(n371), .B(n370), .Z(n476) );
  XOR2_X1 U429 ( .A(n476), .B(KEYINPUT28), .Z(n528) );
  NAND2_X1 U430 ( .A1(n525), .A2(n528), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n372), .B(KEYINPUT99), .ZN(n388) );
  XOR2_X1 U432 ( .A(KEYINPUT20), .B(G183GAT), .Z(n374) );
  XNOR2_X1 U433 ( .A(G15GAT), .B(G176GAT), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n374), .B(n373), .ZN(n385) );
  XOR2_X1 U435 ( .A(G120GAT), .B(G71GAT), .Z(n442) );
  XOR2_X1 U436 ( .A(KEYINPUT81), .B(G99GAT), .Z(n376) );
  XNOR2_X1 U437 ( .A(G43GAT), .B(G190GAT), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U439 ( .A(n442), .B(n377), .Z(n379) );
  NAND2_X1 U440 ( .A1(G227GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U441 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U442 ( .A(n380), .B(KEYINPUT80), .Z(n383) );
  XNOR2_X1 U443 ( .A(n381), .B(KEYINPUT78), .ZN(n382) );
  XNOR2_X1 U444 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U445 ( .A(n385), .B(n384), .Z(n386) );
  XOR2_X2 U446 ( .A(n387), .B(n386), .Z(n530) );
  NAND2_X1 U447 ( .A1(n388), .A2(n530), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n389), .B(KEYINPUT100), .ZN(n400) );
  NAND2_X1 U449 ( .A1(n476), .A2(n530), .ZN(n390) );
  XOR2_X1 U450 ( .A(KEYINPUT26), .B(n390), .Z(n541) );
  INV_X1 U451 ( .A(n541), .ZN(n565) );
  OR2_X1 U452 ( .A1(n565), .A2(n391), .ZN(n397) );
  XOR2_X1 U453 ( .A(KEYINPUT25), .B(KEYINPUT102), .Z(n395) );
  NOR2_X1 U454 ( .A1(n530), .A2(n519), .ZN(n392) );
  NOR2_X1 U455 ( .A1(n476), .A2(n392), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n393), .B(KEYINPUT101), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n395), .B(n394), .ZN(n396) );
  NAND2_X1 U458 ( .A1(n397), .A2(n396), .ZN(n398) );
  NAND2_X1 U459 ( .A1(n398), .A2(n517), .ZN(n399) );
  NAND2_X1 U460 ( .A1(n400), .A2(n399), .ZN(n484) );
  NAND2_X1 U461 ( .A1(n482), .A2(n484), .ZN(n420) );
  XOR2_X1 U462 ( .A(KEYINPUT11), .B(KEYINPUT74), .Z(n402) );
  XNOR2_X1 U463 ( .A(G134GAT), .B(G106GAT), .ZN(n401) );
  XNOR2_X1 U464 ( .A(n402), .B(n401), .ZN(n419) );
  XOR2_X1 U465 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n404) );
  XNOR2_X1 U466 ( .A(G92GAT), .B(KEYINPUT73), .ZN(n403) );
  XNOR2_X1 U467 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U468 ( .A(G99GAT), .B(G85GAT), .Z(n448) );
  XNOR2_X1 U469 ( .A(n405), .B(n448), .ZN(n407) );
  AND2_X1 U470 ( .A1(G232GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U471 ( .A(n407), .B(n406), .ZN(n412) );
  XOR2_X1 U472 ( .A(G29GAT), .B(G43GAT), .Z(n409) );
  XNOR2_X1 U473 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n408) );
  XNOR2_X1 U474 ( .A(n409), .B(n408), .ZN(n426) );
  XNOR2_X1 U475 ( .A(n426), .B(n410), .ZN(n411) );
  XNOR2_X1 U476 ( .A(n412), .B(n411), .ZN(n414) );
  INV_X1 U477 ( .A(KEYINPUT65), .ZN(n413) );
  XNOR2_X1 U478 ( .A(n414), .B(n413), .ZN(n417) );
  XNOR2_X1 U479 ( .A(n415), .B(KEYINPUT72), .ZN(n416) );
  XNOR2_X1 U480 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U481 ( .A(KEYINPUT36), .B(n560), .Z(n579) );
  XNOR2_X1 U482 ( .A(n421), .B(KEYINPUT37), .ZN(n516) );
  XOR2_X1 U483 ( .A(n423), .B(n422), .Z(n425) );
  XNOR2_X1 U484 ( .A(G36GAT), .B(G50GAT), .ZN(n424) );
  XNOR2_X1 U485 ( .A(n425), .B(n424), .ZN(n430) );
  XOR2_X1 U486 ( .A(n426), .B(KEYINPUT30), .Z(n428) );
  NAND2_X1 U487 ( .A1(G229GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n438) );
  XOR2_X1 U490 ( .A(G8GAT), .B(G113GAT), .Z(n432) );
  XNOR2_X1 U491 ( .A(G169GAT), .B(G197GAT), .ZN(n431) );
  XNOR2_X1 U492 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U493 ( .A(KEYINPUT69), .B(KEYINPUT66), .Z(n434) );
  XNOR2_X1 U494 ( .A(KEYINPUT67), .B(KEYINPUT29), .ZN(n433) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n502) );
  INV_X1 U498 ( .A(n502), .ZN(n566) );
  XOR2_X1 U499 ( .A(n440), .B(n439), .Z(n444) );
  XNOR2_X1 U500 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U501 ( .A(n444), .B(n443), .ZN(n452) );
  XOR2_X1 U502 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n446) );
  XNOR2_X1 U503 ( .A(G204GAT), .B(KEYINPUT33), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U505 ( .A(n448), .B(n447), .Z(n450) );
  NAND2_X1 U506 ( .A1(G230GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U508 ( .A(n452), .B(n451), .ZN(n571) );
  NAND2_X1 U509 ( .A1(n566), .A2(n571), .ZN(n486) );
  NOR2_X1 U510 ( .A1(n516), .A2(n486), .ZN(n453) );
  XOR2_X1 U511 ( .A(KEYINPUT104), .B(n453), .Z(n454) );
  XNOR2_X1 U512 ( .A(KEYINPUT38), .B(n454), .ZN(n499) );
  NOR2_X1 U513 ( .A1(n499), .A2(n530), .ZN(n458) );
  XNOR2_X1 U514 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n456) );
  INV_X1 U515 ( .A(G43GAT), .ZN(n455) );
  OR2_X1 U516 ( .A1(n579), .A2(n482), .ZN(n459) );
  XNOR2_X1 U517 ( .A(KEYINPUT45), .B(n459), .ZN(n461) );
  NAND2_X1 U518 ( .A1(n502), .A2(n571), .ZN(n460) );
  OR2_X1 U519 ( .A1(n461), .A2(n460), .ZN(n470) );
  XOR2_X1 U520 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n463) );
  XNOR2_X1 U521 ( .A(KEYINPUT41), .B(n571), .ZN(n555) );
  NAND2_X1 U522 ( .A1(n555), .A2(n566), .ZN(n462) );
  XNOR2_X1 U523 ( .A(n463), .B(n462), .ZN(n464) );
  NOR2_X1 U524 ( .A1(n574), .A2(n464), .ZN(n465) );
  XNOR2_X1 U525 ( .A(n465), .B(KEYINPUT113), .ZN(n466) );
  NOR2_X1 U526 ( .A1(n560), .A2(n466), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n467), .B(KEYINPUT114), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n468), .B(KEYINPUT47), .ZN(n469) );
  NAND2_X1 U529 ( .A1(n470), .A2(n469), .ZN(n472) );
  INV_X1 U530 ( .A(n526), .ZN(n473) );
  NOR2_X1 U531 ( .A1(n473), .A2(n519), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n474), .B(n292), .ZN(n475) );
  NAND2_X1 U533 ( .A1(n475), .A2(n517), .ZN(n564) );
  NOR2_X1 U534 ( .A1(n476), .A2(n564), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n477), .B(KEYINPUT55), .ZN(n478) );
  NAND2_X1 U536 ( .A1(n561), .A2(n566), .ZN(n481) );
  INV_X1 U537 ( .A(G169GAT), .ZN(n479) );
  NOR2_X1 U538 ( .A1(n560), .A2(n482), .ZN(n483) );
  XNOR2_X1 U539 ( .A(n483), .B(KEYINPUT16), .ZN(n485) );
  NAND2_X1 U540 ( .A1(n485), .A2(n484), .ZN(n503) );
  NOR2_X1 U541 ( .A1(n486), .A2(n503), .ZN(n487) );
  XNOR2_X1 U542 ( .A(KEYINPUT103), .B(n487), .ZN(n493) );
  NOR2_X1 U543 ( .A1(n517), .A2(n493), .ZN(n488) );
  XOR2_X1 U544 ( .A(KEYINPUT34), .B(n488), .Z(n489) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(n489), .ZN(G1324GAT) );
  NOR2_X1 U546 ( .A1(n519), .A2(n493), .ZN(n490) );
  XOR2_X1 U547 ( .A(G8GAT), .B(n490), .Z(G1325GAT) );
  NOR2_X1 U548 ( .A1(n530), .A2(n493), .ZN(n492) );
  XNOR2_X1 U549 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n492), .B(n491), .ZN(G1326GAT) );
  NOR2_X1 U551 ( .A1(n528), .A2(n493), .ZN(n494) );
  XOR2_X1 U552 ( .A(G22GAT), .B(n494), .Z(G1327GAT) );
  NOR2_X1 U553 ( .A1(n517), .A2(n499), .ZN(n497) );
  XOR2_X1 U554 ( .A(KEYINPUT39), .B(KEYINPUT105), .Z(n495) );
  XNOR2_X1 U555 ( .A(G29GAT), .B(n495), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n497), .B(n496), .ZN(G1328GAT) );
  NOR2_X1 U557 ( .A1(n519), .A2(n499), .ZN(n498) );
  XOR2_X1 U558 ( .A(G36GAT), .B(n498), .Z(G1329GAT) );
  NOR2_X1 U559 ( .A1(n528), .A2(n499), .ZN(n501) );
  XNOR2_X1 U560 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(G1331GAT) );
  NAND2_X1 U562 ( .A1(n555), .A2(n502), .ZN(n515) );
  NOR2_X1 U563 ( .A1(n503), .A2(n515), .ZN(n504) );
  XOR2_X1 U564 ( .A(KEYINPUT108), .B(n504), .Z(n511) );
  NOR2_X1 U565 ( .A1(n511), .A2(n517), .ZN(n505) );
  XOR2_X1 U566 ( .A(KEYINPUT42), .B(n505), .Z(n506) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NOR2_X1 U568 ( .A1(n519), .A2(n511), .ZN(n507) );
  XOR2_X1 U569 ( .A(G64GAT), .B(n507), .Z(G1333GAT) );
  XNOR2_X1 U570 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n509) );
  NOR2_X1 U571 ( .A1(n530), .A2(n511), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U573 ( .A(G71GAT), .B(n510), .ZN(G1334GAT) );
  XNOR2_X1 U574 ( .A(KEYINPUT43), .B(KEYINPUT111), .ZN(n513) );
  NOR2_X1 U575 ( .A1(n528), .A2(n511), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U577 ( .A(G78GAT), .B(n514), .Z(G1335GAT) );
  OR2_X1 U578 ( .A1(n516), .A2(n515), .ZN(n522) );
  NOR2_X1 U579 ( .A1(n517), .A2(n522), .ZN(n518) );
  XOR2_X1 U580 ( .A(G85GAT), .B(n518), .Z(G1336GAT) );
  NOR2_X1 U581 ( .A1(n519), .A2(n522), .ZN(n520) );
  XOR2_X1 U582 ( .A(G92GAT), .B(n520), .Z(G1337GAT) );
  NOR2_X1 U583 ( .A1(n530), .A2(n522), .ZN(n521) );
  XOR2_X1 U584 ( .A(G99GAT), .B(n521), .Z(G1338GAT) );
  NOR2_X1 U585 ( .A1(n528), .A2(n522), .ZN(n523) );
  XOR2_X1 U586 ( .A(KEYINPUT44), .B(n523), .Z(n524) );
  XNOR2_X1 U587 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  NAND2_X1 U588 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U589 ( .A(KEYINPUT115), .B(n527), .ZN(n542) );
  NAND2_X1 U590 ( .A1(n528), .A2(n542), .ZN(n529) );
  NOR2_X1 U591 ( .A1(n530), .A2(n529), .ZN(n538) );
  NAND2_X1 U592 ( .A1(n538), .A2(n566), .ZN(n531) );
  XNOR2_X1 U593 ( .A(n531), .B(KEYINPUT116), .ZN(n532) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .Z(n534) );
  NAND2_X1 U596 ( .A1(n538), .A2(n555), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n534), .B(n533), .ZN(G1341GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n536) );
  NAND2_X1 U599 ( .A1(n538), .A2(n574), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U603 ( .A1(n538), .A2(n560), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  NAND2_X1 U605 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U606 ( .A(KEYINPUT118), .B(n543), .Z(n550) );
  NAND2_X1 U607 ( .A1(n566), .A2(n550), .ZN(n544) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(n544), .ZN(G1344GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n546) );
  NAND2_X1 U610 ( .A1(n555), .A2(n550), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(n547), .ZN(G1345GAT) );
  XOR2_X1 U613 ( .A(G155GAT), .B(KEYINPUT119), .Z(n549) );
  NAND2_X1 U614 ( .A1(n574), .A2(n550), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(G1346GAT) );
  NAND2_X1 U616 ( .A1(n550), .A2(n560), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n551), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n553) );
  XNOR2_X1 U619 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U621 ( .A(KEYINPUT56), .B(n554), .Z(n557) );
  NAND2_X1 U622 ( .A1(n561), .A2(n555), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1349GAT) );
  NAND2_X1 U624 ( .A1(n561), .A2(n574), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(KEYINPUT124), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G183GAT), .B(n559), .ZN(G1350GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT58), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(n563), .ZN(G1351GAT) );
  XOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT59), .Z(n568) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n575) );
  NAND2_X1 U632 ( .A1(n575), .A2(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n570) );
  XOR2_X1 U634 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(G204GAT), .B(KEYINPUT61), .Z(n573) );
  INV_X1 U637 ( .A(n575), .ZN(n578) );
  OR2_X1 U638 ( .A1(n578), .A2(n571), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(KEYINPUT126), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G211GAT), .B(n577), .ZN(G1354GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

