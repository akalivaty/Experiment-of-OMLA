//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n452), .B(new_n453), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI21_X1  g033(.A(KEYINPUT69), .B1(new_n454), .B2(G2106), .ZN(new_n459));
  AND3_X1   g034(.A1(new_n454), .A2(KEYINPUT69), .A3(G2106), .ZN(new_n460));
  AOI211_X1 g035(.A(new_n459), .B(new_n460), .C1(G567), .C2(new_n456), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(new_n464), .A3(G101), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(G101), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT70), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n466), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n469), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n466), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n473), .A2(new_n476), .ZN(G160));
  AND2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  OR2_X1    g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n466), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n482), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  OAI211_X1 g065(.A(G138), .B(new_n466), .C1(new_n478), .C2(new_n479), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n493), .A2(new_n466), .A3(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT72), .B1(new_n480), .B2(new_n494), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n493), .A2(new_n466), .A3(G138), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT72), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n471), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n492), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n500), .A2(KEYINPUT71), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(KEYINPUT71), .ZN(new_n502));
  OAI21_X1  g077(.A(G2105), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n503), .A2(new_n505), .B1(new_n485), .B2(G126), .ZN(new_n506));
  AND3_X1   g081(.A1(new_n499), .A2(KEYINPUT73), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(KEYINPUT73), .B1(new_n499), .B2(new_n506), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(KEYINPUT75), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT75), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT5), .A3(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT74), .B(G651), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  OAI21_X1  g097(.A(G543), .B1(new_n518), .B2(new_n519), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G50), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n526), .A2(new_n516), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n522), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(G166));
  NAND2_X1  g104(.A1(new_n524), .A2(G51), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n521), .A2(G89), .ZN(new_n531));
  AND2_X1   g106(.A1(G63), .A2(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n515), .A2(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n530), .A2(new_n531), .A3(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  NAND2_X1  g113(.A1(new_n524), .A2(G52), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n521), .A2(G90), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(new_n516), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND2_X1  g119(.A1(new_n524), .A2(G43), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n521), .A2(G81), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n516), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(new_n515), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n521), .A2(G91), .B1(G651), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n524), .B2(G53), .ZN(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  NOR3_X1   g138(.A1(new_n523), .A2(KEYINPUT9), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n560), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT76), .ZN(G299));
  NAND2_X1  g141(.A1(new_n528), .A2(KEYINPUT77), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n522), .A2(new_n525), .A3(new_n568), .A4(new_n527), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n567), .A2(new_n569), .ZN(G303));
  OAI21_X1  g145(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n571));
  INV_X1    g146(.A(G87), .ZN(new_n572));
  INV_X1    g147(.A(G49), .ZN(new_n573));
  OAI221_X1 g148(.A(new_n571), .B1(new_n520), .B2(new_n572), .C1(new_n573), .C2(new_n523), .ZN(G288));
  NAND2_X1  g149(.A1(new_n521), .A2(G86), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n524), .A2(G48), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n557), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n516), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n575), .A2(new_n576), .A3(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(new_n524), .A2(G47), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n521), .A2(G85), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n583), .B(new_n584), .C1(new_n516), .C2(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  OAI211_X1 g162(.A(G92), .B(new_n515), .C1(new_n518), .C2(new_n519), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT10), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(G651), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(new_n593), .B2(new_n592), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n524), .A2(G54), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n590), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n587), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n587), .B1(new_n598), .B2(G868), .ZN(G321));
  NAND2_X1  g175(.A1(G286), .A2(G868), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT76), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n565), .B(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n601), .B1(new_n603), .B2(G868), .ZN(G297));
  OAI21_X1  g179(.A(new_n601), .B1(new_n603), .B2(G868), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n598), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n598), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n485), .A2(G123), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n466), .A2(G111), .ZN(new_n613));
  OAI21_X1  g188(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(G135), .B2(new_n481), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT79), .Z(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(G2096), .Z(new_n618));
  NAND2_X1  g193(.A1(new_n471), .A2(new_n463), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT13), .B(G2100), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n618), .A2(new_n622), .ZN(G156));
  XOR2_X1   g198(.A(KEYINPUT15), .B(G2435), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2438), .ZN(new_n625));
  XOR2_X1   g200(.A(G2427), .B(G2430), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT80), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n625), .A2(new_n627), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n628), .A2(KEYINPUT14), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2451), .B(G2454), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n630), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G14), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n635), .A2(new_n636), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n638), .A2(new_n639), .ZN(G401));
  XNOR2_X1  g215(.A(G2072), .B(G2078), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT81), .ZN(new_n642));
  XOR2_X1   g217(.A(G2067), .B(G2678), .Z(new_n643));
  XNOR2_X1  g218(.A(G2084), .B(G2090), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT18), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n642), .B(KEYINPUT17), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n643), .B(KEYINPUT82), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n649), .A2(new_n644), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n647), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n649), .B1(KEYINPUT83), .B2(new_n642), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(KEYINPUT83), .B2(new_n642), .ZN(new_n653));
  INV_X1    g228(.A(new_n649), .ZN(new_n654));
  OAI211_X1 g229(.A(new_n653), .B(new_n644), .C1(new_n654), .C2(new_n648), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2100), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT84), .B(G2096), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(G227));
  XOR2_X1   g234(.A(G1971), .B(G1976), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  AND2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT20), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n662), .A2(new_n663), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n661), .A2(new_n664), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n661), .B2(new_n667), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT85), .Z(new_n671));
  XOR2_X1   g246(.A(G1981), .B(G1986), .Z(new_n672));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n671), .B(new_n676), .ZN(G229));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G23), .ZN(new_n679));
  INV_X1    g254(.A(G288), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(new_n678), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT33), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT89), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n682), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n681), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(KEYINPUT89), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT87), .B(G16), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n690), .A2(G22), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(G166), .B2(new_n690), .ZN(new_n692));
  INV_X1    g267(.A(G1971), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G6), .B(G305), .S(G16), .Z(new_n695));
  XOR2_X1   g270(.A(KEYINPUT32), .B(G1981), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND4_X1  g272(.A1(new_n685), .A2(new_n688), .A3(new_n694), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT88), .B(KEYINPUT34), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n698), .A2(new_n700), .ZN(new_n702));
  MUX2_X1   g277(.A(G24), .B(G290), .S(new_n690), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1986), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n485), .A2(G119), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n466), .A2(G107), .ZN(new_n706));
  OAI21_X1  g281(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n707));
  INV_X1    g282(.A(G131), .ZN(new_n708));
  OAI221_X1 g283(.A(new_n705), .B1(new_n706), .B2(new_n707), .C1(new_n708), .C2(new_n472), .ZN(new_n709));
  MUX2_X1   g284(.A(G25), .B(new_n709), .S(G29), .Z(new_n710));
  XOR2_X1   g285(.A(KEYINPUT35), .B(G1991), .Z(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT86), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n710), .B(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n704), .A2(new_n713), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n702), .A2(KEYINPUT90), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(KEYINPUT90), .B1(new_n702), .B2(new_n714), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n701), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT92), .Z(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n678), .A2(G4), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n598), .B2(new_n678), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT93), .B(G1348), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g301(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT26), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n463), .A2(G105), .ZN(new_n729));
  INV_X1    g304(.A(G141), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n472), .B2(new_n730), .ZN(new_n731));
  AOI211_X1 g306(.A(new_n728), .B(new_n731), .C1(G129), .C2(new_n485), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT98), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G29), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n735), .B(KEYINPUT99), .C1(G29), .C2(G32), .ZN(new_n736));
  INV_X1    g311(.A(G29), .ZN(new_n737));
  OR3_X1    g312(.A1(new_n733), .A2(KEYINPUT99), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT27), .B(G1996), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n740), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n736), .A2(new_n742), .A3(new_n738), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n726), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G2072), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n737), .A2(G33), .ZN(new_n746));
  INV_X1    g321(.A(G127), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n480), .A2(new_n747), .ZN(new_n748));
  AND2_X1   g323(.A1(G115), .A2(G2104), .ZN(new_n749));
  OAI21_X1  g324(.A(G2105), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT95), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g327(.A(KEYINPUT95), .B(G2105), .C1(new_n748), .C2(new_n749), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT25), .ZN(new_n754));
  NAND2_X1  g329(.A1(G103), .A2(G2104), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(G2105), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n466), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n481), .A2(G139), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n752), .A2(new_n753), .A3(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT96), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n746), .B1(new_n761), .B2(G29), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n724), .A2(new_n725), .B1(new_n745), .B2(new_n762), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n744), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n689), .A2(G20), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT23), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n603), .B2(new_n678), .ZN(new_n767));
  INV_X1    g342(.A(G1956), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n762), .A2(new_n745), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT97), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT103), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n678), .A2(G5), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G171), .B2(new_n678), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(G1961), .Z(new_n777));
  NAND2_X1  g352(.A1(G160), .A2(G29), .ZN(new_n778));
  INV_X1    g353(.A(G34), .ZN(new_n779));
  AOI21_X1  g354(.A(G29), .B1(new_n779), .B2(KEYINPUT24), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(KEYINPUT24), .B2(new_n779), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G2084), .ZN(new_n783));
  OAI22_X1  g358(.A1(new_n617), .A2(new_n737), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT31), .B(G11), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT100), .B(G28), .ZN(new_n787));
  AOI21_X1  g362(.A(G29), .B1(new_n787), .B2(KEYINPUT30), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(KEYINPUT101), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(KEYINPUT101), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(KEYINPUT30), .B2(new_n787), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n785), .B(new_n786), .C1(new_n789), .C2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G29), .A2(G35), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G162), .B2(G29), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT29), .B(G2090), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n784), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n678), .A2(G21), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G168), .B2(new_n678), .ZN(new_n799));
  INV_X1    g374(.A(G1966), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n737), .A2(G27), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT102), .Z(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G164), .B2(new_n737), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(G2078), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n777), .A2(new_n797), .A3(new_n801), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n690), .A2(G19), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n550), .B2(new_n690), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(G1341), .Z(new_n809));
  OR2_X1    g384(.A1(new_n804), .A2(G2078), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n737), .A2(G26), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT28), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n485), .A2(G128), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n466), .A2(G116), .ZN(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n815));
  INV_X1    g390(.A(G140), .ZN(new_n816));
  OAI221_X1 g391(.A(new_n813), .B1(new_n814), .B2(new_n815), .C1(new_n816), .C2(new_n472), .ZN(new_n817));
  AND3_X1   g392(.A1(new_n817), .A2(KEYINPUT94), .A3(G29), .ZN(new_n818));
  AOI21_X1  g393(.A(KEYINPUT94), .B1(new_n817), .B2(G29), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n812), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(G2067), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n809), .A2(new_n810), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n806), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n764), .A2(new_n773), .A3(new_n774), .A4(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n744), .A2(new_n763), .A3(new_n824), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT103), .B1(new_n826), .B2(new_n772), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n701), .B(new_n719), .C1(new_n715), .C2(new_n716), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n721), .A2(new_n828), .A3(new_n829), .ZN(G150));
  INV_X1    g405(.A(G150), .ZN(G311));
  NOR2_X1   g406(.A1(new_n597), .A2(new_n606), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n515), .A2(G67), .ZN(new_n835));
  AND2_X1   g410(.A1(G80), .A2(G543), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n580), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT105), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT106), .B(G55), .Z(new_n841));
  NAND2_X1  g416(.A1(new_n524), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n521), .A2(G93), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n839), .A2(new_n840), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n549), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n834), .B(new_n845), .Z(new_n846));
  AND2_X1   g421(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n847), .A2(new_n848), .A3(G860), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n844), .A2(G860), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT37), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n849), .A2(new_n851), .ZN(G145));
  NAND2_X1  g427(.A1(new_n761), .A2(new_n732), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n734), .B2(new_n761), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n499), .A2(new_n506), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(new_n817), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n854), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n485), .A2(G130), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n466), .A2(G118), .ZN(new_n859));
  OAI21_X1  g434(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n860));
  INV_X1    g435(.A(G142), .ZN(new_n861));
  OAI221_X1 g436(.A(new_n858), .B1(new_n859), .B2(new_n860), .C1(new_n861), .C2(new_n472), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT107), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n620), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n709), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n857), .A2(KEYINPUT108), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(KEYINPUT108), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n867), .B2(new_n857), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n617), .B(new_n489), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(G160), .Z(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(G37), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n870), .B(new_n866), .C1(new_n867), .C2(new_n857), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g451(.A(G868), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n844), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT109), .ZN(new_n879));
  XNOR2_X1  g454(.A(G288), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(G305), .ZN(new_n881));
  XNOR2_X1  g456(.A(G166), .B(G290), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT110), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT42), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n603), .A2(new_n597), .ZN(new_n887));
  NAND2_X1  g462(.A1(G299), .A2(new_n598), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT41), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n887), .A2(new_n888), .A3(KEYINPUT41), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n845), .B(new_n608), .Z(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n889), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n895), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n886), .B(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n878), .B1(new_n898), .B2(new_n877), .ZN(G295));
  OAI21_X1  g474(.A(new_n878), .B1(new_n898), .B2(new_n877), .ZN(G331));
  XNOR2_X1  g475(.A(KEYINPUT111), .B(KEYINPUT44), .ZN(new_n901));
  XNOR2_X1  g476(.A(G301), .B(G286), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n845), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n845), .A2(new_n902), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n905), .A2(KEYINPUT112), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT112), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n907), .B1(new_n845), .B2(new_n902), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n904), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n896), .A2(new_n903), .ZN(new_n910));
  AOI22_X1  g485(.A1(new_n893), .A2(new_n909), .B1(new_n910), .B2(new_n905), .ZN(new_n911));
  INV_X1    g486(.A(new_n883), .ZN(new_n912));
  AOI21_X1  g487(.A(G37), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n906), .A2(new_n908), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n915), .A2(new_n896), .A3(new_n903), .ZN(new_n916));
  AOI22_X1  g491(.A1(new_n891), .A2(new_n892), .B1(new_n904), .B2(new_n905), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n883), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n913), .A2(new_n914), .A3(new_n918), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n911), .A2(new_n912), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n914), .B1(new_n920), .B2(new_n913), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n901), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n914), .A3(new_n913), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n913), .A2(new_n918), .ZN(new_n924));
  OAI211_X1 g499(.A(KEYINPUT44), .B(new_n923), .C1(new_n924), .C2(new_n914), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(G397));
  XOR2_X1   g501(.A(KEYINPUT113), .B(G1384), .Z(new_n927));
  AOI21_X1  g502(.A(KEYINPUT45), .B1(new_n855), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(G40), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n473), .A2(new_n476), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n931), .A2(G1996), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n933), .A2(new_n733), .ZN(new_n934));
  XOR2_X1   g509(.A(new_n934), .B(KEYINPUT114), .Z(new_n935));
  INV_X1    g510(.A(new_n931), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n817), .B(new_n821), .ZN(new_n937));
  INV_X1    g512(.A(G1996), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n937), .B1(new_n732), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n935), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n711), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n709), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n709), .A2(new_n941), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n936), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(G290), .B(G1986), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n945), .B1(new_n936), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT61), .ZN(new_n948));
  XOR2_X1   g523(.A(new_n565), .B(KEYINPUT57), .Z(new_n949));
  AOI21_X1  g524(.A(G1384), .B1(new_n499), .B2(new_n506), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT50), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n930), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT116), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT116), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n954), .B(new_n930), .C1(new_n950), .C2(new_n951), .ZN(new_n955));
  INV_X1    g530(.A(G1384), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n951), .B(new_n956), .C1(new_n507), .C2(new_n508), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n953), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n768), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT120), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT120), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n961), .A3(new_n768), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n956), .B1(new_n507), .B2(new_n508), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n855), .A2(KEYINPUT45), .A3(new_n927), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n967), .A2(new_n930), .ZN(new_n968));
  XNOR2_X1  g543(.A(KEYINPUT56), .B(G2072), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n949), .B1(new_n963), .B2(new_n970), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n958), .A2(new_n961), .A3(new_n768), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n961), .B1(new_n958), .B2(new_n768), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n949), .B(new_n970), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n948), .B1(new_n971), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT59), .ZN(new_n977));
  XNOR2_X1  g552(.A(KEYINPUT121), .B(G1996), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n966), .A2(new_n968), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n930), .A2(new_n950), .ZN(new_n981));
  XOR2_X1   g556(.A(KEYINPUT58), .B(G1341), .Z(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n977), .B1(new_n984), .B2(new_n550), .ZN(new_n985));
  AOI211_X1 g560(.A(KEYINPUT59), .B(new_n549), .C1(new_n980), .C2(new_n983), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n481), .A2(G137), .B1(new_n468), .B2(new_n465), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n474), .A2(new_n475), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n987), .B(G40), .C1(new_n466), .C2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n951), .B2(new_n950), .ZN(new_n990));
  INV_X1    g565(.A(new_n508), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n499), .A2(KEYINPUT73), .A3(new_n506), .ZN(new_n992));
  AOI21_X1  g567(.A(G1384), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n990), .B1(new_n993), .B2(new_n951), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n725), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT60), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(new_n598), .B2(KEYINPUT122), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n930), .A2(new_n950), .A3(new_n821), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n995), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n598), .A2(KEYINPUT122), .ZN(new_n1000));
  OAI22_X1  g575(.A1(new_n985), .A2(new_n986), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n1000), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT60), .B1(new_n995), .B2(new_n998), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(new_n1006));
  INV_X1    g581(.A(new_n949), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1008), .A2(KEYINPUT61), .A3(new_n974), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n976), .A2(new_n1005), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n597), .B1(new_n995), .B2(new_n998), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n974), .B1(new_n971), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT125), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT123), .ZN(new_n1015));
  OAI211_X1 g590(.A(KEYINPUT45), .B(new_n956), .C1(new_n507), .C2(new_n508), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n855), .A2(new_n956), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n989), .B1(new_n1017), .B2(new_n965), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1015), .B1(new_n1019), .B2(G2078), .ZN(new_n1020));
  INV_X1    g595(.A(G2078), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1016), .A2(new_n1018), .A3(KEYINPUT123), .A4(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1020), .A2(KEYINPUT53), .A3(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n966), .A2(new_n1021), .A3(new_n968), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT124), .B(G1961), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1024), .A2(new_n1025), .B1(new_n994), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1014), .B1(new_n1028), .B2(G171), .ZN(new_n1029));
  AOI211_X1 g604(.A(KEYINPUT125), .B(G301), .C1(new_n1023), .C2(new_n1027), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n994), .A2(new_n1026), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n928), .A2(new_n1025), .A3(G2078), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n968), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1031), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(G171), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1029), .A2(new_n1030), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT126), .B1(new_n1037), .B2(KEYINPUT54), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n567), .A2(G8), .A3(new_n569), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n1039), .B(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(G1971), .B1(new_n966), .B2(new_n968), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n1044));
  AOI21_X1  g619(.A(G2090), .B1(new_n958), .B2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n953), .A2(KEYINPUT117), .A3(new_n955), .A4(new_n957), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(G8), .B1(new_n1047), .B2(KEYINPUT118), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n1049));
  AOI211_X1 g624(.A(new_n1049), .B(new_n1043), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1042), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G2090), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1052), .B(new_n990), .C1(new_n993), .C2(new_n951), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT115), .B1(new_n1054), .B2(new_n1043), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n966), .A2(new_n968), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1056), .B(new_n1053), .C1(new_n1057), .C2(G1971), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1041), .A2(new_n1055), .A3(new_n1058), .A4(G8), .ZN(new_n1059));
  NAND2_X1  g634(.A1(G305), .A2(G1981), .ZN(new_n1060));
  INV_X1    g635(.A(G1981), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n575), .A2(new_n576), .A3(new_n1061), .A4(new_n581), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT49), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1060), .A2(KEYINPUT49), .A3(new_n1062), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n981), .A2(G8), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1067), .B1(G1976), .B2(new_n680), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1070), .B(new_n1071), .C1(G1976), .C2(new_n680), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1069), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1059), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1019), .A2(new_n800), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1077), .B(G168), .C1(G2084), .C2(new_n994), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(G8), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n951), .A3(new_n956), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n930), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(KEYINPUT50), .B2(new_n964), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1082), .A2(new_n783), .B1(new_n1019), .B2(new_n800), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(G168), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT51), .B1(new_n1079), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G8), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1086), .B1(new_n1083), .B2(G168), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT51), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n1035), .B2(G171), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(G171), .B2(new_n1028), .ZN(new_n1093));
  AND4_X1   g668(.A1(new_n1051), .A2(new_n1076), .A3(new_n1090), .A4(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT126), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1028), .A2(G171), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT125), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1028), .A2(new_n1014), .A3(G171), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1095), .B(new_n1091), .C1(new_n1099), .C2(new_n1036), .ZN(new_n1100));
  AND4_X1   g675(.A1(new_n1013), .A2(new_n1038), .A3(new_n1094), .A4(new_n1100), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1083), .A2(new_n1086), .A3(G286), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1051), .A2(new_n1076), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT63), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1059), .A2(KEYINPUT63), .A3(new_n1102), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1055), .A2(new_n1058), .A3(G8), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n1042), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1107), .B1(new_n1109), .B2(new_n1075), .ZN(new_n1110));
  AOI211_X1 g685(.A(KEYINPUT119), .B(new_n1074), .C1(new_n1108), .C2(new_n1042), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1106), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1105), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(G288), .A2(G1976), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1069), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1062), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1068), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n1059), .B2(new_n1074), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1077), .B1(new_n994), .B2(G2084), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(G286), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1088), .B1(new_n1087), .B2(new_n1121), .ZN(new_n1122));
  AOI211_X1 g697(.A(KEYINPUT51), .B(new_n1086), .C1(new_n1083), .C2(G168), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1119), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1085), .A2(KEYINPUT62), .A3(new_n1089), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1124), .A2(new_n1125), .B1(new_n1098), .B2(new_n1097), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1059), .A2(new_n1075), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1049), .B1(new_n1128), .B2(new_n1043), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1047), .A2(KEYINPUT118), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(G8), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1127), .B1(new_n1131), .B2(new_n1042), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1118), .B1(new_n1126), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1113), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n947), .B1(new_n1101), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n931), .B1(new_n732), .B2(new_n937), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n933), .A2(KEYINPUT46), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n933), .A2(KEYINPUT46), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT47), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n940), .A2(new_n943), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n817), .A2(G2067), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n931), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n945), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n931), .A2(G290), .A3(G1986), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1145), .B(KEYINPUT48), .Z(new_n1146));
  AOI211_X1 g721(.A(new_n1140), .B(new_n1143), .C1(new_n1144), .C2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1135), .A2(new_n1147), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g723(.A(G319), .B1(new_n638), .B2(new_n639), .ZN(new_n1150));
  OR2_X1    g724(.A1(G229), .A2(new_n1150), .ZN(new_n1151));
  OR3_X1    g725(.A1(new_n1151), .A2(KEYINPUT127), .A3(G227), .ZN(new_n1152));
  OAI21_X1  g726(.A(KEYINPUT127), .B1(new_n1151), .B2(G227), .ZN(new_n1153));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  OAI211_X1 g728(.A(new_n875), .B(new_n1154), .C1(new_n919), .C2(new_n921), .ZN(G225));
  INV_X1    g729(.A(G225), .ZN(G308));
endmodule


