

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U553 ( .A1(n598), .A2(G2104), .ZN(n895) );
  AND2_X1 U554 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U555 ( .A1(n680), .A2(KEYINPUT33), .ZN(n681) );
  NOR2_X1 U556 ( .A1(n696), .A2(n695), .ZN(n704) );
  XOR2_X1 U557 ( .A(n613), .B(KEYINPUT65), .Z(n518) );
  AND2_X1 U558 ( .A1(n600), .A2(n599), .ZN(n519) );
  AND2_X1 U559 ( .A1(n741), .A2(n740), .ZN(n520) );
  AND2_X1 U560 ( .A1(n738), .A2(n754), .ZN(n521) );
  AND2_X1 U561 ( .A1(n650), .A2(n649), .ZN(n522) );
  INV_X1 U562 ( .A(n650), .ZN(n662) );
  NOR2_X1 U563 ( .A1(n982), .A2(n620), .ZN(n625) );
  INV_X1 U564 ( .A(KEYINPUT31), .ZN(n658) );
  INV_X1 U565 ( .A(n981), .ZN(n680) );
  INV_X1 U566 ( .A(KEYINPUT32), .ZN(n670) );
  OR2_X2 U567 ( .A1(n719), .A2(n720), .ZN(n650) );
  NOR2_X1 U568 ( .A1(n739), .A2(n521), .ZN(n740) );
  INV_X1 U569 ( .A(KEYINPUT17), .ZN(n593) );
  XOR2_X1 U570 ( .A(KEYINPUT75), .B(n582), .Z(n972) );
  NAND2_X1 U571 ( .A1(n894), .A2(G138), .ZN(n596) );
  NOR2_X1 U572 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U573 ( .A1(G651), .A2(n555), .ZN(n791) );
  XOR2_X1 U574 ( .A(KEYINPUT1), .B(n529), .Z(n790) );
  XNOR2_X1 U575 ( .A(KEYINPUT9), .B(KEYINPUT71), .ZN(n527) );
  XOR2_X1 U576 ( .A(KEYINPUT0), .B(G543), .Z(n555) );
  INV_X1 U577 ( .A(G651), .ZN(n528) );
  NOR2_X1 U578 ( .A1(n555), .A2(n528), .ZN(n794) );
  NAND2_X1 U579 ( .A1(n794), .A2(G77), .ZN(n523) );
  XNOR2_X1 U580 ( .A(n523), .B(KEYINPUT70), .ZN(n525) );
  NOR2_X1 U581 ( .A1(G651), .A2(G543), .ZN(n796) );
  NAND2_X1 U582 ( .A1(G90), .A2(n796), .ZN(n524) );
  NAND2_X1 U583 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U584 ( .A(n527), .B(n526), .ZN(n534) );
  NOR2_X1 U585 ( .A1(G543), .A2(n528), .ZN(n529) );
  NAND2_X1 U586 ( .A1(G64), .A2(n790), .ZN(n531) );
  NAND2_X1 U587 ( .A1(G52), .A2(n791), .ZN(n530) );
  NAND2_X1 U588 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U589 ( .A(KEYINPUT69), .B(n532), .Z(n533) );
  NOR2_X1 U590 ( .A1(n534), .A2(n533), .ZN(G171) );
  NAND2_X1 U591 ( .A1(n796), .A2(G89), .ZN(n535) );
  XNOR2_X1 U592 ( .A(n535), .B(KEYINPUT4), .ZN(n537) );
  NAND2_X1 U593 ( .A1(G76), .A2(n794), .ZN(n536) );
  NAND2_X1 U594 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U595 ( .A(KEYINPUT5), .B(n538), .ZN(n544) );
  NAND2_X1 U596 ( .A1(n790), .A2(G63), .ZN(n539) );
  XOR2_X1 U597 ( .A(KEYINPUT77), .B(n539), .Z(n541) );
  NAND2_X1 U598 ( .A1(n791), .A2(G51), .ZN(n540) );
  NAND2_X1 U599 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U600 ( .A(KEYINPUT6), .B(n542), .Z(n543) );
  NAND2_X1 U601 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U602 ( .A(KEYINPUT7), .B(n545), .ZN(G168) );
  XOR2_X1 U603 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U604 ( .A1(G75), .A2(n794), .ZN(n547) );
  NAND2_X1 U605 ( .A1(G88), .A2(n796), .ZN(n546) );
  NAND2_X1 U606 ( .A1(n547), .A2(n546), .ZN(n551) );
  NAND2_X1 U607 ( .A1(G62), .A2(n790), .ZN(n549) );
  NAND2_X1 U608 ( .A1(G50), .A2(n791), .ZN(n548) );
  NAND2_X1 U609 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U610 ( .A1(n551), .A2(n550), .ZN(G166) );
  INV_X1 U611 ( .A(G166), .ZN(G303) );
  NAND2_X1 U612 ( .A1(G49), .A2(n791), .ZN(n553) );
  NAND2_X1 U613 ( .A1(G74), .A2(G651), .ZN(n552) );
  NAND2_X1 U614 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U615 ( .A1(n790), .A2(n554), .ZN(n557) );
  NAND2_X1 U616 ( .A1(n555), .A2(G87), .ZN(n556) );
  NAND2_X1 U617 ( .A1(n557), .A2(n556), .ZN(G288) );
  NAND2_X1 U618 ( .A1(G86), .A2(n796), .ZN(n559) );
  NAND2_X1 U619 ( .A1(G61), .A2(n790), .ZN(n558) );
  NAND2_X1 U620 ( .A1(n559), .A2(n558), .ZN(n562) );
  NAND2_X1 U621 ( .A1(n794), .A2(G73), .ZN(n560) );
  XOR2_X1 U622 ( .A(KEYINPUT2), .B(n560), .Z(n561) );
  NOR2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n564) );
  NAND2_X1 U624 ( .A1(n791), .A2(G48), .ZN(n563) );
  NAND2_X1 U625 ( .A1(n564), .A2(n563), .ZN(G305) );
  NAND2_X1 U626 ( .A1(n794), .A2(G72), .ZN(n565) );
  XNOR2_X1 U627 ( .A(n565), .B(KEYINPUT66), .ZN(n567) );
  NAND2_X1 U628 ( .A1(G85), .A2(n796), .ZN(n566) );
  NAND2_X1 U629 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U630 ( .A(KEYINPUT67), .B(n568), .ZN(n573) );
  NAND2_X1 U631 ( .A1(G60), .A2(n790), .ZN(n570) );
  NAND2_X1 U632 ( .A1(G47), .A2(n791), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U634 ( .A(KEYINPUT68), .B(n571), .Z(n572) );
  NAND2_X1 U635 ( .A1(n573), .A2(n572), .ZN(G290) );
  NAND2_X1 U636 ( .A1(G54), .A2(n791), .ZN(n580) );
  NAND2_X1 U637 ( .A1(G79), .A2(n794), .ZN(n575) );
  NAND2_X1 U638 ( .A1(G66), .A2(n790), .ZN(n574) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n796), .A2(G92), .ZN(n576) );
  XOR2_X1 U641 ( .A(KEYINPUT74), .B(n576), .Z(n577) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U643 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U644 ( .A(n581), .B(KEYINPUT15), .ZN(n582) );
  NAND2_X1 U645 ( .A1(n796), .A2(G81), .ZN(n583) );
  XNOR2_X1 U646 ( .A(n583), .B(KEYINPUT12), .ZN(n585) );
  NAND2_X1 U647 ( .A1(G68), .A2(n794), .ZN(n584) );
  NAND2_X1 U648 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U649 ( .A(KEYINPUT13), .B(n586), .Z(n590) );
  NAND2_X1 U650 ( .A1(G56), .A2(n790), .ZN(n587) );
  XNOR2_X1 U651 ( .A(n587), .B(KEYINPUT14), .ZN(n588) );
  XNOR2_X1 U652 ( .A(n588), .B(KEYINPUT73), .ZN(n589) );
  NOR2_X1 U653 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U654 ( .A1(n791), .A2(G43), .ZN(n591) );
  NAND2_X1 U655 ( .A1(n592), .A2(n591), .ZN(n982) );
  NOR2_X1 U656 ( .A1(G2105), .A2(G2104), .ZN(n594) );
  XNOR2_X2 U657 ( .A(n594), .B(n593), .ZN(n894) );
  INV_X1 U658 ( .A(KEYINPUT90), .ZN(n595) );
  XNOR2_X1 U659 ( .A(n596), .B(n595), .ZN(n603) );
  AND2_X1 U660 ( .A1(G2105), .A2(G2104), .ZN(n710) );
  NAND2_X1 U661 ( .A1(G114), .A2(n710), .ZN(n597) );
  XOR2_X1 U662 ( .A(KEYINPUT89), .B(n597), .Z(n601) );
  INV_X1 U663 ( .A(G2105), .ZN(n598) );
  NOR2_X1 U664 ( .A1(n598), .A2(G2104), .ZN(n607) );
  BUF_X1 U665 ( .A(n607), .Z(n899) );
  NAND2_X1 U666 ( .A1(G126), .A2(n899), .ZN(n600) );
  NAND2_X1 U667 ( .A1(G102), .A2(n895), .ZN(n599) );
  NAND2_X1 U668 ( .A1(n601), .A2(n519), .ZN(n602) );
  NOR2_X1 U669 ( .A1(n603), .A2(n602), .ZN(n761) );
  NOR2_X1 U670 ( .A1(n761), .A2(G1384), .ZN(n604) );
  INV_X1 U671 ( .A(n604), .ZN(n719) );
  NAND2_X1 U672 ( .A1(G113), .A2(n710), .ZN(n606) );
  NAND2_X1 U673 ( .A1(G137), .A2(n894), .ZN(n605) );
  AND2_X1 U674 ( .A1(n606), .A2(n605), .ZN(n760) );
  AND2_X1 U675 ( .A1(n760), .A2(G40), .ZN(n614) );
  INV_X1 U676 ( .A(KEYINPUT64), .ZN(n609) );
  NAND2_X1 U677 ( .A1(n607), .A2(G125), .ZN(n608) );
  XNOR2_X1 U678 ( .A(n609), .B(n608), .ZN(n612) );
  NAND2_X1 U679 ( .A1(n895), .A2(G101), .ZN(n610) );
  XNOR2_X1 U680 ( .A(KEYINPUT23), .B(n610), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n614), .A2(n518), .ZN(n720) );
  INV_X1 U682 ( .A(n650), .ZN(n615) );
  NAND2_X1 U683 ( .A1(G1996), .A2(n615), .ZN(n616) );
  XNOR2_X1 U684 ( .A(n616), .B(KEYINPUT26), .ZN(n618) );
  NAND2_X1 U685 ( .A1(G1341), .A2(n650), .ZN(n617) );
  NAND2_X1 U686 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U687 ( .A(n619), .B(KEYINPUT100), .ZN(n620) );
  NAND2_X1 U688 ( .A1(n972), .A2(n625), .ZN(n624) );
  NOR2_X1 U689 ( .A1(n662), .A2(G1348), .ZN(n622) );
  NOR2_X1 U690 ( .A1(G2067), .A2(n650), .ZN(n621) );
  NOR2_X1 U691 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U692 ( .A1(n624), .A2(n623), .ZN(n627) );
  OR2_X1 U693 ( .A1(n972), .A2(n625), .ZN(n626) );
  NAND2_X1 U694 ( .A1(n627), .A2(n626), .ZN(n638) );
  NAND2_X1 U695 ( .A1(G65), .A2(n790), .ZN(n629) );
  NAND2_X1 U696 ( .A1(G53), .A2(n791), .ZN(n628) );
  NAND2_X1 U697 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U698 ( .A1(G78), .A2(n794), .ZN(n631) );
  NAND2_X1 U699 ( .A1(G91), .A2(n796), .ZN(n630) );
  NAND2_X1 U700 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U701 ( .A1(n633), .A2(n632), .ZN(n983) );
  NAND2_X1 U702 ( .A1(n662), .A2(G2072), .ZN(n634) );
  XNOR2_X1 U703 ( .A(n634), .B(KEYINPUT27), .ZN(n636) );
  INV_X1 U704 ( .A(G1956), .ZN(n847) );
  NOR2_X1 U705 ( .A1(n847), .A2(n662), .ZN(n635) );
  NOR2_X1 U706 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U707 ( .A1(n983), .A2(n639), .ZN(n637) );
  NAND2_X1 U708 ( .A1(n638), .A2(n637), .ZN(n642) );
  NOR2_X1 U709 ( .A1(n983), .A2(n639), .ZN(n640) );
  XOR2_X1 U710 ( .A(n640), .B(KEYINPUT28), .Z(n641) );
  NAND2_X1 U711 ( .A1(n642), .A2(n641), .ZN(n644) );
  INV_X1 U712 ( .A(KEYINPUT29), .ZN(n643) );
  XNOR2_X1 U713 ( .A(n644), .B(n643), .ZN(n648) );
  XNOR2_X1 U714 ( .A(G2078), .B(KEYINPUT25), .ZN(n957) );
  NOR2_X1 U715 ( .A1(n650), .A2(n957), .ZN(n646) );
  INV_X1 U716 ( .A(G1961), .ZN(n971) );
  NOR2_X1 U717 ( .A1(n662), .A2(n971), .ZN(n645) );
  NOR2_X1 U718 ( .A1(n646), .A2(n645), .ZN(n655) );
  NAND2_X1 U719 ( .A1(G171), .A2(n655), .ZN(n647) );
  NAND2_X1 U720 ( .A1(n648), .A2(n647), .ZN(n661) );
  NOR2_X1 U721 ( .A1(n667), .A2(G1966), .ZN(n649) );
  NOR2_X1 U722 ( .A1(G2084), .A2(n650), .ZN(n672) );
  NOR2_X1 U723 ( .A1(n522), .A2(n672), .ZN(n651) );
  NAND2_X1 U724 ( .A1(G8), .A2(n651), .ZN(n652) );
  XNOR2_X1 U725 ( .A(KEYINPUT101), .B(n652), .ZN(n653) );
  XOR2_X1 U726 ( .A(KEYINPUT30), .B(n653), .Z(n654) );
  NOR2_X1 U727 ( .A1(G168), .A2(n654), .ZN(n657) );
  NOR2_X1 U728 ( .A1(G171), .A2(n655), .ZN(n656) );
  NOR2_X1 U729 ( .A1(n657), .A2(n656), .ZN(n659) );
  XNOR2_X1 U730 ( .A(n659), .B(n658), .ZN(n660) );
  NAND2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n673) );
  NAND2_X1 U732 ( .A1(n673), .A2(G286), .ZN(n669) );
  INV_X1 U733 ( .A(G8), .ZN(n667) );
  OR2_X1 U734 ( .A1(n667), .A2(n662), .ZN(n702) );
  NOR2_X1 U735 ( .A1(G1971), .A2(n702), .ZN(n664) );
  NOR2_X1 U736 ( .A1(G2090), .A2(n650), .ZN(n663) );
  NOR2_X1 U737 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U738 ( .A1(n665), .A2(G303), .ZN(n666) );
  OR2_X1 U739 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U740 ( .A1(n669), .A2(n668), .ZN(n671) );
  XNOR2_X1 U741 ( .A(n671), .B(n670), .ZN(n678) );
  NAND2_X1 U742 ( .A1(n672), .A2(G8), .ZN(n676) );
  INV_X1 U743 ( .A(n673), .ZN(n674) );
  NOR2_X1 U744 ( .A1(n522), .A2(n674), .ZN(n675) );
  NAND2_X1 U745 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U746 ( .A1(n678), .A2(n677), .ZN(n699) );
  NOR2_X1 U747 ( .A1(G1976), .A2(G288), .ZN(n685) );
  NOR2_X1 U748 ( .A1(G1971), .A2(G303), .ZN(n679) );
  NOR2_X1 U749 ( .A1(n685), .A2(n679), .ZN(n987) );
  NAND2_X1 U750 ( .A1(n699), .A2(n987), .ZN(n682) );
  NAND2_X1 U751 ( .A1(G1976), .A2(G288), .ZN(n981) );
  INV_X1 U752 ( .A(n702), .ZN(n684) );
  NAND2_X1 U753 ( .A1(n683), .A2(n684), .ZN(n688) );
  NAND2_X1 U754 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U755 ( .A1(n686), .A2(KEYINPUT33), .ZN(n687) );
  NAND2_X1 U756 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U757 ( .A(KEYINPUT102), .B(n689), .ZN(n690) );
  XOR2_X1 U758 ( .A(G1981), .B(G305), .Z(n977) );
  NAND2_X1 U759 ( .A1(n690), .A2(n977), .ZN(n691) );
  XNOR2_X1 U760 ( .A(n691), .B(KEYINPUT103), .ZN(n696) );
  NOR2_X1 U761 ( .A1(G1981), .A2(G305), .ZN(n692) );
  XNOR2_X1 U762 ( .A(n692), .B(KEYINPUT24), .ZN(n693) );
  XNOR2_X1 U763 ( .A(n693), .B(KEYINPUT99), .ZN(n694) );
  NOR2_X1 U764 ( .A1(n702), .A2(n694), .ZN(n695) );
  NOR2_X1 U765 ( .A1(G2090), .A2(G303), .ZN(n697) );
  NAND2_X1 U766 ( .A1(G8), .A2(n697), .ZN(n698) );
  NAND2_X1 U767 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U768 ( .A(KEYINPUT104), .B(n700), .ZN(n701) );
  NAND2_X1 U769 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n741) );
  XNOR2_X1 U771 ( .A(KEYINPUT37), .B(G2067), .ZN(n752) );
  XNOR2_X1 U772 ( .A(KEYINPUT95), .B(KEYINPUT36), .ZN(n718) );
  NAND2_X1 U773 ( .A1(n894), .A2(G140), .ZN(n705) );
  XNOR2_X1 U774 ( .A(n705), .B(KEYINPUT92), .ZN(n707) );
  NAND2_X1 U775 ( .A1(G104), .A2(n895), .ZN(n706) );
  NAND2_X1 U776 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U777 ( .A(n708), .B(KEYINPUT93), .ZN(n709) );
  XNOR2_X1 U778 ( .A(n709), .B(KEYINPUT34), .ZN(n716) );
  XNOR2_X1 U779 ( .A(KEYINPUT94), .B(KEYINPUT35), .ZN(n714) );
  NAND2_X1 U780 ( .A1(G128), .A2(n899), .ZN(n712) );
  NAND2_X1 U781 ( .A1(G116), .A2(n710), .ZN(n711) );
  NAND2_X1 U782 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U783 ( .A(n714), .B(n713), .ZN(n715) );
  NAND2_X1 U784 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U785 ( .A(n718), .B(n717), .ZN(n874) );
  NOR2_X1 U786 ( .A1(n752), .A2(n874), .ZN(n943) );
  NOR2_X1 U787 ( .A1(n604), .A2(n720), .ZN(n721) );
  XOR2_X1 U788 ( .A(KEYINPUT91), .B(n721), .Z(n754) );
  NAND2_X1 U789 ( .A1(n943), .A2(n754), .ZN(n750) );
  INV_X1 U790 ( .A(n750), .ZN(n739) );
  NAND2_X1 U791 ( .A1(n895), .A2(G105), .ZN(n723) );
  XNOR2_X1 U792 ( .A(KEYINPUT98), .B(KEYINPUT38), .ZN(n722) );
  XNOR2_X1 U793 ( .A(n723), .B(n722), .ZN(n730) );
  NAND2_X1 U794 ( .A1(G129), .A2(n899), .ZN(n725) );
  NAND2_X1 U795 ( .A1(G141), .A2(n894), .ZN(n724) );
  NAND2_X1 U796 ( .A1(n725), .A2(n724), .ZN(n728) );
  NAND2_X1 U797 ( .A1(G117), .A2(n710), .ZN(n726) );
  XNOR2_X1 U798 ( .A(KEYINPUT97), .B(n726), .ZN(n727) );
  NOR2_X1 U799 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U800 ( .A1(n730), .A2(n729), .ZN(n877) );
  AND2_X1 U801 ( .A1(n877), .A2(G1996), .ZN(n929) );
  NAND2_X1 U802 ( .A1(G119), .A2(n899), .ZN(n732) );
  NAND2_X1 U803 ( .A1(G131), .A2(n894), .ZN(n731) );
  NAND2_X1 U804 ( .A1(n732), .A2(n731), .ZN(n735) );
  NAND2_X1 U805 ( .A1(n895), .A2(G95), .ZN(n733) );
  XOR2_X1 U806 ( .A(KEYINPUT96), .B(n733), .Z(n734) );
  NOR2_X1 U807 ( .A1(n735), .A2(n734), .ZN(n737) );
  NAND2_X1 U808 ( .A1(n710), .A2(G107), .ZN(n736) );
  NAND2_X1 U809 ( .A1(n737), .A2(n736), .ZN(n873) );
  AND2_X1 U810 ( .A1(n873), .A2(G1991), .ZN(n931) );
  OR2_X1 U811 ( .A1(n929), .A2(n931), .ZN(n738) );
  XNOR2_X1 U812 ( .A(G1986), .B(G290), .ZN(n993) );
  NAND2_X1 U813 ( .A1(n993), .A2(n754), .ZN(n742) );
  NAND2_X1 U814 ( .A1(n520), .A2(n742), .ZN(n757) );
  XOR2_X1 U815 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n749) );
  NOR2_X1 U816 ( .A1(G1996), .A2(n877), .ZN(n743) );
  XOR2_X1 U817 ( .A(KEYINPUT105), .B(n743), .Z(n926) );
  NOR2_X1 U818 ( .A1(G1986), .A2(G290), .ZN(n744) );
  XNOR2_X1 U819 ( .A(n744), .B(KEYINPUT106), .ZN(n745) );
  NOR2_X1 U820 ( .A1(G1991), .A2(n873), .ZN(n930) );
  NOR2_X1 U821 ( .A1(n745), .A2(n930), .ZN(n746) );
  NOR2_X1 U822 ( .A1(n521), .A2(n746), .ZN(n747) );
  NOR2_X1 U823 ( .A1(n926), .A2(n747), .ZN(n748) );
  XNOR2_X1 U824 ( .A(n749), .B(n748), .ZN(n751) );
  NAND2_X1 U825 ( .A1(n751), .A2(n750), .ZN(n753) );
  NAND2_X1 U826 ( .A1(n752), .A2(n874), .ZN(n940) );
  NAND2_X1 U827 ( .A1(n753), .A2(n940), .ZN(n755) );
  NAND2_X1 U828 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U829 ( .A1(n757), .A2(n756), .ZN(n759) );
  XNOR2_X1 U830 ( .A(KEYINPUT40), .B(KEYINPUT108), .ZN(n758) );
  XNOR2_X1 U831 ( .A(n759), .B(n758), .ZN(G329) );
  AND2_X1 U832 ( .A1(n760), .A2(n518), .ZN(G160) );
  INV_X1 U833 ( .A(G57), .ZN(G237) );
  INV_X1 U834 ( .A(G132), .ZN(G219) );
  INV_X1 U835 ( .A(G82), .ZN(G220) );
  INV_X1 U836 ( .A(n983), .ZN(G299) );
  BUF_X1 U837 ( .A(n761), .Z(G164) );
  NAND2_X1 U838 ( .A1(G94), .A2(G452), .ZN(n762) );
  XOR2_X1 U839 ( .A(KEYINPUT72), .B(n762), .Z(G173) );
  NAND2_X1 U840 ( .A1(G7), .A2(G661), .ZN(n763) );
  XOR2_X1 U841 ( .A(n763), .B(KEYINPUT10), .Z(n919) );
  NAND2_X1 U842 ( .A1(n919), .A2(G567), .ZN(n764) );
  XOR2_X1 U843 ( .A(KEYINPUT11), .B(n764), .Z(G234) );
  INV_X1 U844 ( .A(G860), .ZN(n772) );
  OR2_X1 U845 ( .A1(n982), .A2(n772), .ZN(G153) );
  INV_X1 U846 ( .A(G171), .ZN(G301) );
  INV_X1 U847 ( .A(G868), .ZN(n768) );
  AND2_X1 U848 ( .A1(n768), .A2(n972), .ZN(n766) );
  NOR2_X1 U849 ( .A1(n768), .A2(G301), .ZN(n765) );
  NOR2_X1 U850 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U851 ( .A(KEYINPUT76), .B(n767), .ZN(G284) );
  NOR2_X1 U852 ( .A1(G286), .A2(n768), .ZN(n769) );
  XNOR2_X1 U853 ( .A(n769), .B(KEYINPUT78), .ZN(n771) );
  NOR2_X1 U854 ( .A1(G299), .A2(G868), .ZN(n770) );
  NOR2_X1 U855 ( .A1(n771), .A2(n770), .ZN(G297) );
  NAND2_X1 U856 ( .A1(n772), .A2(G559), .ZN(n773) );
  NAND2_X1 U857 ( .A1(n773), .A2(n972), .ZN(n774) );
  XNOR2_X1 U858 ( .A(n774), .B(KEYINPUT16), .ZN(n776) );
  XOR2_X1 U859 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n775) );
  XNOR2_X1 U860 ( .A(n776), .B(n775), .ZN(G148) );
  NOR2_X1 U861 ( .A1(G868), .A2(n982), .ZN(n779) );
  NAND2_X1 U862 ( .A1(n972), .A2(G868), .ZN(n777) );
  NOR2_X1 U863 ( .A1(G559), .A2(n777), .ZN(n778) );
  NOR2_X1 U864 ( .A1(n779), .A2(n778), .ZN(G282) );
  NAND2_X1 U865 ( .A1(n899), .A2(G123), .ZN(n780) );
  XNOR2_X1 U866 ( .A(n780), .B(KEYINPUT18), .ZN(n782) );
  NAND2_X1 U867 ( .A1(G111), .A2(n710), .ZN(n781) );
  NAND2_X1 U868 ( .A1(n782), .A2(n781), .ZN(n786) );
  NAND2_X1 U869 ( .A1(G135), .A2(n894), .ZN(n784) );
  NAND2_X1 U870 ( .A1(G99), .A2(n895), .ZN(n783) );
  NAND2_X1 U871 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U872 ( .A1(n786), .A2(n785), .ZN(n928) );
  XOR2_X1 U873 ( .A(G2096), .B(n928), .Z(n787) );
  NOR2_X1 U874 ( .A1(G2100), .A2(n787), .ZN(n788) );
  XNOR2_X1 U875 ( .A(KEYINPUT81), .B(n788), .ZN(G156) );
  NAND2_X1 U876 ( .A1(n972), .A2(G559), .ZN(n814) );
  XNOR2_X1 U877 ( .A(n982), .B(n814), .ZN(n789) );
  NOR2_X1 U878 ( .A1(n789), .A2(G860), .ZN(n802) );
  NAND2_X1 U879 ( .A1(G67), .A2(n790), .ZN(n793) );
  NAND2_X1 U880 ( .A1(G55), .A2(n791), .ZN(n792) );
  NAND2_X1 U881 ( .A1(n793), .A2(n792), .ZN(n801) );
  NAND2_X1 U882 ( .A1(n794), .A2(G80), .ZN(n795) );
  XNOR2_X1 U883 ( .A(n795), .B(KEYINPUT82), .ZN(n798) );
  NAND2_X1 U884 ( .A1(G93), .A2(n796), .ZN(n797) );
  NAND2_X1 U885 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U886 ( .A(KEYINPUT83), .B(n799), .Z(n800) );
  NOR2_X1 U887 ( .A1(n801), .A2(n800), .ZN(n812) );
  XNOR2_X1 U888 ( .A(n802), .B(n812), .ZN(G145) );
  NOR2_X1 U889 ( .A1(G868), .A2(n812), .ZN(n803) );
  XNOR2_X1 U890 ( .A(n803), .B(KEYINPUT87), .ZN(n817) );
  XNOR2_X1 U891 ( .A(KEYINPUT85), .B(KEYINPUT19), .ZN(n805) );
  XNOR2_X1 U892 ( .A(G305), .B(KEYINPUT84), .ZN(n804) );
  XNOR2_X1 U893 ( .A(n805), .B(n804), .ZN(n808) );
  XOR2_X1 U894 ( .A(G299), .B(n982), .Z(n806) );
  XNOR2_X1 U895 ( .A(n806), .B(G288), .ZN(n807) );
  XNOR2_X1 U896 ( .A(n808), .B(n807), .ZN(n810) );
  XOR2_X1 U897 ( .A(G290), .B(G303), .Z(n809) );
  XNOR2_X1 U898 ( .A(n810), .B(n809), .ZN(n811) );
  XNOR2_X1 U899 ( .A(n812), .B(n811), .ZN(n910) );
  XOR2_X1 U900 ( .A(KEYINPUT86), .B(n910), .Z(n813) );
  XNOR2_X1 U901 ( .A(n814), .B(n813), .ZN(n815) );
  NAND2_X1 U902 ( .A1(G868), .A2(n815), .ZN(n816) );
  NAND2_X1 U903 ( .A1(n817), .A2(n816), .ZN(G295) );
  NAND2_X1 U904 ( .A1(G2078), .A2(G2084), .ZN(n818) );
  XOR2_X1 U905 ( .A(KEYINPUT20), .B(n818), .Z(n819) );
  NAND2_X1 U906 ( .A1(G2090), .A2(n819), .ZN(n821) );
  XNOR2_X1 U907 ( .A(KEYINPUT21), .B(KEYINPUT88), .ZN(n820) );
  XNOR2_X1 U908 ( .A(n821), .B(n820), .ZN(n822) );
  NAND2_X1 U909 ( .A1(G2072), .A2(n822), .ZN(G158) );
  XNOR2_X1 U910 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U911 ( .A1(G220), .A2(G219), .ZN(n823) );
  XOR2_X1 U912 ( .A(KEYINPUT22), .B(n823), .Z(n824) );
  NOR2_X1 U913 ( .A1(G218), .A2(n824), .ZN(n825) );
  NAND2_X1 U914 ( .A1(G96), .A2(n825), .ZN(n834) );
  NAND2_X1 U915 ( .A1(n834), .A2(G2106), .ZN(n829) );
  NAND2_X1 U916 ( .A1(G108), .A2(G120), .ZN(n826) );
  NOR2_X1 U917 ( .A1(G237), .A2(n826), .ZN(n827) );
  NAND2_X1 U918 ( .A1(G69), .A2(n827), .ZN(n835) );
  NAND2_X1 U919 ( .A1(n835), .A2(G567), .ZN(n828) );
  NAND2_X1 U920 ( .A1(n829), .A2(n828), .ZN(n918) );
  NAND2_X1 U921 ( .A1(G661), .A2(G483), .ZN(n830) );
  NOR2_X1 U922 ( .A1(n918), .A2(n830), .ZN(n833) );
  NAND2_X1 U923 ( .A1(n833), .A2(G36), .ZN(G176) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n919), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U926 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(G188) );
  XNOR2_X1 U929 ( .A(G120), .B(KEYINPUT111), .ZN(G236) );
  INV_X1 U931 ( .A(G108), .ZN(G238) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  NOR2_X1 U933 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  XOR2_X1 U935 ( .A(G2430), .B(G2451), .Z(n837) );
  XNOR2_X1 U936 ( .A(G2446), .B(G2427), .ZN(n836) );
  XNOR2_X1 U937 ( .A(n837), .B(n836), .ZN(n844) );
  XOR2_X1 U938 ( .A(G2438), .B(G2435), .Z(n839) );
  XNOR2_X1 U939 ( .A(G2443), .B(KEYINPUT109), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U941 ( .A(n840), .B(G2454), .Z(n842) );
  XNOR2_X1 U942 ( .A(G1348), .B(G1341), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n845) );
  NAND2_X1 U945 ( .A1(n845), .A2(G14), .ZN(n846) );
  XOR2_X1 U946 ( .A(KEYINPUT110), .B(n846), .Z(G401) );
  XOR2_X1 U947 ( .A(n847), .B(KEYINPUT41), .Z(n857) );
  XOR2_X1 U948 ( .A(G1976), .B(G1981), .Z(n849) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1971), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n971), .B(G1966), .ZN(n851) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U954 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U955 ( .A(KEYINPUT112), .B(G2474), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(G229) );
  XOR2_X1 U958 ( .A(G2100), .B(G2096), .Z(n859) );
  XNOR2_X1 U959 ( .A(KEYINPUT42), .B(G2678), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U961 ( .A(KEYINPUT43), .B(G2090), .Z(n861) );
  XNOR2_X1 U962 ( .A(G2067), .B(G2072), .ZN(n860) );
  XNOR2_X1 U963 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U964 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U965 ( .A(G2078), .B(G2084), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(G227) );
  NAND2_X1 U967 ( .A1(n899), .A2(G124), .ZN(n866) );
  XNOR2_X1 U968 ( .A(n866), .B(KEYINPUT44), .ZN(n868) );
  NAND2_X1 U969 ( .A1(G112), .A2(n710), .ZN(n867) );
  NAND2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G136), .A2(n894), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G100), .A2(n895), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U974 ( .A1(n872), .A2(n871), .ZN(G162) );
  XOR2_X1 U975 ( .A(G160), .B(n873), .Z(n876) );
  XNOR2_X1 U976 ( .A(n874), .B(G164), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n876), .B(n875), .ZN(n880) );
  XOR2_X1 U978 ( .A(n877), .B(G162), .Z(n878) );
  XNOR2_X1 U979 ( .A(n878), .B(n928), .ZN(n879) );
  XOR2_X1 U980 ( .A(n880), .B(n879), .Z(n885) );
  XOR2_X1 U981 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n882) );
  XNOR2_X1 U982 ( .A(KEYINPUT117), .B(KEYINPUT46), .ZN(n881) );
  XNOR2_X1 U983 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U984 ( .A(KEYINPUT48), .B(n883), .ZN(n884) );
  XNOR2_X1 U985 ( .A(n885), .B(n884), .ZN(n907) );
  NAND2_X1 U986 ( .A1(G139), .A2(n894), .ZN(n887) );
  NAND2_X1 U987 ( .A1(G103), .A2(n895), .ZN(n886) );
  NAND2_X1 U988 ( .A1(n887), .A2(n886), .ZN(n893) );
  NAND2_X1 U989 ( .A1(n899), .A2(G127), .ZN(n888) );
  XNOR2_X1 U990 ( .A(n888), .B(KEYINPUT116), .ZN(n890) );
  NAND2_X1 U991 ( .A1(G115), .A2(n710), .ZN(n889) );
  NAND2_X1 U992 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U993 ( .A(KEYINPUT47), .B(n891), .Z(n892) );
  NOR2_X1 U994 ( .A1(n893), .A2(n892), .ZN(n920) );
  NAND2_X1 U995 ( .A1(G142), .A2(n894), .ZN(n897) );
  NAND2_X1 U996 ( .A1(G106), .A2(n895), .ZN(n896) );
  NAND2_X1 U997 ( .A1(n897), .A2(n896), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n898), .B(KEYINPUT45), .ZN(n901) );
  NAND2_X1 U999 ( .A1(G130), .A2(n899), .ZN(n900) );
  NAND2_X1 U1000 ( .A1(n901), .A2(n900), .ZN(n904) );
  NAND2_X1 U1001 ( .A1(G118), .A2(n710), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(KEYINPUT113), .B(n902), .ZN(n903) );
  NOR2_X1 U1003 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n920), .B(n905), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n908), .ZN(G395) );
  XOR2_X1 U1007 ( .A(G301), .B(n972), .Z(n909) );
  XNOR2_X1 U1008 ( .A(n909), .B(G286), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n912), .ZN(G397) );
  OR2_X1 U1011 ( .A1(n918), .A2(G401), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(G229), .A2(G227), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1014 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(n918), .ZN(G319) );
  INV_X1 U1019 ( .A(G69), .ZN(G235) );
  INV_X1 U1020 ( .A(n919), .ZN(G223) );
  INV_X1 U1021 ( .A(G29), .ZN(n968) );
  XNOR2_X1 U1022 ( .A(G2072), .B(n920), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(G164), .B(G2078), .ZN(n921) );
  XNOR2_X1 U1024 ( .A(n921), .B(KEYINPUT118), .ZN(n922) );
  NAND2_X1 U1025 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1026 ( .A(n924), .B(KEYINPUT50), .ZN(n939) );
  XOR2_X1 U1027 ( .A(G2090), .B(G162), .Z(n925) );
  NOR2_X1 U1028 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1029 ( .A(KEYINPUT51), .B(n927), .Z(n937) );
  NOR2_X1 U1030 ( .A1(n929), .A2(n928), .ZN(n933) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n935) );
  XOR2_X1 U1033 ( .A(G160), .B(G2084), .Z(n934) );
  NOR2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n941) );
  NAND2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1039 ( .A(KEYINPUT52), .B(n944), .Z(n945) );
  NOR2_X1 U1040 ( .A1(KEYINPUT55), .A2(n945), .ZN(n946) );
  NOR2_X1 U1041 ( .A1(n968), .A2(n946), .ZN(n947) );
  XNOR2_X1 U1042 ( .A(n947), .B(KEYINPUT119), .ZN(n970) );
  XOR2_X1 U1043 ( .A(G2084), .B(G34), .Z(n948) );
  XNOR2_X1 U1044 ( .A(KEYINPUT54), .B(n948), .ZN(n964) );
  XNOR2_X1 U1045 ( .A(G2090), .B(G35), .ZN(n962) );
  XNOR2_X1 U1046 ( .A(G1991), .B(G25), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(G33), .B(G2072), .ZN(n949) );
  NOR2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n956) );
  XOR2_X1 U1049 ( .A(G32), .B(G1996), .Z(n951) );
  NAND2_X1 U1050 ( .A1(n951), .A2(G28), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(KEYINPUT120), .B(G2067), .ZN(n952) );
  XNOR2_X1 U1052 ( .A(G26), .B(n952), .ZN(n953) );
  NOR2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n959) );
  XOR2_X1 U1055 ( .A(G27), .B(n957), .Z(n958) );
  NOR2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1057 ( .A(KEYINPUT53), .B(n960), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(n965), .B(KEYINPUT121), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(KEYINPUT55), .B(n966), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n1027) );
  INV_X1 U1064 ( .A(G16), .ZN(n1022) );
  XOR2_X1 U1065 ( .A(n1022), .B(KEYINPUT56), .Z(n997) );
  XOR2_X1 U1066 ( .A(G171), .B(n971), .Z(n975) );
  XNOR2_X1 U1067 ( .A(G1348), .B(n972), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(n973), .B(KEYINPUT122), .ZN(n974) );
  NAND2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(n976), .B(KEYINPUT123), .ZN(n995) );
  XNOR2_X1 U1071 ( .A(G1966), .B(G168), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(n979), .B(KEYINPUT57), .ZN(n991) );
  NAND2_X1 U1074 ( .A1(G1971), .A2(G303), .ZN(n980) );
  NAND2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(n982), .B(G1341), .ZN(n985) );
  XOR2_X1 U1077 ( .A(n983), .B(G1956), .Z(n984) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1084 ( .A1(n997), .A2(n996), .ZN(n1024) );
  XOR2_X1 U1085 ( .A(G4), .B(KEYINPUT124), .Z(n999) );
  XNOR2_X1 U1086 ( .A(G1348), .B(KEYINPUT59), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(n999), .B(n998), .ZN(n1005) );
  XOR2_X1 U1088 ( .A(G20), .B(G1956), .Z(n1003) );
  XNOR2_X1 U1089 ( .A(G1341), .B(G19), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(G6), .B(G1981), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(KEYINPUT125), .B(KEYINPUT60), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(n1007), .B(n1006), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(G21), .B(G1966), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(KEYINPUT126), .B(n1010), .ZN(n1012) );
  XOR2_X1 U1099 ( .A(G1961), .B(G5), .Z(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1019) );
  XNOR2_X1 U1101 ( .A(G1971), .B(G22), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(G23), .B(G1976), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XOR2_X1 U1104 ( .A(G1986), .B(G24), .Z(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(KEYINPUT58), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1108 ( .A(KEYINPUT61), .B(n1020), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1111 ( .A(KEYINPUT127), .B(n1025), .Z(n1026) );
  NOR2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1113 ( .A1(n1028), .A2(G11), .ZN(n1029) );
  XNOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1029), .ZN(G150) );
  INV_X1 U1115 ( .A(G150), .ZN(G311) );
endmodule

