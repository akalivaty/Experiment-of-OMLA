

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(n709), .A2(n708), .ZN(n713) );
  NAND2_X1 U553 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U554 ( .A1(n720), .A2(n719), .ZN(n721) );
  OR2_X1 U555 ( .A1(n791), .A2(n696), .ZN(n697) );
  NOR2_X2 U556 ( .A1(n791), .A2(n696), .ZN(n707) );
  NOR2_X1 U557 ( .A1(n537), .A2(n536), .ZN(G160) );
  XOR2_X1 U558 ( .A(KEYINPUT29), .B(n723), .Z(n518) );
  OR2_X1 U559 ( .A1(n959), .A2(n762), .ZN(n519) );
  OR2_X1 U560 ( .A1(n770), .A2(n769), .ZN(n520) );
  NAND2_X1 U561 ( .A1(n702), .A2(n701), .ZN(n715) );
  NOR2_X1 U562 ( .A1(n715), .A2(n971), .ZN(n703) );
  XNOR2_X1 U563 ( .A(n748), .B(KEYINPUT98), .ZN(n749) );
  AND2_X1 U564 ( .A1(n771), .A2(n520), .ZN(n772) );
  NOR2_X2 U565 ( .A1(G2105), .A2(n525), .ZN(n881) );
  NOR2_X1 U566 ( .A1(G651), .A2(n647), .ZN(n660) );
  INV_X1 U567 ( .A(G2104), .ZN(n525) );
  INV_X1 U568 ( .A(G2105), .ZN(n521) );
  NOR2_X1 U569 ( .A1(n525), .A2(n521), .ZN(n886) );
  NAND2_X1 U570 ( .A1(G114), .A2(n886), .ZN(n523) );
  NOR2_X2 U571 ( .A1(G2104), .A2(n521), .ZN(n884) );
  NAND2_X1 U572 ( .A1(G126), .A2(n884), .ZN(n522) );
  NAND2_X1 U573 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U574 ( .A(KEYINPUT88), .B(n524), .ZN(n530) );
  NAND2_X1 U575 ( .A1(G102), .A2(n881), .ZN(n528) );
  NOR2_X1 U576 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XOR2_X2 U577 ( .A(KEYINPUT17), .B(n526), .Z(n879) );
  NAND2_X1 U578 ( .A1(G138), .A2(n879), .ZN(n527) );
  NAND2_X1 U579 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X2 U580 ( .A1(n530), .A2(n529), .ZN(G164) );
  NAND2_X1 U581 ( .A1(n886), .A2(G113), .ZN(n533) );
  NAND2_X1 U582 ( .A1(G101), .A2(n881), .ZN(n531) );
  XOR2_X1 U583 ( .A(KEYINPUT23), .B(n531), .Z(n532) );
  NAND2_X1 U584 ( .A1(n533), .A2(n532), .ZN(n537) );
  NAND2_X1 U585 ( .A1(G137), .A2(n879), .ZN(n535) );
  NAND2_X1 U586 ( .A1(G125), .A2(n884), .ZN(n534) );
  NAND2_X1 U587 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U588 ( .A(G2451), .B(G2454), .Z(n539) );
  XNOR2_X1 U589 ( .A(G2430), .B(KEYINPUT104), .ZN(n538) );
  XNOR2_X1 U590 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U591 ( .A(n540), .B(G2446), .Z(n542) );
  XNOR2_X1 U592 ( .A(G1341), .B(G1348), .ZN(n541) );
  XNOR2_X1 U593 ( .A(n542), .B(n541), .ZN(n546) );
  XOR2_X1 U594 ( .A(G2438), .B(G2427), .Z(n544) );
  XNOR2_X1 U595 ( .A(G2443), .B(G2435), .ZN(n543) );
  XNOR2_X1 U596 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U597 ( .A(n546), .B(n545), .Z(n547) );
  AND2_X1 U598 ( .A1(G14), .A2(n547), .ZN(G401) );
  INV_X1 U599 ( .A(G651), .ZN(n551) );
  NOR2_X1 U600 ( .A1(G543), .A2(n551), .ZN(n548) );
  XOR2_X1 U601 ( .A(KEYINPUT1), .B(n548), .Z(n656) );
  NAND2_X1 U602 ( .A1(G64), .A2(n656), .ZN(n550) );
  XOR2_X1 U603 ( .A(G543), .B(KEYINPUT0), .Z(n647) );
  NAND2_X1 U604 ( .A1(G52), .A2(n660), .ZN(n549) );
  NAND2_X1 U605 ( .A1(n550), .A2(n549), .ZN(n556) );
  NOR2_X1 U606 ( .A1(G651), .A2(G543), .ZN(n652) );
  NAND2_X1 U607 ( .A1(G90), .A2(n652), .ZN(n553) );
  NOR2_X1 U608 ( .A1(n647), .A2(n551), .ZN(n653) );
  NAND2_X1 U609 ( .A1(G77), .A2(n653), .ZN(n552) );
  NAND2_X1 U610 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U611 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  NOR2_X1 U612 ( .A1(n556), .A2(n555), .ZN(G171) );
  AND2_X1 U613 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U614 ( .A(G57), .ZN(G237) );
  INV_X1 U615 ( .A(G132), .ZN(G219) );
  INV_X1 U616 ( .A(G82), .ZN(G220) );
  NAND2_X1 U617 ( .A1(G7), .A2(G661), .ZN(n557) );
  XNOR2_X1 U618 ( .A(n557), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U619 ( .A(G223), .ZN(n827) );
  NAND2_X1 U620 ( .A1(n827), .A2(G567), .ZN(n558) );
  XOR2_X1 U621 ( .A(KEYINPUT11), .B(n558), .Z(G234) );
  XNOR2_X1 U622 ( .A(KEYINPUT67), .B(KEYINPUT13), .ZN(n563) );
  NAND2_X1 U623 ( .A1(n652), .A2(G81), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n559), .B(KEYINPUT12), .ZN(n561) );
  NAND2_X1 U625 ( .A1(G68), .A2(n653), .ZN(n560) );
  NAND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n563), .B(n562), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n656), .A2(G56), .ZN(n564) );
  XOR2_X1 U629 ( .A(KEYINPUT14), .B(n564), .Z(n565) );
  NOR2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n660), .A2(G43), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n974) );
  INV_X1 U633 ( .A(G860), .ZN(n626) );
  OR2_X1 U634 ( .A1(n974), .A2(n626), .ZN(G153) );
  INV_X1 U635 ( .A(G171), .ZN(G301) );
  NAND2_X1 U636 ( .A1(G301), .A2(G868), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n569), .B(KEYINPUT68), .ZN(n579) );
  INV_X1 U638 ( .A(G868), .ZN(n599) );
  NAND2_X1 U639 ( .A1(G66), .A2(n656), .ZN(n571) );
  NAND2_X1 U640 ( .A1(G54), .A2(n660), .ZN(n570) );
  NAND2_X1 U641 ( .A1(n571), .A2(n570), .ZN(n575) );
  NAND2_X1 U642 ( .A1(G92), .A2(n652), .ZN(n573) );
  NAND2_X1 U643 ( .A1(G79), .A2(n653), .ZN(n572) );
  NAND2_X1 U644 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U645 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U646 ( .A(KEYINPUT15), .B(n576), .Z(n577) );
  XNOR2_X1 U647 ( .A(KEYINPUT69), .B(n577), .ZN(n971) );
  NAND2_X1 U648 ( .A1(n599), .A2(n971), .ZN(n578) );
  NAND2_X1 U649 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U650 ( .A(KEYINPUT70), .B(n580), .ZN(G284) );
  NAND2_X1 U651 ( .A1(G63), .A2(n656), .ZN(n582) );
  NAND2_X1 U652 ( .A1(G51), .A2(n660), .ZN(n581) );
  NAND2_X1 U653 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U654 ( .A(KEYINPUT6), .B(n583), .ZN(n589) );
  NAND2_X1 U655 ( .A1(n652), .A2(G89), .ZN(n584) );
  XNOR2_X1 U656 ( .A(n584), .B(KEYINPUT4), .ZN(n586) );
  NAND2_X1 U657 ( .A1(G76), .A2(n653), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U659 ( .A(n587), .B(KEYINPUT5), .Z(n588) );
  NOR2_X1 U660 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U661 ( .A(KEYINPUT71), .B(n590), .Z(n591) );
  XOR2_X1 U662 ( .A(KEYINPUT7), .B(n591), .Z(G168) );
  XOR2_X1 U663 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U664 ( .A1(n656), .A2(G65), .ZN(n594) );
  NAND2_X1 U665 ( .A1(G78), .A2(n653), .ZN(n592) );
  XOR2_X1 U666 ( .A(KEYINPUT65), .B(n592), .Z(n593) );
  NAND2_X1 U667 ( .A1(n594), .A2(n593), .ZN(n598) );
  NAND2_X1 U668 ( .A1(G91), .A2(n652), .ZN(n596) );
  NAND2_X1 U669 ( .A1(G53), .A2(n660), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U671 ( .A1(n598), .A2(n597), .ZN(n964) );
  XOR2_X1 U672 ( .A(n964), .B(KEYINPUT66), .Z(G299) );
  NOR2_X1 U673 ( .A1(G286), .A2(n599), .ZN(n601) );
  NOR2_X1 U674 ( .A1(G299), .A2(G868), .ZN(n600) );
  NOR2_X1 U675 ( .A1(n601), .A2(n600), .ZN(G297) );
  NAND2_X1 U676 ( .A1(n626), .A2(G559), .ZN(n602) );
  INV_X1 U677 ( .A(n971), .ZN(n901) );
  NAND2_X1 U678 ( .A1(n602), .A2(n901), .ZN(n603) );
  XNOR2_X1 U679 ( .A(n603), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U680 ( .A1(G868), .A2(n974), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n901), .A2(G868), .ZN(n604) );
  NOR2_X1 U682 ( .A1(G559), .A2(n604), .ZN(n605) );
  NOR2_X1 U683 ( .A1(n606), .A2(n605), .ZN(G282) );
  NAND2_X1 U684 ( .A1(G123), .A2(n884), .ZN(n607) );
  XNOR2_X1 U685 ( .A(n607), .B(KEYINPUT18), .ZN(n608) );
  XNOR2_X1 U686 ( .A(KEYINPUT72), .B(n608), .ZN(n611) );
  NAND2_X1 U687 ( .A1(G111), .A2(n886), .ZN(n609) );
  XOR2_X1 U688 ( .A(KEYINPUT73), .B(n609), .Z(n610) );
  NAND2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U690 ( .A1(G99), .A2(n881), .ZN(n613) );
  NAND2_X1 U691 ( .A1(G135), .A2(n879), .ZN(n612) );
  NAND2_X1 U692 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n997) );
  XNOR2_X1 U694 ( .A(n997), .B(G2096), .ZN(n617) );
  INV_X1 U695 ( .A(G2100), .ZN(n616) );
  NAND2_X1 U696 ( .A1(n617), .A2(n616), .ZN(G156) );
  NAND2_X1 U697 ( .A1(G93), .A2(n652), .ZN(n619) );
  NAND2_X1 U698 ( .A1(G80), .A2(n653), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n624) );
  NAND2_X1 U700 ( .A1(G55), .A2(n660), .ZN(n620) );
  XNOR2_X1 U701 ( .A(n620), .B(KEYINPUT74), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n656), .A2(G67), .ZN(n621) );
  NAND2_X1 U703 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n664) );
  NAND2_X1 U705 ( .A1(G559), .A2(n901), .ZN(n625) );
  XOR2_X1 U706 ( .A(n974), .B(n625), .Z(n671) );
  NAND2_X1 U707 ( .A1(n626), .A2(n671), .ZN(n627) );
  XNOR2_X1 U708 ( .A(n627), .B(KEYINPUT75), .ZN(n628) );
  XNOR2_X1 U709 ( .A(n664), .B(n628), .ZN(G145) );
  NAND2_X1 U710 ( .A1(G60), .A2(n656), .ZN(n630) );
  NAND2_X1 U711 ( .A1(G47), .A2(n660), .ZN(n629) );
  NAND2_X1 U712 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U713 ( .A(KEYINPUT64), .B(n631), .Z(n635) );
  NAND2_X1 U714 ( .A1(G85), .A2(n652), .ZN(n633) );
  NAND2_X1 U715 ( .A1(G72), .A2(n653), .ZN(n632) );
  AND2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U717 ( .A1(n635), .A2(n634), .ZN(G290) );
  NAND2_X1 U718 ( .A1(G86), .A2(n652), .ZN(n637) );
  NAND2_X1 U719 ( .A1(G61), .A2(n656), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U721 ( .A(KEYINPUT78), .B(n638), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n653), .A2(G73), .ZN(n639) );
  XOR2_X1 U723 ( .A(KEYINPUT2), .B(n639), .Z(n640) );
  NOR2_X1 U724 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U725 ( .A1(n660), .A2(G48), .ZN(n642) );
  NAND2_X1 U726 ( .A1(n643), .A2(n642), .ZN(G305) );
  NAND2_X1 U727 ( .A1(G49), .A2(n660), .ZN(n645) );
  NAND2_X1 U728 ( .A1(G74), .A2(G651), .ZN(n644) );
  NAND2_X1 U729 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U730 ( .A(KEYINPUT76), .B(n646), .Z(n649) );
  NAND2_X1 U731 ( .A1(n647), .A2(G87), .ZN(n648) );
  NAND2_X1 U732 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U733 ( .A1(n650), .A2(n656), .ZN(n651) );
  XNOR2_X1 U734 ( .A(n651), .B(KEYINPUT77), .ZN(G288) );
  NAND2_X1 U735 ( .A1(G88), .A2(n652), .ZN(n655) );
  NAND2_X1 U736 ( .A1(G75), .A2(n653), .ZN(n654) );
  NAND2_X1 U737 ( .A1(n655), .A2(n654), .ZN(n659) );
  NAND2_X1 U738 ( .A1(G62), .A2(n656), .ZN(n657) );
  XNOR2_X1 U739 ( .A(KEYINPUT79), .B(n657), .ZN(n658) );
  NOR2_X1 U740 ( .A1(n659), .A2(n658), .ZN(n662) );
  NAND2_X1 U741 ( .A1(n660), .A2(G50), .ZN(n661) );
  NAND2_X1 U742 ( .A1(n662), .A2(n661), .ZN(G303) );
  INV_X1 U743 ( .A(G303), .ZN(G166) );
  NOR2_X1 U744 ( .A1(G868), .A2(n664), .ZN(n663) );
  XNOR2_X1 U745 ( .A(n663), .B(KEYINPUT81), .ZN(n674) );
  XNOR2_X1 U746 ( .A(n664), .B(G305), .ZN(n665) );
  XNOR2_X1 U747 ( .A(n665), .B(G288), .ZN(n666) );
  XOR2_X1 U748 ( .A(n666), .B(KEYINPUT80), .Z(n668) );
  XNOR2_X1 U749 ( .A(G166), .B(KEYINPUT19), .ZN(n667) );
  XNOR2_X1 U750 ( .A(n668), .B(n667), .ZN(n669) );
  XOR2_X1 U751 ( .A(G299), .B(n669), .Z(n670) );
  XNOR2_X1 U752 ( .A(G290), .B(n670), .ZN(n900) );
  XNOR2_X1 U753 ( .A(n900), .B(n671), .ZN(n672) );
  NAND2_X1 U754 ( .A1(G868), .A2(n672), .ZN(n673) );
  NAND2_X1 U755 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U756 ( .A1(G2078), .A2(G2084), .ZN(n676) );
  XOR2_X1 U757 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n675) );
  XNOR2_X1 U758 ( .A(n676), .B(n675), .ZN(n677) );
  NAND2_X1 U759 ( .A1(G2090), .A2(n677), .ZN(n678) );
  XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n678), .ZN(n679) );
  NAND2_X1 U761 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U763 ( .A1(G220), .A2(G219), .ZN(n680) );
  XOR2_X1 U764 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U765 ( .A1(G218), .A2(n681), .ZN(n682) );
  XOR2_X1 U766 ( .A(KEYINPUT83), .B(n682), .Z(n683) );
  NAND2_X1 U767 ( .A1(G96), .A2(n683), .ZN(n832) );
  NAND2_X1 U768 ( .A1(G2106), .A2(n832), .ZN(n684) );
  XNOR2_X1 U769 ( .A(n684), .B(KEYINPUT84), .ZN(n688) );
  NAND2_X1 U770 ( .A1(G69), .A2(G120), .ZN(n685) );
  NOR2_X1 U771 ( .A1(G237), .A2(n685), .ZN(n686) );
  NAND2_X1 U772 ( .A1(G108), .A2(n686), .ZN(n831) );
  NAND2_X1 U773 ( .A1(G567), .A2(n831), .ZN(n687) );
  NAND2_X1 U774 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U775 ( .A(KEYINPUT85), .B(n689), .ZN(G319) );
  NAND2_X1 U776 ( .A1(G661), .A2(G483), .ZN(n690) );
  XOR2_X1 U777 ( .A(KEYINPUT86), .B(n690), .Z(n691) );
  NAND2_X1 U778 ( .A1(n691), .A2(G319), .ZN(n692) );
  XNOR2_X1 U779 ( .A(n692), .B(KEYINPUT87), .ZN(n830) );
  NAND2_X1 U780 ( .A1(n830), .A2(G36), .ZN(G176) );
  XNOR2_X1 U781 ( .A(G1981), .B(G305), .ZN(n959) );
  XOR2_X1 U782 ( .A(G2078), .B(KEYINPUT25), .Z(n938) );
  NAND2_X1 U783 ( .A1(G160), .A2(G40), .ZN(n791) );
  NOR2_X2 U784 ( .A1(G164), .A2(G1384), .ZN(n792) );
  INV_X1 U785 ( .A(n792), .ZN(n696) );
  INV_X1 U786 ( .A(n707), .ZN(n734) );
  NOR2_X1 U787 ( .A1(n938), .A2(n734), .ZN(n693) );
  XNOR2_X1 U788 ( .A(n693), .B(KEYINPUT95), .ZN(n695) );
  INV_X1 U789 ( .A(G1961), .ZN(n912) );
  NAND2_X1 U790 ( .A1(n912), .A2(n734), .ZN(n694) );
  NAND2_X1 U791 ( .A1(n695), .A2(n694), .ZN(n728) );
  NAND2_X1 U792 ( .A1(n728), .A2(G171), .ZN(n724) );
  NAND2_X1 U793 ( .A1(n697), .A2(G1341), .ZN(n698) );
  XOR2_X1 U794 ( .A(KEYINPUT96), .B(n698), .Z(n699) );
  NOR2_X1 U795 ( .A1(n974), .A2(n699), .ZN(n702) );
  NAND2_X1 U796 ( .A1(n707), .A2(G1996), .ZN(n700) );
  XNOR2_X1 U797 ( .A(KEYINPUT26), .B(n700), .ZN(n701) );
  XNOR2_X1 U798 ( .A(n703), .B(KEYINPUT97), .ZN(n712) );
  NOR2_X1 U799 ( .A1(G2067), .A2(n734), .ZN(n705) );
  NOR2_X1 U800 ( .A1(n707), .A2(G1348), .ZN(n704) );
  NOR2_X1 U801 ( .A1(n705), .A2(n704), .ZN(n710) );
  NAND2_X1 U802 ( .A1(n707), .A2(G2072), .ZN(n706) );
  XNOR2_X1 U803 ( .A(n706), .B(KEYINPUT27), .ZN(n709) );
  INV_X1 U804 ( .A(G1956), .ZN(n913) );
  NOR2_X1 U805 ( .A1(n913), .A2(n707), .ZN(n708) );
  NAND2_X1 U806 ( .A1(n964), .A2(n713), .ZN(n716) );
  AND2_X1 U807 ( .A1(n710), .A2(n716), .ZN(n711) );
  NAND2_X1 U808 ( .A1(n712), .A2(n711), .ZN(n722) );
  NOR2_X1 U809 ( .A1(n964), .A2(n713), .ZN(n714) );
  XOR2_X1 U810 ( .A(n714), .B(KEYINPUT28), .Z(n720) );
  NAND2_X1 U811 ( .A1(n715), .A2(n971), .ZN(n718) );
  INV_X1 U812 ( .A(n716), .ZN(n717) );
  OR2_X1 U813 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U814 ( .A1(n724), .A2(n518), .ZN(n733) );
  NAND2_X1 U815 ( .A1(n734), .A2(G8), .ZN(n769) );
  NOR2_X1 U816 ( .A1(G1966), .A2(n769), .ZN(n742) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n734), .ZN(n745) );
  NOR2_X1 U818 ( .A1(n742), .A2(n745), .ZN(n725) );
  NAND2_X1 U819 ( .A1(G8), .A2(n725), .ZN(n726) );
  XNOR2_X1 U820 ( .A(KEYINPUT30), .B(n726), .ZN(n727) );
  NOR2_X1 U821 ( .A1(G168), .A2(n727), .ZN(n730) );
  NOR2_X1 U822 ( .A1(G171), .A2(n728), .ZN(n729) );
  NOR2_X1 U823 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U824 ( .A(KEYINPUT31), .B(n731), .Z(n732) );
  NAND2_X1 U825 ( .A1(n733), .A2(n732), .ZN(n743) );
  NAND2_X1 U826 ( .A1(G286), .A2(n743), .ZN(n739) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n769), .ZN(n736) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n734), .ZN(n735) );
  NOR2_X1 U829 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U830 ( .A1(n737), .A2(G303), .ZN(n738) );
  NAND2_X1 U831 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U832 ( .A1(n740), .A2(G8), .ZN(n741) );
  XNOR2_X1 U833 ( .A(KEYINPUT32), .B(n741), .ZN(n750) );
  INV_X1 U834 ( .A(n742), .ZN(n744) );
  AND2_X1 U835 ( .A1(n744), .A2(n743), .ZN(n747) );
  NAND2_X1 U836 ( .A1(G8), .A2(n745), .ZN(n746) );
  NAND2_X1 U837 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U838 ( .A1(n750), .A2(n749), .ZN(n765) );
  NOR2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n757) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n751) );
  NOR2_X1 U841 ( .A1(n757), .A2(n751), .ZN(n965) );
  NAND2_X1 U842 ( .A1(n765), .A2(n965), .ZN(n753) );
  NAND2_X1 U843 ( .A1(G288), .A2(G1976), .ZN(n752) );
  XOR2_X1 U844 ( .A(KEYINPUT99), .B(n752), .Z(n977) );
  NAND2_X1 U845 ( .A1(n753), .A2(n977), .ZN(n754) );
  NOR2_X1 U846 ( .A1(KEYINPUT33), .A2(n754), .ZN(n755) );
  INV_X1 U847 ( .A(n769), .ZN(n756) );
  NAND2_X1 U848 ( .A1(n755), .A2(n756), .ZN(n760) );
  NAND2_X1 U849 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U850 ( .A1(n758), .A2(KEYINPUT33), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U852 ( .A(KEYINPUT100), .B(n761), .Z(n762) );
  NOR2_X1 U853 ( .A1(G2090), .A2(G303), .ZN(n763) );
  NAND2_X1 U854 ( .A1(G8), .A2(n763), .ZN(n764) );
  NAND2_X1 U855 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U856 ( .A1(n769), .A2(n766), .ZN(n771) );
  NOR2_X1 U857 ( .A1(G1981), .A2(G305), .ZN(n767) );
  XOR2_X1 U858 ( .A(n767), .B(KEYINPUT24), .Z(n768) );
  XNOR2_X1 U859 ( .A(KEYINPUT94), .B(n768), .ZN(n770) );
  NAND2_X1 U860 ( .A1(n519), .A2(n772), .ZN(n807) );
  NAND2_X1 U861 ( .A1(G107), .A2(n886), .ZN(n774) );
  NAND2_X1 U862 ( .A1(G119), .A2(n884), .ZN(n773) );
  NAND2_X1 U863 ( .A1(n774), .A2(n773), .ZN(n778) );
  NAND2_X1 U864 ( .A1(G95), .A2(n881), .ZN(n776) );
  NAND2_X1 U865 ( .A1(G131), .A2(n879), .ZN(n775) );
  NAND2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n777) );
  OR2_X1 U867 ( .A1(n778), .A2(n777), .ZN(n876) );
  NAND2_X1 U868 ( .A1(G1991), .A2(n876), .ZN(n779) );
  XNOR2_X1 U869 ( .A(n779), .B(KEYINPUT91), .ZN(n790) );
  NAND2_X1 U870 ( .A1(G129), .A2(n884), .ZN(n780) );
  XNOR2_X1 U871 ( .A(n780), .B(KEYINPUT92), .ZN(n784) );
  XOR2_X1 U872 ( .A(KEYINPUT93), .B(KEYINPUT38), .Z(n782) );
  NAND2_X1 U873 ( .A1(G105), .A2(n881), .ZN(n781) );
  XNOR2_X1 U874 ( .A(n782), .B(n781), .ZN(n783) );
  NAND2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n788) );
  NAND2_X1 U876 ( .A1(G117), .A2(n886), .ZN(n786) );
  NAND2_X1 U877 ( .A1(G141), .A2(n879), .ZN(n785) );
  NAND2_X1 U878 ( .A1(n786), .A2(n785), .ZN(n787) );
  OR2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n894) );
  AND2_X1 U880 ( .A1(G1996), .A2(n894), .ZN(n789) );
  NOR2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n988) );
  XOR2_X1 U882 ( .A(G1986), .B(G290), .Z(n973) );
  NAND2_X1 U883 ( .A1(n988), .A2(n973), .ZN(n793) );
  NOR2_X1 U884 ( .A1(n792), .A2(n791), .ZN(n818) );
  NAND2_X1 U885 ( .A1(n793), .A2(n818), .ZN(n805) );
  XNOR2_X1 U886 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n798) );
  NAND2_X1 U887 ( .A1(G116), .A2(n886), .ZN(n795) );
  NAND2_X1 U888 ( .A1(G128), .A2(n884), .ZN(n794) );
  NAND2_X1 U889 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U890 ( .A(n796), .B(KEYINPUT35), .ZN(n797) );
  XNOR2_X1 U891 ( .A(n798), .B(n797), .ZN(n803) );
  NAND2_X1 U892 ( .A1(G104), .A2(n881), .ZN(n800) );
  NAND2_X1 U893 ( .A1(G140), .A2(n879), .ZN(n799) );
  NAND2_X1 U894 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U895 ( .A(KEYINPUT34), .B(n801), .ZN(n802) );
  NOR2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n804) );
  XOR2_X1 U897 ( .A(KEYINPUT36), .B(n804), .Z(n897) );
  XOR2_X1 U898 ( .A(G2067), .B(KEYINPUT37), .Z(n808) );
  AND2_X1 U899 ( .A1(n897), .A2(n808), .ZN(n986) );
  NAND2_X1 U900 ( .A1(n986), .A2(n818), .ZN(n809) );
  AND2_X1 U901 ( .A1(n805), .A2(n809), .ZN(n806) );
  NAND2_X1 U902 ( .A1(n807), .A2(n806), .ZN(n825) );
  NOR2_X1 U903 ( .A1(n897), .A2(n808), .ZN(n985) );
  NAND2_X1 U904 ( .A1(n985), .A2(n818), .ZN(n823) );
  INV_X1 U905 ( .A(n809), .ZN(n821) );
  NOR2_X1 U906 ( .A1(G1996), .A2(n894), .ZN(n990) );
  INV_X1 U907 ( .A(n988), .ZN(n814) );
  NOR2_X1 U908 ( .A1(G1986), .A2(G290), .ZN(n811) );
  NOR2_X1 U909 ( .A1(G1991), .A2(n876), .ZN(n810) );
  XOR2_X1 U910 ( .A(KEYINPUT101), .B(n810), .Z(n998) );
  NOR2_X1 U911 ( .A1(n811), .A2(n998), .ZN(n812) );
  XNOR2_X1 U912 ( .A(n812), .B(KEYINPUT102), .ZN(n813) );
  NOR2_X1 U913 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U914 ( .A1(n990), .A2(n815), .ZN(n816) );
  XOR2_X1 U915 ( .A(KEYINPUT39), .B(n816), .Z(n817) );
  XNOR2_X1 U916 ( .A(KEYINPUT103), .B(n817), .ZN(n819) );
  NAND2_X1 U917 ( .A1(n819), .A2(n818), .ZN(n820) );
  OR2_X1 U918 ( .A1(n821), .A2(n820), .ZN(n822) );
  AND2_X1 U919 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U921 ( .A(n826), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n827), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U924 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U926 ( .A1(n830), .A2(n829), .ZN(G188) );
  XNOR2_X1 U927 ( .A(G96), .B(KEYINPUT105), .ZN(G221) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G69), .ZN(G235) );
  NOR2_X1 U931 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U932 ( .A(n833), .B(KEYINPUT106), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  XOR2_X1 U934 ( .A(KEYINPUT41), .B(G1981), .Z(n835) );
  XNOR2_X1 U935 ( .A(G1966), .B(G1956), .ZN(n834) );
  XNOR2_X1 U936 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U937 ( .A(n836), .B(KEYINPUT108), .Z(n838) );
  XNOR2_X1 U938 ( .A(G1996), .B(G1991), .ZN(n837) );
  XNOR2_X1 U939 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U940 ( .A(G1986), .B(G1976), .Z(n840) );
  XNOR2_X1 U941 ( .A(G1961), .B(G1971), .ZN(n839) );
  XNOR2_X1 U942 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U943 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U944 ( .A(KEYINPUT107), .B(G2474), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(G229) );
  XOR2_X1 U946 ( .A(G2100), .B(G2096), .Z(n846) );
  XNOR2_X1 U947 ( .A(KEYINPUT42), .B(G2678), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U949 ( .A(KEYINPUT43), .B(G2090), .Z(n848) );
  XNOR2_X1 U950 ( .A(G2072), .B(G2067), .ZN(n847) );
  XNOR2_X1 U951 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U952 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2084), .ZN(n851) );
  XNOR2_X1 U954 ( .A(n852), .B(n851), .ZN(G227) );
  NAND2_X1 U955 ( .A1(G100), .A2(n881), .ZN(n854) );
  NAND2_X1 U956 ( .A1(G112), .A2(n886), .ZN(n853) );
  NAND2_X1 U957 ( .A1(n854), .A2(n853), .ZN(n860) );
  NAND2_X1 U958 ( .A1(n884), .A2(G124), .ZN(n855) );
  XNOR2_X1 U959 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U960 ( .A1(G136), .A2(n879), .ZN(n856) );
  NAND2_X1 U961 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U962 ( .A(KEYINPUT109), .B(n858), .Z(n859) );
  NOR2_X1 U963 ( .A1(n860), .A2(n859), .ZN(G162) );
  XOR2_X1 U964 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n862) );
  XNOR2_X1 U965 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n861) );
  XNOR2_X1 U966 ( .A(n862), .B(n861), .ZN(n865) );
  XNOR2_X1 U967 ( .A(G160), .B(n997), .ZN(n863) );
  XNOR2_X1 U968 ( .A(n863), .B(G162), .ZN(n864) );
  XNOR2_X1 U969 ( .A(n865), .B(n864), .ZN(n878) );
  NAND2_X1 U970 ( .A1(G118), .A2(n886), .ZN(n867) );
  NAND2_X1 U971 ( .A1(G130), .A2(n884), .ZN(n866) );
  NAND2_X1 U972 ( .A1(n867), .A2(n866), .ZN(n874) );
  NAND2_X1 U973 ( .A1(n879), .A2(G142), .ZN(n868) );
  XNOR2_X1 U974 ( .A(n868), .B(KEYINPUT110), .ZN(n870) );
  NAND2_X1 U975 ( .A1(G106), .A2(n881), .ZN(n869) );
  NAND2_X1 U976 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U977 ( .A(KEYINPUT45), .B(n871), .ZN(n872) );
  XNOR2_X1 U978 ( .A(KEYINPUT111), .B(n872), .ZN(n873) );
  NOR2_X1 U979 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U980 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U981 ( .A(n878), .B(n877), .ZN(n893) );
  NAND2_X1 U982 ( .A1(n879), .A2(G139), .ZN(n880) );
  XNOR2_X1 U983 ( .A(n880), .B(KEYINPUT112), .ZN(n883) );
  NAND2_X1 U984 ( .A1(G103), .A2(n881), .ZN(n882) );
  NAND2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n892) );
  NAND2_X1 U986 ( .A1(n884), .A2(G127), .ZN(n885) );
  XOR2_X1 U987 ( .A(KEYINPUT113), .B(n885), .Z(n888) );
  NAND2_X1 U988 ( .A1(n886), .A2(G115), .ZN(n887) );
  NAND2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U990 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  XNOR2_X1 U991 ( .A(KEYINPUT114), .B(n890), .ZN(n891) );
  NOR2_X1 U992 ( .A1(n892), .A2(n891), .ZN(n992) );
  XOR2_X1 U993 ( .A(n893), .B(n992), .Z(n896) );
  XOR2_X1 U994 ( .A(G164), .B(n894), .Z(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n898) );
  XOR2_X1 U996 ( .A(n898), .B(n897), .Z(n899) );
  NOR2_X1 U997 ( .A1(G37), .A2(n899), .ZN(G395) );
  XOR2_X1 U998 ( .A(KEYINPUT117), .B(n900), .Z(n903) );
  XNOR2_X1 U999 ( .A(n901), .B(G286), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(n974), .B(G171), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n906), .ZN(G397) );
  NOR2_X1 U1004 ( .A1(G229), .A2(G227), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n907), .ZN(n908) );
  NOR2_X1 U1006 ( .A1(G401), .A2(n908), .ZN(n909) );
  AND2_X1 U1007 ( .A1(G319), .A2(n909), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n910) );
  NAND2_X1 U1009 ( .A1(n911), .A2(n910), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1012 ( .A(n912), .B(G5), .ZN(n933) );
  XOR2_X1 U1013 ( .A(G1966), .B(G21), .Z(n924) );
  XNOR2_X1 U1014 ( .A(G20), .B(n913), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(G1341), .B(G19), .ZN(n915) );
  XNOR2_X1 U1016 ( .A(G6), .B(G1981), .ZN(n914) );
  NOR2_X1 U1017 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1018 ( .A(KEYINPUT125), .B(n916), .Z(n917) );
  NAND2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n921) );
  XOR2_X1 U1020 ( .A(KEYINPUT59), .B(G1348), .Z(n919) );
  XNOR2_X1 U1021 ( .A(G4), .B(n919), .ZN(n920) );
  NOR2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1023 ( .A(KEYINPUT60), .B(n922), .ZN(n923) );
  NAND2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n931) );
  XNOR2_X1 U1025 ( .A(G1971), .B(G22), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(G23), .B(G1976), .ZN(n925) );
  NOR2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n928) );
  XOR2_X1 U1028 ( .A(G1986), .B(G24), .Z(n927) );
  NAND2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(KEYINPUT58), .B(n929), .ZN(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(n934), .B(KEYINPUT126), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(n935), .B(KEYINPUT61), .ZN(n936) );
  NOR2_X1 U1035 ( .A1(G16), .A2(n936), .ZN(n937) );
  XNOR2_X1 U1036 ( .A(n937), .B(KEYINPUT127), .ZN(n957) );
  XNOR2_X1 U1037 ( .A(G2090), .B(G35), .ZN(n952) );
  XOR2_X1 U1038 ( .A(n938), .B(G27), .Z(n940) );
  XOR2_X1 U1039 ( .A(G1996), .B(G32), .Z(n939) );
  NAND2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(G26), .B(G2067), .ZN(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n945) );
  XOR2_X1 U1043 ( .A(G2072), .B(KEYINPUT122), .Z(n943) );
  XNOR2_X1 U1044 ( .A(G33), .B(n943), .ZN(n944) );
  NAND2_X1 U1045 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1046 ( .A(KEYINPUT123), .B(n946), .ZN(n947) );
  NAND2_X1 U1047 ( .A1(n947), .A2(G28), .ZN(n949) );
  XNOR2_X1 U1048 ( .A(G25), .B(G1991), .ZN(n948) );
  NOR2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1050 ( .A(KEYINPUT53), .B(n950), .ZN(n951) );
  NOR2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n955) );
  XOR2_X1 U1052 ( .A(G2084), .B(G34), .Z(n953) );
  XNOR2_X1 U1053 ( .A(KEYINPUT54), .B(n953), .ZN(n954) );
  NAND2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n1017) );
  XOR2_X1 U1055 ( .A(KEYINPUT55), .B(KEYINPUT121), .Z(n1015) );
  INV_X1 U1056 ( .A(n1015), .ZN(n1010) );
  OR2_X1 U1057 ( .A1(n1017), .A2(n1010), .ZN(n956) );
  NAND2_X1 U1058 ( .A1(n957), .A2(n956), .ZN(n984) );
  XOR2_X1 U1059 ( .A(G16), .B(KEYINPUT56), .Z(n982) );
  XOR2_X1 U1060 ( .A(G168), .B(G1966), .Z(n958) );
  NOR2_X1 U1061 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1062 ( .A(KEYINPUT124), .B(n960), .Z(n961) );
  XNOR2_X1 U1063 ( .A(KEYINPUT57), .B(n961), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(G171), .B(G1961), .ZN(n963) );
  NAND2_X1 U1065 ( .A1(G1971), .A2(G303), .ZN(n962) );
  NAND2_X1 U1066 ( .A1(n963), .A2(n962), .ZN(n968) );
  XNOR2_X1 U1067 ( .A(n964), .B(G1956), .ZN(n966) );
  NAND2_X1 U1068 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1069 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1070 ( .A1(n970), .A2(n969), .ZN(n980) );
  XOR2_X1 U1071 ( .A(G1348), .B(n971), .Z(n972) );
  NAND2_X1 U1072 ( .A1(n973), .A2(n972), .ZN(n976) );
  XNOR2_X1 U1073 ( .A(G1341), .B(n974), .ZN(n975) );
  NOR2_X1 U1074 ( .A1(n976), .A2(n975), .ZN(n978) );
  NAND2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n1014) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n1008) );
  XOR2_X1 U1081 ( .A(G2090), .B(G162), .Z(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1083 ( .A(KEYINPUT51), .B(n991), .Z(n1006) );
  XOR2_X1 U1084 ( .A(G164), .B(G2078), .Z(n995) );
  XOR2_X1 U1085 ( .A(n992), .B(KEYINPUT120), .Z(n993) );
  XNOR2_X1 U1086 ( .A(G2072), .B(n993), .ZN(n994) );
  NOR2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1088 ( .A(KEYINPUT50), .B(n996), .Z(n1004) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1090 ( .A(KEYINPUT118), .B(n999), .Z(n1001) );
  XOR2_X1 U1091 ( .A(G160), .B(G2084), .Z(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(KEYINPUT119), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(KEYINPUT52), .B(n1009), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(G29), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1020) );
  NOR2_X1 U1101 ( .A1(G29), .A2(n1015), .ZN(n1016) );
  NAND2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1103 ( .A1(G11), .A2(n1018), .ZN(n1019) );
  NOR2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1105 ( .A(n1021), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

