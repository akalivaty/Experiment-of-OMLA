//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT64), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n463), .A3(G137), .ZN(new_n464));
  NAND2_X1  g039(.A1(G101), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n468), .B1(new_n469), .B2(G125), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT65), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n461), .A2(new_n463), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(new_n467), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n474), .A2(new_n475), .A3(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n466), .B1(new_n472), .B2(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n469), .A2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n469), .A2(new_n471), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n480), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND3_X1  g062(.A1(new_n461), .A2(new_n463), .A3(G126), .ZN(new_n488));
  NAND2_X1  g063(.A1(G114), .A2(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT66), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n471), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n490), .A2(G2105), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(G102), .A2(G2104), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT66), .A2(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n493), .A2(G138), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n461), .A2(new_n463), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(new_n471), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(KEYINPUT67), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT67), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .A3(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(new_n512), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n510), .A2(G88), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n506), .B1(new_n515), .B2(new_n516), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G50), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT68), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n518), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n521), .B1(new_n518), .B2(new_n520), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n513), .B1(new_n522), .B2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND2_X1  g100(.A1(new_n519), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n510), .A2(new_n517), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n526), .B(new_n528), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n510), .A2(KEYINPUT69), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n510), .A2(KEYINPUT69), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n534), .A2(G63), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n531), .B1(new_n535), .B2(G651), .ZN(G168));
  NAND2_X1  g111(.A1(new_n519), .A2(G52), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n529), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n534), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n541), .B2(new_n512), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  AOI22_X1  g118(.A1(new_n534), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n512), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n519), .A2(G43), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n529), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(new_n519), .A2(G53), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n519), .A2(KEYINPUT9), .A3(G53), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g135(.A1(G78), .A2(G543), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n510), .B2(G65), .ZN(new_n562));
  INV_X1    g137(.A(G91), .ZN(new_n563));
  OAI22_X1  g138(.A1(new_n562), .A2(new_n512), .B1(new_n529), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT70), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G299));
  INV_X1    g142(.A(G168), .ZN(G286));
  OAI21_X1  g143(.A(G651), .B1(new_n534), .B2(G74), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n510), .A2(new_n517), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n570), .A2(G87), .B1(G49), .B2(new_n519), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT71), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT71), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n569), .A2(new_n574), .A3(new_n571), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(G288));
  NAND3_X1  g151(.A1(new_n510), .A2(G86), .A3(new_n517), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT72), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT73), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n519), .A2(new_n579), .A3(G48), .ZN(new_n580));
  INV_X1    g155(.A(new_n516), .ZN(new_n581));
  NOR2_X1   g156(.A1(KEYINPUT6), .A2(G651), .ZN(new_n582));
  OAI211_X1 g157(.A(G48), .B(G543), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(KEYINPUT73), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n512), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n578), .A2(new_n585), .A3(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n570), .A2(G85), .B1(G47), .B2(new_n519), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n534), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n591), .B2(new_n512), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n519), .A2(G54), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n510), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(new_n512), .ZN(new_n596));
  XOR2_X1   g171(.A(new_n596), .B(KEYINPUT74), .Z(new_n597));
  NAND2_X1  g172(.A1(new_n570), .A2(G92), .ZN(new_n598));
  XOR2_X1   g173(.A(new_n598), .B(KEYINPUT10), .Z(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n593), .B1(new_n601), .B2(G868), .ZN(G321));
  XNOR2_X1  g177(.A(G321), .B(KEYINPUT75), .ZN(G284));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(new_n566), .B2(G868), .ZN(G297));
  OAI21_X1  g180(.A(new_n604), .B1(new_n566), .B2(G868), .ZN(G280));
  NOR2_X1   g181(.A1(new_n600), .A2(G559), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n607), .B1(G860), .B2(new_n601), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT76), .Z(G148));
  INV_X1    g184(.A(new_n549), .ZN(new_n610));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n607), .B2(new_n611), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR3_X1    g189(.A1(new_n481), .A2(KEYINPUT12), .A3(new_n460), .ZN(new_n615));
  OAI21_X1  g190(.A(KEYINPUT12), .B1(new_n481), .B2(new_n460), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2100), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n479), .A2(G123), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n482), .A2(G135), .ZN(new_n621));
  NOR2_X1   g196(.A1(G99), .A2(G2105), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(new_n471), .B2(G111), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n620), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  NAND2_X1  g200(.A1(new_n619), .A2(new_n625), .ZN(G156));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2435), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2438), .ZN(new_n628));
  XOR2_X1   g203(.A(G2427), .B(G2430), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT78), .B(KEYINPUT14), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2451), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n632), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n638), .B(new_n639), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G14), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(G401));
  XNOR2_X1  g217(.A(G2084), .B(G2090), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT79), .ZN(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n644), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT18), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n645), .B(KEYINPUT17), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(KEYINPUT80), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(new_n644), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n645), .ZN(new_n653));
  INV_X1    g228(.A(new_n644), .ZN(new_n654));
  OAI211_X1 g229(.A(new_n653), .B(new_n654), .C1(new_n650), .C2(new_n651), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n649), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2096), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2100), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G227));
  XOR2_X1   g234(.A(G1956), .B(G2474), .Z(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n660), .A2(new_n661), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT20), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n666), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n663), .A2(new_n665), .A3(new_n667), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n670), .B(new_n671), .C1(new_n669), .C2(new_n668), .ZN(new_n672));
  XOR2_X1   g247(.A(G1981), .B(G1986), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1991), .B(G1996), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT81), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n676), .B(new_n678), .Z(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G229));
  NAND2_X1  g255(.A1(G168), .A2(G16), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n681), .B(KEYINPUT88), .C1(G16), .C2(G21), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(KEYINPUT88), .B2(new_n681), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT89), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G1966), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT90), .B(KEYINPUT31), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G11), .ZN(new_n687));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G20), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT95), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT23), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(new_n566), .B2(new_n688), .ZN(new_n692));
  INV_X1    g267(.A(G1956), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n685), .A2(new_n687), .A3(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G1961), .ZN(new_n696));
  NOR2_X1   g271(.A1(G171), .A2(new_n688), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n688), .A2(G5), .ZN(new_n698));
  OR3_X1    g273(.A1(new_n697), .A2(KEYINPUT92), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(KEYINPUT92), .B1(new_n697), .B2(new_n698), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n696), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(G29), .A2(G32), .ZN(new_n702));
  AOI22_X1  g277(.A1(new_n469), .A2(G141), .B1(G105), .B2(G2104), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n703), .A2(G2105), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G129), .B2(new_n479), .ZN(new_n705));
  NAND3_X1  g280(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT26), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n702), .B1(new_n710), .B2(G29), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT27), .B(G1996), .Z(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n624), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT91), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT30), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(G28), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(G28), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n718), .A2(new_n719), .A3(new_n714), .ZN(new_n720));
  OR2_X1    g295(.A1(G29), .A2(G33), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n482), .A2(G139), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT25), .Z(new_n724));
  AOI22_X1  g299(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT86), .Z(new_n726));
  OAI211_X1 g301(.A(new_n722), .B(new_n724), .C1(new_n726), .C2(new_n471), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n721), .B1(new_n727), .B2(new_n714), .ZN(new_n728));
  INV_X1    g303(.A(G2072), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n720), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR4_X1   g305(.A1(new_n701), .A2(new_n713), .A3(new_n716), .A4(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n728), .A2(new_n729), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  NOR3_X1   g309(.A1(new_n695), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n714), .A2(G35), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G162), .B2(new_n714), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT94), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT29), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(G2090), .ZN(new_n740));
  INV_X1    g315(.A(new_n684), .ZN(new_n741));
  INV_X1    g316(.A(G1966), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT24), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n714), .B1(new_n744), .B2(G34), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT87), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n744), .A2(G34), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n745), .A2(new_n746), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G160), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(new_n714), .ZN(new_n752));
  INV_X1    g327(.A(G2084), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n739), .A2(G2090), .ZN(new_n755));
  AND3_X1   g330(.A1(new_n743), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n699), .A2(new_n696), .A3(new_n700), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n711), .A2(new_n712), .B1(new_n753), .B2(new_n752), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT93), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n714), .A2(G27), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G164), .B2(new_n714), .ZN(new_n762));
  INV_X1    g337(.A(G2078), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n735), .A2(new_n756), .A3(new_n760), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(G16), .A2(G23), .ZN(new_n766));
  INV_X1    g341(.A(new_n572), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT33), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1976), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n688), .A2(G22), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G166), .B2(new_n688), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT83), .B(G1971), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  MUX2_X1   g349(.A(G6), .B(G305), .S(G16), .Z(new_n775));
  XOR2_X1   g350(.A(KEYINPUT32), .B(G1981), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n770), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT82), .B(KEYINPUT34), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n778), .A2(new_n780), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(G290), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n784), .A2(new_n688), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n688), .B2(G24), .ZN(new_n786));
  INV_X1    g361(.A(G1986), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n479), .A2(G119), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n482), .A2(G131), .ZN(new_n791));
  NOR2_X1   g366(.A1(G95), .A2(G2105), .ZN(new_n792));
  OAI21_X1  g367(.A(G2104), .B1(new_n471), .B2(G107), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n790), .B(new_n791), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  MUX2_X1   g369(.A(G25), .B(new_n794), .S(G29), .Z(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT35), .B(G1991), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n795), .B(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n788), .A2(new_n789), .A3(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n783), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(KEYINPUT36), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT36), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n783), .A2(new_n803), .A3(new_n800), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n765), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n688), .A2(G4), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n601), .B2(new_n688), .ZN(new_n807));
  INV_X1    g382(.A(G1348), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n688), .A2(G19), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n549), .B2(new_n688), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G1341), .Z(new_n812));
  XOR2_X1   g387(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n714), .A2(G26), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n479), .A2(G128), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n482), .A2(G140), .ZN(new_n817));
  OR2_X1    g392(.A1(G104), .A2(G2105), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n818), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n815), .B1(new_n821), .B2(new_n714), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT85), .B(G2067), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n805), .A2(new_n809), .A3(new_n812), .A4(new_n824), .ZN(G150));
  NAND2_X1  g400(.A1(G150), .A2(KEYINPUT96), .ZN(new_n826));
  INV_X1    g401(.A(new_n695), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n827), .A2(new_n764), .A3(new_n733), .A4(new_n731), .ZN(new_n828));
  INV_X1    g403(.A(new_n760), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n743), .A2(new_n754), .A3(new_n755), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n803), .B1(new_n783), .B2(new_n800), .ZN(new_n832));
  AOI211_X1 g407(.A(KEYINPUT36), .B(new_n799), .C1(new_n781), .C2(new_n782), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n831), .B(new_n824), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT96), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n835), .A2(new_n836), .A3(new_n809), .A4(new_n812), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n826), .A2(new_n837), .ZN(G311));
  NAND2_X1  g413(.A1(new_n534), .A2(G67), .ZN(new_n839));
  NAND2_X1  g414(.A1(G80), .A2(G543), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n839), .A2(KEYINPUT97), .A3(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT97), .ZN(new_n842));
  INV_X1    g417(.A(G67), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n532), .B2(new_n533), .ZN(new_n844));
  INV_X1    g419(.A(new_n840), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n841), .A2(G651), .A3(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT98), .B(G93), .ZN(new_n848));
  AOI22_X1  g423(.A1(new_n570), .A2(new_n848), .B1(G55), .B2(new_n519), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT100), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n847), .A2(new_n852), .A3(new_n849), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(G860), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n601), .A2(G559), .ZN(new_n858));
  XNOR2_X1  g433(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n850), .A2(new_n549), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n853), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n852), .B1(new_n847), .B2(new_n849), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n610), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n850), .A2(new_n549), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(KEYINPUT99), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n863), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n860), .B(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n857), .B1(new_n870), .B2(G860), .ZN(G145));
  INV_X1    g446(.A(G142), .ZN(new_n872));
  NOR2_X1   g447(.A1(G106), .A2(G2105), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(new_n471), .B2(G118), .ZN(new_n874));
  OAI22_X1  g449(.A1(new_n481), .A2(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(G130), .B2(new_n479), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n617), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n794), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT102), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n820), .B(new_n503), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n710), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n727), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n878), .A2(KEYINPUT102), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n883), .B1(new_n884), .B2(new_n882), .ZN(new_n885));
  XNOR2_X1  g460(.A(G160), .B(new_n624), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n486), .B(KEYINPUT101), .Z(new_n888));
  OR2_X1    g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(G37), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n888), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(KEYINPUT103), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n889), .A2(new_n894), .A3(new_n890), .A4(new_n891), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT40), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n893), .A2(new_n895), .A3(KEYINPUT40), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(G395));
  NAND2_X1  g475(.A1(new_n855), .A2(new_n611), .ZN(new_n901));
  XNOR2_X1  g476(.A(G299), .B(new_n600), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(KEYINPUT41), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n600), .B(new_n566), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT104), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n903), .B(new_n906), .Z(new_n907));
  XOR2_X1   g482(.A(new_n869), .B(new_n607), .Z(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n902), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n909), .B1(new_n910), .B2(KEYINPUT105), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(KEYINPUT105), .B2(new_n909), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n572), .B(G303), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(new_n784), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(G305), .ZN(new_n915));
  XOR2_X1   g490(.A(new_n915), .B(KEYINPUT42), .Z(new_n916));
  XNOR2_X1  g491(.A(new_n912), .B(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n901), .B1(new_n917), .B2(new_n611), .ZN(G295));
  OAI21_X1  g493(.A(new_n901), .B1(new_n917), .B2(new_n611), .ZN(G331));
  NOR2_X1   g494(.A1(new_n869), .A2(G171), .ZN(new_n920));
  AOI22_X1  g495(.A1(new_n854), .A2(new_n610), .B1(new_n861), .B2(new_n862), .ZN(new_n921));
  AOI21_X1  g496(.A(G301), .B1(new_n921), .B2(new_n868), .ZN(new_n922));
  OAI21_X1  g497(.A(G286), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n869), .A2(G171), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(G301), .A3(new_n868), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n925), .A3(G168), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(new_n926), .A3(new_n904), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT106), .ZN(new_n928));
  INV_X1    g503(.A(new_n915), .ZN(new_n929));
  INV_X1    g504(.A(new_n926), .ZN(new_n930));
  AOI21_X1  g505(.A(G168), .B1(new_n924), .B2(new_n925), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n907), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n923), .A2(new_n926), .A3(new_n933), .A4(new_n904), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n928), .A2(new_n929), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n935), .A2(new_n890), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n928), .A2(new_n932), .A3(new_n934), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n915), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT43), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n927), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n904), .A2(new_n905), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(KEYINPUT107), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n923), .A2(new_n926), .B1(new_n903), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n915), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  AND4_X1   g519(.A1(KEYINPUT43), .A2(new_n935), .A3(new_n890), .A4(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT44), .B1(new_n939), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n948), .B1(new_n936), .B2(new_n938), .ZN(new_n949));
  AND4_X1   g524(.A1(new_n948), .A2(new_n935), .A3(new_n890), .A4(new_n944), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n946), .A2(new_n951), .ZN(G397));
  INV_X1    g527(.A(G8), .ZN(new_n953));
  INV_X1    g528(.A(G1384), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n495), .A2(new_n494), .ZN(new_n955));
  INV_X1    g530(.A(new_n489), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n956), .B1(new_n469), .B2(G126), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n955), .B1(new_n957), .B2(new_n471), .ZN(new_n958));
  INV_X1    g533(.A(G138), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(KEYINPUT66), .B2(KEYINPUT4), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n469), .A2(new_n493), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(G2105), .B1(new_n961), .B2(new_n497), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n954), .B1(new_n958), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT112), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n503), .A2(new_n965), .A3(new_n954), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g542(.A(KEYINPUT108), .B(G40), .Z(new_n968));
  AOI211_X1 g543(.A(new_n466), .B(new_n968), .C1(new_n472), .C2(new_n476), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n953), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G1981), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n578), .A2(new_n588), .A3(new_n971), .A4(new_n585), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT49), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n585), .A2(KEYINPUT115), .A3(new_n577), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT115), .B1(new_n585), .B2(new_n577), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n975), .A2(new_n976), .A3(new_n587), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n972), .B(new_n973), .C1(new_n977), .C2(new_n971), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n976), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n980), .A2(new_n588), .A3(new_n974), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(G1981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n973), .B1(new_n982), .B2(new_n972), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n970), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n767), .A2(G1976), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n970), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT52), .ZN(new_n987));
  INV_X1    g562(.A(G1976), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT52), .B1(G288), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n989), .A2(new_n970), .A3(new_n985), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n984), .A2(new_n987), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT50), .B1(new_n964), .B2(new_n966), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n993));
  AOI21_X1  g568(.A(G1384), .B1(new_n496), .B2(new_n502), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n969), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n992), .A2(new_n995), .A3(G2090), .ZN(new_n996));
  INV_X1    g571(.A(new_n466), .ZN(new_n997));
  INV_X1    g572(.A(new_n968), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n475), .B1(new_n474), .B2(G2105), .ZN(new_n999));
  AOI211_X1 g574(.A(KEYINPUT65), .B(new_n471), .C1(new_n473), .C2(new_n467), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n997), .B(new_n998), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1001), .B1(KEYINPUT45), .B2(new_n994), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n963), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1971), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(G8), .B1(new_n996), .B2(new_n1005), .ZN(new_n1006));
  NOR4_X1   g581(.A1(G166), .A2(KEYINPUT113), .A3(KEYINPUT55), .A4(new_n953), .ZN(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1009), .B1(G303), .B2(G8), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT114), .B1(new_n1006), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1005), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n965), .B1(new_n503), .B2(new_n954), .ZN(new_n1015));
  AOI211_X1 g590(.A(KEYINPUT112), .B(G1384), .C1(new_n496), .C2(new_n502), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n993), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G2090), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1001), .B1(KEYINPUT50), .B2(new_n963), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n953), .B1(new_n1014), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n1022), .A3(new_n1011), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n991), .B1(new_n1013), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n964), .A2(KEYINPUT50), .A3(new_n966), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n994), .A2(new_n993), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n969), .A3(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(G2090), .ZN(new_n1028));
  OAI21_X1  g603(.A(G8), .B1(new_n1028), .B2(new_n1005), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n1012), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1024), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n964), .A2(new_n1003), .A3(new_n966), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n1002), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n742), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1017), .A2(new_n753), .A3(new_n1019), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(G168), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(G168), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT51), .ZN(new_n1038));
  OAI211_X1 g613(.A(G8), .B(new_n1036), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n992), .A2(new_n995), .A3(G2084), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1966), .B1(new_n1032), .B2(new_n1002), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1040), .A2(new_n1041), .A3(G286), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT51), .B1(new_n1042), .B2(new_n953), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(G301), .B(KEYINPUT54), .ZN(new_n1045));
  OAI211_X1 g620(.A(KEYINPUT45), .B(new_n954), .C1(new_n958), .C2(new_n962), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1004), .A2(KEYINPUT53), .A3(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n466), .B(KEYINPUT123), .ZN(new_n1048));
  INV_X1    g623(.A(G40), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n470), .A2(new_n471), .ZN(new_n1050));
  NOR4_X1   g625(.A1(new_n1048), .A2(new_n1049), .A3(G2078), .A4(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1045), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n696), .B1(new_n992), .B2(new_n995), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1002), .A2(new_n763), .A3(new_n1004), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(KEYINPUT122), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT122), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1052), .A2(new_n1053), .A3(new_n1056), .A4(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1032), .A2(new_n763), .A3(new_n1002), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT53), .B1(new_n1061), .B2(KEYINPUT121), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(KEYINPUT121), .B2(new_n1061), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1059), .A2(new_n1053), .A3(new_n1056), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1045), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1044), .A2(new_n1060), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1027), .A2(new_n693), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT56), .B(G2072), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1002), .A2(new_n1004), .A3(new_n1068), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n510), .A2(G65), .ZN(new_n1071));
  OAI21_X1  g646(.A(G651), .B1(new_n1071), .B2(new_n561), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n570), .A2(G91), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1072), .A2(new_n558), .A3(new_n559), .A4(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT118), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n565), .A2(new_n1077), .A3(KEYINPUT57), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n559), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT9), .B1(new_n519), .B2(G53), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT116), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n558), .A2(new_n1083), .A3(new_n559), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1082), .A2(new_n1084), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1085), .A2(new_n1086), .A3(new_n1075), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1086), .B1(new_n1085), .B2(new_n1075), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1079), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n1070), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1067), .A2(new_n1089), .A3(new_n1069), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n808), .B1(new_n992), .B2(new_n995), .ZN(new_n1092));
  INV_X1    g667(.A(G2067), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n967), .A2(new_n1093), .A3(new_n969), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1095), .A2(KEYINPUT119), .A3(new_n601), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT119), .B1(new_n1095), .B2(new_n601), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1091), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1091), .A2(KEYINPUT61), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT61), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1067), .A2(new_n1089), .A3(new_n1100), .A4(new_n1069), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n969), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT58), .B(G1341), .Z(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G1996), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1004), .A2(new_n969), .A3(new_n1105), .A4(new_n1046), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT120), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1002), .A2(new_n1108), .A3(new_n1105), .A4(new_n1004), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1104), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1110), .A2(new_n1111), .A3(new_n549), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1111), .B1(new_n1110), .B2(new_n549), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1099), .B(new_n1101), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT60), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n601), .B1(new_n1095), .B2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1092), .A2(new_n1094), .A3(KEYINPUT60), .A4(new_n600), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1116), .A2(new_n1117), .B1(new_n1115), .B2(new_n1095), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1090), .B(new_n1098), .C1(new_n1114), .C2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1066), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT63), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1121), .B1(new_n1006), .B2(new_n1012), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1024), .A2(new_n1122), .ZN(new_n1123));
  AOI211_X1 g698(.A(new_n953), .B(G286), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1031), .B1(new_n1120), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1013), .A2(new_n1023), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1127), .A2(new_n991), .ZN(new_n1128));
  INV_X1    g703(.A(new_n991), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1127), .A2(new_n1129), .A3(new_n1122), .A4(new_n1124), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1128), .B1(new_n1130), .B2(KEYINPUT63), .ZN(new_n1131));
  INV_X1    g706(.A(new_n970), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n979), .A2(new_n983), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1133), .A2(new_n988), .A3(new_n573), .A4(new_n575), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1132), .B1(new_n1134), .B2(new_n972), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1131), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT124), .B1(new_n1126), .B2(new_n1137), .ZN(new_n1138));
  AOI211_X1 g713(.A(new_n1135), .B(new_n1128), .C1(new_n1130), .C2(KEYINPUT63), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1119), .A2(new_n1066), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1139), .B(new_n1140), .C1(new_n1141), .C2(new_n1031), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1044), .A2(KEYINPUT62), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1144), .A2(G301), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1143), .A2(new_n1024), .A3(new_n1030), .A4(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT125), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1044), .A2(KEYINPUT62), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1031), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1150), .A2(KEYINPUT125), .A3(new_n1145), .A4(new_n1143), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1148), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1138), .A2(new_n1142), .A3(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1004), .A2(new_n1001), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n820), .B(new_n1093), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT110), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n709), .B(G1996), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1154), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT111), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1154), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n794), .B(new_n797), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n784), .A2(new_n1154), .A3(new_n787), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1154), .A2(G1986), .A3(G290), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT109), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1162), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1153), .A2(new_n1167), .ZN(new_n1168));
  XOR2_X1   g743(.A(new_n1163), .B(KEYINPUT48), .Z(new_n1169));
  NOR2_X1   g744(.A1(new_n1162), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n794), .A2(new_n796), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1159), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n821), .A2(new_n1093), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1160), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1154), .B1(new_n1156), .B2(new_n709), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT46), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1176), .B1(new_n1160), .B2(G1996), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1154), .A2(KEYINPUT46), .A3(new_n1105), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1175), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1179), .B(KEYINPUT47), .Z(new_n1180));
  NOR3_X1   g755(.A1(new_n1170), .A2(new_n1174), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1168), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1168), .A2(KEYINPUT126), .A3(new_n1181), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g761(.A1(new_n641), .A2(G319), .A3(new_n658), .ZN(new_n1188));
  XNOR2_X1  g762(.A(new_n1188), .B(KEYINPUT127), .ZN(new_n1189));
  NAND2_X1  g763(.A1(new_n892), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g764(.A(new_n938), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n935), .A2(new_n890), .ZN(new_n1192));
  OAI21_X1  g766(.A(KEYINPUT43), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g767(.A1(new_n936), .A2(new_n948), .A3(new_n944), .ZN(new_n1194));
  AOI211_X1 g768(.A(G229), .B(new_n1190), .C1(new_n1193), .C2(new_n1194), .ZN(G308));
  AOI21_X1  g769(.A(G229), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1196));
  NAND3_X1  g770(.A1(new_n1196), .A2(new_n892), .A3(new_n1189), .ZN(G225));
endmodule


