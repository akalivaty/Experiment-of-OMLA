//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT64), .ZN(new_n458));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n459), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n458), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(KEYINPUT64), .A3(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n462), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G101), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n473), .B1(new_n465), .B2(G2105), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n461), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g051(.A(KEYINPUT65), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(new_n463), .A3(G2104), .ZN(new_n479));
  AND4_X1   g054(.A1(new_n461), .A2(new_n477), .A3(new_n479), .A4(new_n466), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n476), .B1(new_n480), .B2(G137), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n471), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n477), .A2(new_n479), .A3(G2105), .A4(new_n466), .ZN(new_n486));
  INV_X1    g061(.A(G124), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(G136), .B2(new_n480), .ZN(G162));
  AND3_X1   g064(.A1(new_n477), .A2(new_n479), .A3(new_n466), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n490), .A2(KEYINPUT67), .A3(G126), .A4(G2105), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n492));
  INV_X1    g067(.A(G126), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n486), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n477), .A2(new_n479), .A3(new_n461), .A4(new_n466), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT4), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n497), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n459), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n495), .A2(new_n501), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT68), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT68), .A3(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n508), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n520), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n511), .A2(new_n513), .B1(KEYINPUT5), .B2(new_n510), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n523), .A2(new_n520), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT69), .B(G88), .Z(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n519), .A2(new_n522), .A3(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n520), .A2(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT71), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT71), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n520), .A2(new_n532), .A3(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n524), .A2(G89), .ZN(new_n536));
  XNOR2_X1  g111(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n537), .B(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n535), .A2(new_n536), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT70), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n542), .B(new_n543), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n529), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n542), .B(KEYINPUT70), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n539), .B1(new_n534), .B2(G51), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n546), .A2(new_n547), .A3(KEYINPUT73), .A4(new_n536), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n545), .A2(new_n548), .ZN(G168));
  NAND2_X1  g124(.A1(new_n534), .A2(G52), .ZN(new_n550));
  INV_X1    g125(.A(G90), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n523), .A2(new_n520), .ZN(new_n552));
  NAND2_X1  g127(.A1(G77), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G64), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n516), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n555), .A2(new_n556), .ZN(new_n559));
  OAI221_X1 g134(.A(new_n550), .B1(new_n551), .B2(new_n552), .C1(new_n558), .C2(new_n559), .ZN(G301));
  INV_X1    g135(.A(G301), .ZN(G171));
  AOI22_X1  g136(.A1(new_n534), .A2(G43), .B1(new_n524), .B2(G81), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G651), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  INV_X1    g147(.A(KEYINPUT9), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n521), .A2(new_n573), .A3(G53), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT9), .B1(new_n530), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(G91), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n578), .B2(new_n552), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n514), .A2(G65), .A3(new_n515), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT75), .ZN(new_n582));
  NAND2_X1  g157(.A1(G78), .A2(G543), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G651), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n582), .B1(new_n581), .B2(new_n583), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n580), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n581), .A2(new_n583), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT75), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n589), .A2(KEYINPUT76), .A3(G651), .A4(new_n584), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n579), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G299));
  INV_X1    g167(.A(G168), .ZN(G286));
  NAND2_X1  g168(.A1(new_n524), .A2(G87), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n521), .A2(G49), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G288));
  NAND4_X1  g172(.A1(new_n514), .A2(G86), .A3(new_n515), .A4(new_n520), .ZN(new_n598));
  INV_X1    g173(.A(G48), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n523), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n600));
  OAI221_X1 g175(.A(new_n598), .B1(new_n599), .B2(new_n530), .C1(new_n600), .C2(new_n564), .ZN(G305));
  AOI22_X1  g176(.A1(new_n534), .A2(G47), .B1(new_n524), .B2(G85), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n564), .B2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  AND3_X1   g180(.A1(new_n523), .A2(G92), .A3(new_n520), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(KEYINPUT10), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n523), .A2(G66), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G651), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n534), .A2(G54), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n610), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n564), .B1(new_n611), .B2(new_n612), .ZN(new_n617));
  INV_X1    g192(.A(G54), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n618), .B1(new_n531), .B2(new_n533), .ZN(new_n619));
  NOR3_X1   g194(.A1(new_n617), .A2(new_n619), .A3(KEYINPUT77), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n609), .B1(new_n616), .B2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n605), .B1(new_n622), .B2(G868), .ZN(G284));
  OAI21_X1  g198(.A(new_n605), .B1(new_n622), .B2(G868), .ZN(G321));
  NOR2_X1   g199(.A1(G299), .A2(G868), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n625), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g201(.A(new_n625), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n622), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n622), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G868), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(G868), .B2(new_n567), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g208(.A(new_n474), .ZN(new_n634));
  INV_X1    g209(.A(new_n475), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n459), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2100), .ZN(new_n639));
  OR2_X1    g214(.A1(G99), .A2(G2105), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n640), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n641));
  INV_X1    g216(.A(G123), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n641), .B1(new_n486), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(G135), .B2(new_n480), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n639), .A2(new_n645), .ZN(G156));
  INV_X1    g221(.A(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2427), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n647), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(new_n650), .B2(new_n649), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n652), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  AND3_X1   g235(.A1(new_n659), .A2(G14), .A3(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT17), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n663), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT78), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n663), .A2(new_n664), .ZN(new_n669));
  INV_X1    g244(.A(new_n662), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n669), .B(new_n666), .C1(new_n670), .C2(new_n664), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(new_n664), .A3(new_n665), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT18), .Z(new_n673));
  NAND3_X1  g248(.A1(new_n668), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2096), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT79), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1956), .B(G2474), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT20), .Z(new_n685));
  NOR2_X1   g260(.A1(new_n678), .A2(new_n680), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n687), .A2(new_n683), .A3(new_n681), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n685), .B(new_n688), .C1(new_n683), .C2(new_n687), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n693), .B(new_n694), .Z(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  NOR2_X1   g271(.A1(G6), .A2(G16), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n600), .A2(new_n564), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n598), .B1(new_n599), .B2(new_n530), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n697), .B1(new_n700), .B2(G16), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT32), .ZN(new_n702));
  INV_X1    g277(.A(G1981), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G22), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G166), .B2(new_n705), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT82), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n708), .A2(G1971), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(G1971), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n705), .A2(G23), .ZN(new_n711));
  INV_X1    g286(.A(G288), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(new_n705), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT33), .B(G1976), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  AND4_X1   g290(.A1(new_n704), .A2(new_n709), .A3(new_n710), .A4(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT34), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  MUX2_X1   g294(.A(G24), .B(G290), .S(G16), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G1986), .ZN(new_n721));
  OR2_X1    g296(.A1(G25), .A2(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n480), .A2(G131), .ZN(new_n723));
  INV_X1    g298(.A(G95), .ZN(new_n724));
  AND3_X1   g299(.A1(new_n724), .A2(new_n461), .A3(KEYINPUT80), .ZN(new_n725));
  AOI21_X1  g300(.A(KEYINPUT80), .B1(new_n724), .B2(new_n461), .ZN(new_n726));
  OAI221_X1 g301(.A(G2104), .B1(G107), .B2(new_n461), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G119), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n723), .B(new_n727), .C1(new_n728), .C2(new_n486), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT81), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(KEYINPUT81), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n722), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT35), .B(G1991), .Z(new_n736));
  AND2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NOR3_X1   g313(.A1(new_n721), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n718), .A2(new_n719), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT36), .ZN(new_n741));
  NOR2_X1   g316(.A1(G171), .A2(new_n705), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G5), .B2(new_n705), .ZN(new_n743));
  INV_X1    g318(.A(G1961), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(G164), .A2(G29), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G27), .B2(G29), .ZN(new_n747));
  INV_X1    g322(.A(G2078), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n734), .A2(G35), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G162), .B2(new_n734), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT29), .Z(new_n752));
  INV_X1    g327(.A(G2090), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n745), .A2(new_n749), .A3(new_n754), .ZN(new_n755));
  OAI22_X1  g330(.A1(new_n743), .A2(new_n744), .B1(new_n747), .B2(new_n748), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n705), .A2(G4), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n622), .B2(new_n705), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(G1348), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n734), .A2(G32), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n480), .A2(G141), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n490), .A2(G129), .A3(G2105), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT26), .Z(new_n764));
  OAI21_X1  g339(.A(G105), .B1(new_n634), .B2(new_n635), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n761), .A2(new_n762), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT89), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n760), .B1(new_n767), .B2(new_n734), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT27), .B(G1996), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n758), .A2(G1348), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n759), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(G16), .A2(G19), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n567), .B2(G16), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT83), .B(G1341), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT24), .ZN(new_n777));
  INV_X1    g352(.A(G34), .ZN(new_n778));
  AOI21_X1  g353(.A(G29), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n777), .B2(new_n778), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G160), .B2(new_n734), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G2084), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n734), .A2(G26), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(G104), .ZN(new_n786));
  AND3_X1   g361(.A1(new_n786), .A2(new_n461), .A3(KEYINPUT84), .ZN(new_n787));
  AOI21_X1  g362(.A(KEYINPUT84), .B1(new_n786), .B2(new_n461), .ZN(new_n788));
  OAI221_X1 g363(.A(G2104), .B1(G116), .B2(new_n461), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G128), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(new_n486), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n480), .A2(G140), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n785), .B1(new_n793), .B2(new_n734), .ZN(new_n794));
  INV_X1    g369(.A(G2067), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n644), .A2(G29), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT31), .B(G11), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT30), .B(G28), .Z(new_n799));
  OAI211_X1 g374(.A(new_n797), .B(new_n798), .C1(G29), .C2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n781), .ZN(new_n801));
  INV_X1    g376(.A(G2084), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n776), .A2(new_n782), .A3(new_n796), .A4(new_n803), .ZN(new_n804));
  NOR4_X1   g379(.A1(new_n755), .A2(new_n756), .A3(new_n772), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n752), .A2(new_n753), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT93), .ZN(new_n807));
  NOR2_X1   g382(.A1(G29), .A2(G33), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT25), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G139), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(new_n496), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT86), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n459), .A2(G127), .ZN(new_n817));
  INV_X1    g392(.A(G115), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n465), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n815), .A2(new_n816), .B1(G2105), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n808), .B1(new_n820), .B2(G29), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(G2072), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT87), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(G2072), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT88), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n807), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n805), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n705), .A2(G20), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT23), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n591), .B2(new_n705), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G1956), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n705), .A2(G21), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(G168), .B2(new_n705), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT90), .B(G1966), .Z(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT91), .Z(new_n837));
  NOR2_X1   g412(.A1(new_n833), .A2(new_n835), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT92), .ZN(new_n839));
  NOR4_X1   g414(.A1(new_n827), .A2(new_n831), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n741), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(G311));
  XNOR2_X1  g417(.A(new_n841), .B(KEYINPUT94), .ZN(G150));
  NOR2_X1   g418(.A1(new_n621), .A2(new_n628), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n534), .A2(G55), .B1(new_n524), .B2(G93), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n847), .A2(new_n564), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n566), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n562), .A2(new_n846), .A3(new_n565), .A4(new_n848), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n845), .B(new_n852), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n853), .A2(KEYINPUT39), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n853), .A2(KEYINPUT39), .ZN(new_n855));
  NOR3_X1   g430(.A1(new_n854), .A2(new_n855), .A3(G860), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n849), .A2(G860), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT37), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n856), .A2(new_n858), .ZN(G145));
  INV_X1    g434(.A(KEYINPUT96), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n820), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n506), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n793), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(new_n767), .ZN(new_n864));
  INV_X1    g439(.A(new_n793), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n862), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n767), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G130), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n461), .A2(G118), .ZN(new_n870));
  OAI21_X1  g445(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n871));
  OAI22_X1  g446(.A1(new_n486), .A2(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n872), .B1(G142), .B2(new_n480), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n637), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n733), .B(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n864), .A2(new_n868), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT97), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n864), .A2(new_n868), .ZN(new_n879));
  INV_X1    g454(.A(new_n875), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n878), .B(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n644), .B(KEYINPUT95), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(G162), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n482), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n885), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n876), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(G37), .B1(new_n888), .B2(new_n881), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n886), .A2(KEYINPUT40), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT40), .B1(new_n886), .B2(new_n889), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(G395));
  NOR2_X1   g467(.A1(new_n849), .A2(G868), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n630), .B(new_n852), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n621), .A2(new_n591), .A3(KEYINPUT98), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT98), .B1(new_n621), .B2(new_n591), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n621), .A2(new_n591), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n894), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT99), .ZN(new_n902));
  OAI21_X1  g477(.A(KEYINPUT100), .B1(new_n895), .B2(new_n896), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n621), .A2(new_n591), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT98), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT100), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n621), .A2(new_n591), .A3(KEYINPUT98), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n903), .A2(new_n909), .A3(new_n899), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n898), .A2(new_n911), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n910), .A2(new_n911), .B1(new_n897), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n902), .B1(new_n894), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT102), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(G290), .B(new_n700), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n712), .B(G303), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n921), .B(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(new_n914), .B2(new_n915), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n916), .B(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n893), .B1(new_n925), .B2(G868), .ZN(G295));
  AOI21_X1  g501(.A(new_n893), .B1(new_n925), .B2(G868), .ZN(G331));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n545), .A2(new_n928), .A3(new_n548), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(G301), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n928), .B1(new_n545), .B2(new_n548), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n931), .A2(new_n852), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n852), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n931), .A2(new_n852), .ZN(new_n935));
  INV_X1    g510(.A(new_n930), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n931), .A2(new_n852), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n934), .A2(new_n900), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n938), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  OAI211_X1 g516(.A(KEYINPUT104), .B(new_n939), .C1(new_n913), .C2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n910), .A2(new_n911), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n897), .A2(new_n912), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(new_n946), .A3(new_n940), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n942), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n921), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n921), .B(KEYINPUT105), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n942), .A2(new_n947), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G37), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n903), .A2(new_n909), .A3(new_n912), .ZN(new_n956));
  INV_X1    g531(.A(new_n900), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n956), .B1(new_n957), .B2(KEYINPUT41), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n940), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n941), .A2(KEYINPUT106), .A3(new_n900), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n939), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(G37), .B1(new_n963), .B2(new_n952), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n949), .A2(new_n964), .ZN(new_n965));
  OAI221_X1 g540(.A(KEYINPUT44), .B1(new_n951), .B2(new_n955), .C1(new_n965), .C2(new_n950), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n942), .A2(new_n947), .B1(new_n919), .B2(new_n920), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT43), .B1(new_n955), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n949), .A2(new_n964), .A3(new_n950), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT107), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n973));
  AOI211_X1 g548(.A(new_n973), .B(KEYINPUT44), .C1(new_n968), .C2(new_n969), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n966), .B1(new_n972), .B2(new_n974), .ZN(G397));
  INV_X1    g550(.A(G1384), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n506), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n471), .A2(new_n978), .A3(G40), .A4(new_n481), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT64), .B1(new_n469), .B2(G2105), .ZN(new_n980));
  AOI211_X1 g555(.A(new_n458), .B(new_n461), .C1(new_n467), .C2(new_n468), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n481), .B(G40), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT109), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n977), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(KEYINPUT113), .B(G8), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT114), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n983), .A2(new_n979), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n504), .B1(new_n491), .B2(new_n494), .ZN(new_n988));
  AOI21_X1  g563(.A(G1384), .B1(new_n988), .B2(new_n501), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT114), .ZN(new_n991));
  INV_X1    g566(.A(new_n985), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n986), .A2(new_n993), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n698), .A2(new_n699), .A3(G1981), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT49), .B1(new_n995), .B2(KEYINPUT117), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT49), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n997), .B(new_n998), .C1(G305), .C2(G1981), .ZN(new_n999));
  NAND2_X1  g574(.A1(G305), .A2(G1981), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n996), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1000), .B1(new_n996), .B2(new_n999), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n994), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1976), .ZN(new_n1005));
  NOR2_X1   g580(.A1(G288), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT116), .B(G1976), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT52), .B1(G288), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n991), .B1(new_n990), .B2(new_n992), .ZN(new_n1010));
  AOI211_X1 g585(.A(KEYINPUT114), .B(new_n985), .C1(new_n987), .C2(new_n989), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1007), .B(new_n1009), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1004), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1007), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1014), .B1(new_n1015), .B2(KEYINPUT115), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1006), .B1(new_n986), .B2(new_n993), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1013), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G8), .ZN(new_n1021));
  NAND3_X1  g596(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n977), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n989), .A2(KEYINPUT45), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n987), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1971), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI22_X1  g606(.A1(KEYINPUT50), .A2(new_n977), .B1(new_n983), .B2(new_n979), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n989), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(new_n753), .A3(new_n1034), .ZN(new_n1035));
  AOI211_X1 g610(.A(new_n1021), .B(new_n1025), .C1(new_n1031), .C2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1004), .A2(new_n1005), .A3(new_n712), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(G1981), .B2(G305), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1020), .A2(new_n1036), .B1(new_n1038), .B2(new_n994), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n977), .A2(KEYINPUT50), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1040), .A2(new_n987), .A3(new_n1034), .ZN(new_n1041));
  INV_X1    g616(.A(G1956), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT56), .B(G2072), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT120), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1027), .A2(new_n987), .A3(new_n1028), .A4(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n591), .A2(new_n1048), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n1043), .A2(new_n1046), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G1348), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1041), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n984), .A2(new_n795), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n621), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1043), .A2(new_n1047), .A3(new_n1049), .A4(new_n1046), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1050), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT61), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1058));
  AOI21_X1  g633(.A(G1956), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1059));
  AND4_X1   g634(.A1(new_n987), .A2(new_n1027), .A3(new_n1028), .A4(new_n1045), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1057), .B1(new_n1061), .B2(new_n1050), .ZN(new_n1062));
  AOI21_X1  g637(.A(G1348), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n990), .A2(G2067), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1063), .A2(new_n1064), .A3(new_n622), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT60), .B1(new_n1065), .B2(new_n1054), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n621), .A2(KEYINPUT60), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1070), .A2(new_n1055), .A3(KEYINPUT61), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1062), .A2(new_n1066), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  XOR2_X1   g647(.A(KEYINPUT58), .B(G1341), .Z(new_n1073));
  NAND2_X1  g648(.A1(new_n990), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1996), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1027), .A2(new_n987), .A3(new_n1028), .A4(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n566), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT122), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1074), .A2(KEYINPUT121), .A3(new_n1076), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1079), .A2(new_n1080), .A3(KEYINPUT59), .A4(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1081), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT121), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1083), .A2(new_n1084), .A3(new_n566), .ZN(new_n1085));
  XOR2_X1   g660(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1086));
  OAI21_X1  g661(.A(new_n1082), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1056), .B1(new_n1072), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1029), .A2(new_n834), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT118), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1032), .A2(new_n802), .A3(new_n1034), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1029), .A2(new_n1092), .A3(new_n834), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1090), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(G168), .A2(new_n985), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1094), .B2(G8), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1098), .B1(G168), .B2(new_n985), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1100), .B1(new_n1094), .B2(new_n992), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1096), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1088), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT124), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1017), .A2(new_n1009), .B1(new_n994), .B2(new_n1003), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT52), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1015), .A2(KEYINPUT115), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1025), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(new_n1110), .B2(new_n992), .ZN(new_n1111));
  OR2_X1    g686(.A1(new_n1111), .A2(new_n1036), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1104), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1027), .A2(new_n987), .A3(new_n1028), .A4(new_n748), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT123), .B(G1961), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1041), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n469), .A2(G2105), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1116), .A2(G2078), .ZN(new_n1121));
  AND4_X1   g696(.A1(G40), .A2(new_n481), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT108), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n989), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1026), .B1(new_n989), .B2(new_n1123), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1028), .B(new_n1122), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1117), .A2(new_n1119), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1114), .B1(new_n1128), .B2(G171), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1027), .A2(new_n987), .A3(new_n1028), .A4(new_n1121), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1117), .A2(new_n1119), .A3(G301), .A4(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT125), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1115), .A2(new_n1116), .B1(new_n1041), .B2(new_n1118), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1134), .A2(KEYINPUT125), .A3(G301), .A4(new_n1130), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1129), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(G301), .B1(new_n1134), .B2(new_n1130), .ZN(new_n1137));
  AND4_X1   g712(.A1(G301), .A2(new_n1117), .A3(new_n1119), .A4(new_n1127), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1114), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1015), .A2(KEYINPUT115), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1141), .A2(new_n1019), .A3(KEYINPUT52), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1111), .A2(new_n1036), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1142), .A2(new_n1143), .A3(KEYINPUT124), .A4(new_n1105), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1113), .A2(new_n1140), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1039), .B1(new_n1103), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1093), .A2(new_n1091), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1092), .B1(new_n1029), .B2(new_n834), .ZN(new_n1148));
  OAI211_X1 g723(.A(G168), .B(new_n992), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1109), .B1(new_n1110), .B2(G8), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1110), .A2(G8), .A3(new_n1109), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT63), .ZN(new_n1152));
  NOR4_X1   g727(.A1(new_n1108), .A2(new_n1149), .A3(new_n1150), .A4(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1149), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1142), .A2(new_n1143), .A3(new_n1154), .A4(new_n1105), .ZN(new_n1155));
  AOI21_X1  g730(.A(KEYINPUT63), .B1(new_n1155), .B2(KEYINPUT119), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT119), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1020), .A2(new_n1157), .A3(new_n1143), .A4(new_n1154), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1153), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(KEYINPUT126), .B1(new_n1146), .B2(new_n1159), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1113), .A2(new_n1144), .A3(new_n1140), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1080), .A2(KEYINPUT59), .ZN(new_n1162));
  NOR4_X1   g737(.A1(new_n1083), .A2(new_n1084), .A3(new_n566), .A4(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1086), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AND3_X1   g740(.A1(new_n1070), .A2(KEYINPUT61), .A3(new_n1055), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT61), .B1(new_n1070), .B2(new_n1055), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n622), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1052), .A2(new_n621), .A3(new_n1053), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AOI22_X1  g746(.A1(new_n1171), .A2(KEYINPUT60), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1165), .A2(new_n1168), .A3(new_n1172), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n1094), .A2(new_n992), .ZN(new_n1174));
  OAI22_X1  g749(.A1(new_n1174), .A2(new_n1100), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1173), .A2(new_n1056), .B1(new_n1175), .B2(new_n1096), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1161), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1155), .A2(KEYINPUT119), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT63), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1178), .A2(new_n1179), .A3(new_n1158), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1153), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1177), .A2(new_n1182), .A3(new_n1183), .A4(new_n1039), .ZN(new_n1184));
  OR2_X1    g759(.A1(new_n1102), .A2(KEYINPUT62), .ZN(new_n1185));
  AND2_X1   g760(.A1(new_n1113), .A2(new_n1144), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1102), .A2(KEYINPUT62), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1185), .A2(new_n1186), .A3(new_n1137), .A4(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1160), .A2(new_n1184), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(KEYINPUT45), .B1(new_n977), .B2(KEYINPUT108), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1190), .A2(new_n987), .A3(new_n1124), .ZN(new_n1191));
  XOR2_X1   g766(.A(new_n1191), .B(KEYINPUT110), .Z(new_n1192));
  XNOR2_X1  g767(.A(new_n793), .B(new_n795), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  XOR2_X1   g769(.A(new_n1194), .B(KEYINPUT111), .Z(new_n1195));
  NAND2_X1  g770(.A1(new_n1192), .A2(new_n867), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1191), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1197), .A2(new_n1075), .ZN(new_n1198));
  AOI22_X1  g773(.A1(new_n1196), .A2(new_n1198), .B1(new_n1075), .B2(new_n867), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1192), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n733), .B(new_n736), .ZN(new_n1202));
  XOR2_X1   g777(.A(new_n1202), .B(KEYINPUT112), .Z(new_n1203));
  OAI21_X1  g778(.A(new_n1200), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g779(.A(G290), .B(G1986), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1204), .B1(new_n1197), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1189), .A2(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1198), .B(KEYINPUT46), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1208), .A2(new_n1196), .A3(new_n1194), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(KEYINPUT47), .ZN(new_n1210));
  NOR3_X1   g785(.A1(new_n1191), .A2(G1986), .A3(G290), .ZN(new_n1211));
  XNOR2_X1  g786(.A(new_n1211), .B(KEYINPUT48), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1210), .B1(new_n1204), .B2(new_n1212), .ZN(new_n1213));
  NAND4_X1  g788(.A1(new_n1200), .A2(new_n731), .A3(new_n732), .A4(new_n736), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1214), .B1(G2067), .B2(new_n865), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1213), .B1(new_n1192), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1207), .A2(new_n1216), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g792(.A(G319), .ZN(new_n1219));
  NOR3_X1   g793(.A1(G227), .A2(G401), .A3(new_n1219), .ZN(new_n1220));
  NAND2_X1  g794(.A1(new_n695), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n1222));
  NAND2_X1  g796(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g797(.A1(new_n695), .A2(KEYINPUT127), .A3(new_n1220), .ZN(new_n1224));
  NAND2_X1  g798(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g799(.A1(new_n886), .A2(new_n889), .ZN(new_n1226));
  NAND3_X1  g800(.A1(new_n1225), .A2(new_n1226), .A3(new_n970), .ZN(G225));
  INV_X1    g801(.A(G225), .ZN(G308));
endmodule


