//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n996, new_n997, new_n998;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  AND2_X1   g001(.A1(new_n202), .A2(KEYINPUT83), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(KEYINPUT83), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT15), .ZN(new_n205));
  NOR3_X1   g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(KEYINPUT84), .B(G29gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(G29gat), .A2(G36gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT14), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n206), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(KEYINPUT85), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n214), .A2(new_n211), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT85), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n208), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n213), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n212), .B1(new_n206), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT17), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n220), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G15gat), .B(G22gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(G1gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(G1gat), .B2(new_n224), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n227), .B(G8gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n223), .A2(KEYINPUT86), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n221), .A2(new_n229), .A3(new_n222), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT86), .B1(new_n219), .B2(new_n228), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n230), .A2(new_n233), .B1(G229gat), .B2(G233gat), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n234), .A2(KEYINPUT18), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n229), .B(new_n219), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238));
  XOR2_X1   g037(.A(new_n238), .B(KEYINPUT13), .Z(new_n239));
  AOI22_X1  g038(.A1(new_n234), .A2(KEYINPUT18), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(KEYINPUT87), .ZN(new_n242));
  XNOR2_X1  g041(.A(G113gat), .B(G141gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT82), .B(G197gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT11), .B(G169gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n247), .B(KEYINPUT12), .Z(new_n248));
  NAND3_X1  g047(.A1(new_n241), .A2(new_n242), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n248), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n235), .B(new_n240), .C1(KEYINPUT87), .C2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT74), .ZN(new_n254));
  AND2_X1   g053(.A1(G141gat), .A2(G148gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(G141gat), .A2(G148gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G141gat), .ZN(new_n258));
  INV_X1    g057(.A(G148gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(KEYINPUT74), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT2), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT75), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT75), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT2), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n257), .A2(new_n262), .A3(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(G155gat), .B(G162gat), .Z(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G113gat), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n271), .A2(KEYINPUT68), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(KEYINPUT68), .ZN(new_n273));
  OAI21_X1  g072(.A(G120gat), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G120gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G127gat), .B(G134gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n274), .A2(new_n276), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G141gat), .B(G148gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G155gat), .ZN(new_n282));
  INV_X1    g081(.A(G162gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n263), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G134gat), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n288), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G127gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(G134gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(G127gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(new_n293), .A3(KEYINPUT67), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT1), .B1(G113gat), .B2(G120gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n276), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n290), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n270), .A2(new_n279), .A3(new_n287), .A4(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n277), .A2(new_n278), .A3(new_n276), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT68), .B(G113gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(new_n275), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n297), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT76), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT76), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n279), .A2(new_n305), .A3(new_n297), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n268), .A2(new_n269), .B1(new_n281), .B2(new_n286), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n299), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G225gat), .A2(G233gat), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT5), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT4), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT77), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n276), .A2(new_n292), .A3(new_n293), .ZN(new_n316));
  AND2_X1   g115(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n317));
  NOR2_X1   g116(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n289), .B1(new_n277), .B2(KEYINPUT67), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n274), .A2(new_n320), .B1(new_n321), .B2(new_n296), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT4), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(new_n308), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n314), .A2(new_n315), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n269), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n280), .A2(new_n254), .B1(new_n264), .B2(new_n266), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n326), .B1(new_n327), .B2(new_n262), .ZN(new_n328));
  INV_X1    g127(.A(new_n287), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT3), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n308), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n330), .A2(new_n332), .A3(new_n304), .A4(new_n306), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n298), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n325), .A2(new_n311), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n335), .A2(KEYINPUT78), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(KEYINPUT78), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n313), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G1gat), .B(G29gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT0), .ZN(new_n340));
  XNOR2_X1  g139(.A(G57gat), .B(G85gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n340), .B(new_n341), .Z(new_n342));
  AND2_X1   g141(.A1(new_n333), .A2(new_n311), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT5), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n314), .A2(new_n324), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n338), .A2(new_n342), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n342), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT78), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n343), .A2(new_n349), .A3(new_n325), .A4(new_n334), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT78), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n312), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n346), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n348), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT6), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n347), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  OAI211_X1 g155(.A(KEYINPUT6), .B(new_n348), .C1(new_n352), .C2(new_n353), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT27), .B(G183gat), .ZN(new_n359));
  INV_X1    g158(.A(G190gat), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(KEYINPUT28), .A3(new_n360), .ZN(new_n361));
  AND2_X1   g160(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT27), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OR2_X1    g163(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n365));
  AOI21_X1  g164(.A(G190gat), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n361), .B1(new_n366), .B2(KEYINPUT28), .ZN(new_n367));
  NOR2_X1   g166(.A1(G169gat), .A2(G176gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT26), .ZN(new_n369));
  NAND2_X1  g168(.A1(G183gat), .A2(G190gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G169gat), .A2(G176gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n368), .A2(KEYINPUT26), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n367), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n362), .A2(new_n363), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n370), .A2(KEYINPUT24), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT24), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n378), .A2(G183gat), .A3(G190gat), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n376), .A2(new_n360), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(G169gat), .ZN(new_n381));
  INV_X1    g180(.A(G176gat), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(new_n382), .A3(KEYINPUT23), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT23), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n384), .B1(G169gat), .B2(G176gat), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n383), .A2(new_n385), .A3(KEYINPUT25), .A4(new_n372), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT66), .B1(new_n380), .B2(new_n386), .ZN(new_n387));
  OR2_X1    g186(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(new_n360), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n377), .A2(new_n379), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n372), .B1(new_n368), .B2(KEYINPUT23), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n384), .A2(G169gat), .A3(G176gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT66), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n392), .A2(new_n395), .A3(new_n396), .A4(KEYINPUT25), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n387), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n385), .A3(new_n372), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT64), .ZN(new_n400));
  OR2_X1    g199(.A1(G183gat), .A2(G190gat), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n399), .A2(new_n400), .B1(new_n391), .B2(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n383), .A2(new_n385), .A3(KEYINPUT64), .A4(new_n372), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT25), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n375), .B1(new_n398), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G226gat), .A2(G233gat), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  OR2_X1    g207(.A1(G197gat), .A2(G204gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(G197gat), .A2(G204gat), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT22), .ZN(new_n411));
  NAND2_X1  g210(.A1(G211gat), .A2(G218gat), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n409), .A2(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n413), .A2(KEYINPUT70), .ZN(new_n414));
  XOR2_X1   g213(.A(G211gat), .B(G218gat), .Z(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n415), .B1(new_n413), .B2(KEYINPUT70), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n400), .B1(new_n393), .B2(new_n394), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n391), .A2(new_n401), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n403), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT25), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(new_n387), .A3(new_n397), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT29), .B1(new_n426), .B2(new_n375), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n408), .B(new_n420), .C1(new_n427), .C2(new_n407), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT72), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT29), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n405), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n406), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT72), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n420), .A4(new_n408), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n407), .B1(new_n405), .B2(new_n430), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT71), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n408), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n406), .B1(new_n426), .B2(new_n375), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT71), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n435), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n429), .B(new_n434), .C1(new_n440), .C2(new_n420), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G8gat), .B(G36gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(G64gat), .B(G92gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n443), .B(new_n444), .Z(new_n445));
  NAND4_X1  g244(.A1(new_n442), .A2(KEYINPUT73), .A3(KEYINPUT30), .A4(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT73), .ZN(new_n447));
  AOI211_X1 g246(.A(new_n436), .B(new_n406), .C1(new_n426), .C2(new_n375), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT71), .B1(new_n405), .B2(new_n407), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n432), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n419), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n451), .A2(new_n445), .A3(new_n429), .A4(new_n434), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT30), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n447), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n446), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n452), .A2(new_n453), .ZN(new_n456));
  INV_X1    g255(.A(new_n445), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n358), .A2(new_n455), .A3(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(KEYINPUT31), .B(G50gat), .ZN(new_n462));
  INV_X1    g261(.A(G228gat), .ZN(new_n463));
  INV_X1    g262(.A(G233gat), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n420), .B1(new_n430), .B2(new_n332), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n417), .A2(new_n430), .A3(new_n418), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n308), .B1(new_n467), .B2(new_n331), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n465), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n332), .A2(new_n430), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n419), .ZN(new_n471));
  INV_X1    g270(.A(new_n413), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT29), .B1(new_n472), .B2(new_n416), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n413), .A2(new_n415), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT3), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n475), .A2(new_n308), .ZN(new_n476));
  INV_X1    g275(.A(new_n465), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n471), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT79), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n469), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n479), .B1(new_n469), .B2(new_n478), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n462), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G78gat), .B(G106gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(G22gat), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n471), .A2(new_n476), .A3(new_n477), .ZN(new_n485));
  INV_X1    g284(.A(new_n468), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n477), .B1(new_n486), .B2(new_n471), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT79), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n469), .A2(new_n478), .A3(new_n479), .ZN(new_n489));
  INV_X1    g288(.A(new_n462), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n482), .A2(new_n484), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n484), .B1(new_n482), .B2(new_n491), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n461), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n405), .A2(new_n322), .ZN(new_n497));
  INV_X1    g296(.A(G227gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(new_n464), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n426), .A2(new_n303), .A3(new_n375), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT33), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XOR2_X1   g302(.A(G15gat), .B(G43gat), .Z(new_n504));
  XNOR2_X1  g303(.A(G71gat), .B(G99gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  AOI211_X1 g306(.A(KEYINPUT34), .B(new_n499), .C1(new_n497), .C2(new_n500), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n497), .A2(new_n500), .ZN(new_n510));
  INV_X1    g309(.A(new_n499), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT34), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n507), .A2(new_n509), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT34), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n515), .B1(new_n510), .B2(new_n511), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n503), .B(new_n506), .C1(new_n516), .C2(new_n508), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n501), .A2(KEYINPUT32), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n514), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(new_n514), .B2(new_n517), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT36), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n459), .B1(new_n454), .B2(new_n446), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n311), .B1(new_n345), .B2(new_n333), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n524), .A2(KEYINPUT80), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT80), .ZN(new_n526));
  AOI211_X1 g325(.A(new_n526), .B(new_n311), .C1(new_n345), .C2(new_n333), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT39), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(new_n310), .B2(new_n311), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n529), .B1(new_n525), .B2(new_n527), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n532), .A3(new_n342), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT40), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT40), .A4(new_n342), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(new_n354), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n494), .B1(new_n523), .B2(new_n537), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n445), .A2(KEYINPUT38), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n450), .A2(new_n420), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT37), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n435), .A2(new_n438), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n541), .B1(new_n542), .B2(new_n419), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n539), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n451), .A2(new_n541), .A3(new_n429), .A4(new_n434), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n445), .A2(new_n442), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n546), .A2(new_n356), .A3(new_n357), .ZN(new_n547));
  INV_X1    g346(.A(new_n545), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n445), .B1(new_n441), .B2(KEYINPUT37), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n548), .B1(new_n549), .B2(KEYINPUT81), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT81), .ZN(new_n551));
  NOR3_X1   g350(.A1(new_n435), .A2(new_n419), .A3(new_n438), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n419), .A2(new_n450), .B1(new_n552), .B2(new_n433), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n541), .B1(new_n553), .B2(new_n429), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n551), .B1(new_n554), .B2(new_n445), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n547), .B1(KEYINPUT38), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n496), .B(new_n522), .C1(new_n538), .C2(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n494), .A2(new_n455), .A3(new_n460), .A4(new_n521), .ZN(new_n559));
  INV_X1    g358(.A(new_n358), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT35), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n494), .A2(new_n521), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT35), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n562), .A2(new_n523), .A3(new_n563), .A4(new_n358), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n253), .B1(new_n558), .B2(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(G183gat), .B(G211gat), .Z(new_n567));
  XNOR2_X1  g366(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n568));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G57gat), .B(G64gat), .Z(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n573));
  INV_X1    g372(.A(G71gat), .ZN(new_n574));
  INV_X1    g373(.A(G78gat), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(new_n575), .A3(KEYINPUT88), .ZN(new_n576));
  NAND2_X1  g375(.A1(G71gat), .A2(G78gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n574), .A2(new_n575), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT88), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n573), .A2(new_n576), .A3(new_n577), .A4(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT89), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n572), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT9), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n577), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G57gat), .B(G64gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT89), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n583), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n581), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT90), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT21), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT91), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT92), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT91), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n591), .A2(new_n596), .A3(new_n592), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n595), .B1(new_n594), .B2(new_n597), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n571), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n600), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(new_n598), .A3(new_n570), .ZN(new_n603));
  XNOR2_X1  g402(.A(G127gat), .B(G155gat), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n601), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n605), .B1(new_n601), .B2(new_n603), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n567), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n601), .A2(new_n603), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n604), .ZN(new_n611));
  INV_X1    g410(.A(new_n567), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(new_n612), .A3(new_n606), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT95), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n591), .B(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n228), .B1(new_n616), .B2(KEYINPUT21), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n617), .A2(KEYINPUT96), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(KEYINPUT21), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n619), .A2(KEYINPUT96), .A3(new_n229), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n622), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n618), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n614), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n623), .A2(new_n625), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n628), .A2(new_n609), .A3(new_n613), .ZN(new_n629));
  NAND2_X1  g428(.A1(G85gat), .A2(G92gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT7), .ZN(new_n631));
  NAND2_X1  g430(.A1(G99gat), .A2(G106gat), .ZN(new_n632));
  INV_X1    g431(.A(G85gat), .ZN(new_n633));
  INV_X1    g432(.A(G92gat), .ZN(new_n634));
  AOI22_X1  g433(.A1(KEYINPUT8), .A2(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G99gat), .B(G106gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT98), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n640));
  INV_X1    g439(.A(new_n637), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n636), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT99), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n223), .ZN(new_n645));
  AND2_X1   g444(.A1(G232gat), .A2(G233gat), .ZN(new_n646));
  AOI22_X1  g445(.A1(new_n643), .A2(new_n219), .B1(KEYINPUT41), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(G190gat), .B(G218gat), .Z(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n649), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n645), .A2(new_n651), .A3(new_n647), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n646), .A2(KEYINPUT41), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT97), .ZN(new_n655));
  XOR2_X1   g454(.A(G134gat), .B(G162gat), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n653), .B1(KEYINPUT100), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(KEYINPUT100), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n650), .A2(new_n652), .A3(new_n659), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n643), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT10), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n616), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(new_n591), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n638), .A2(new_n581), .A3(new_n588), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(new_n663), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(G230gat), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n464), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n666), .A2(new_n667), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n671), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(G120gat), .B(G148gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(G176gat), .B(G204gat), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n677), .B(new_n678), .Z(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n676), .A2(new_n680), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n627), .A2(new_n629), .A3(new_n661), .A4(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n566), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n560), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G1gat), .ZN(G1324gat));
  INV_X1    g488(.A(new_n687), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(new_n523), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT16), .B(G8gat), .Z(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(G8gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n693), .B1(new_n694), .B2(new_n691), .ZN(new_n695));
  MUX2_X1   g494(.A(new_n693), .B(new_n695), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g495(.A(new_n521), .ZN(new_n697));
  OR3_X1    g496(.A1(new_n690), .A2(G15gat), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G15gat), .B1(new_n690), .B2(new_n522), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(G1326gat));
  NAND2_X1  g499(.A1(new_n566), .A2(new_n495), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n685), .ZN(new_n702));
  XOR2_X1   g501(.A(KEYINPUT43), .B(G22gat), .Z(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1327gat));
  NAND2_X1  g503(.A1(new_n627), .A2(new_n629), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n684), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n253), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n661), .B1(new_n558), .B2(new_n565), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(new_n358), .A3(new_n207), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT45), .Z(new_n711));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n558), .A2(new_n565), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n658), .A2(new_n660), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n712), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n455), .A2(new_n460), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n535), .A2(new_n354), .A3(new_n536), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n495), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n441), .A2(KEYINPUT37), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(KEYINPUT81), .A3(new_n457), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n545), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n549), .A2(KEYINPUT81), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT38), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n547), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n719), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT101), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n496), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n461), .A2(KEYINPUT101), .A3(new_n495), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n727), .A2(new_n729), .A3(new_n522), .A4(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n716), .B1(new_n731), .B2(new_n565), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n715), .A2(new_n732), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n733), .A2(new_n253), .A3(new_n706), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n560), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n207), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n711), .A2(new_n736), .ZN(G1328gat));
  NOR3_X1   g536(.A1(new_n709), .A2(G36gat), .A3(new_n523), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT46), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n734), .A2(new_n717), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(G36gat), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(G1329gat));
  INV_X1    g541(.A(KEYINPUT36), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n521), .B(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n734), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G43gat), .ZN(new_n746));
  OR3_X1    g545(.A1(new_n709), .A2(G43gat), .A3(new_n697), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT47), .B1(new_n747), .B2(KEYINPUT102), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1330gat));
  NOR4_X1   g549(.A1(new_n701), .A2(G50gat), .A3(new_n661), .A4(new_n706), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n495), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n751), .B1(new_n752), .B2(G50gat), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT103), .B(KEYINPUT48), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1331gat));
  INV_X1    g554(.A(new_n629), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n628), .B1(new_n609), .B2(new_n613), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n684), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n758), .A2(new_n253), .A3(new_n661), .A4(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n730), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT101), .B1(new_n461), .B2(new_n495), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n744), .B1(new_n726), .B2(new_n719), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n763), .A2(new_n764), .B1(new_n561), .B2(new_n564), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n560), .ZN(new_n767));
  XOR2_X1   g566(.A(KEYINPUT104), .B(G57gat), .Z(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(G1332gat));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n770));
  INV_X1    g569(.A(G64gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n717), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT105), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n766), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n770), .A2(new_n771), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(G1333gat));
  AOI21_X1  g575(.A(new_n574), .B1(new_n766), .B2(new_n744), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n697), .A2(G71gat), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n766), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g579(.A1(new_n766), .A2(new_n495), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g581(.A1(new_n705), .A2(new_n253), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n783), .A2(new_n684), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n715), .B2(new_n732), .ZN(new_n785));
  OAI21_X1  g584(.A(G85gat), .B1(new_n785), .B2(new_n358), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n661), .B1(new_n731), .B2(new_n565), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT106), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(KEYINPUT106), .B1(new_n765), .B2(new_n661), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n789), .A2(KEYINPUT51), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT51), .B1(new_n789), .B2(new_n790), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n759), .A2(new_n633), .A3(new_n560), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n786), .B1(new_n793), .B2(new_n794), .ZN(G1336gat));
  INV_X1    g594(.A(new_n785), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n717), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT107), .B1(new_n797), .B2(G92gat), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n759), .A2(new_n634), .A3(new_n717), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n793), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g600(.A(G99gat), .B1(new_n785), .B2(new_n522), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n684), .A2(G99gat), .A3(new_n697), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n793), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT108), .ZN(G1338gat));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n495), .B(new_n784), .C1(new_n715), .C2(new_n732), .ZN(new_n809));
  XOR2_X1   g608(.A(KEYINPUT109), .B(G106gat), .Z(new_n810));
  AND3_X1   g609(.A1(new_n809), .A2(KEYINPUT110), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT110), .B1(new_n809), .B2(new_n810), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n684), .A2(G106gat), .A3(new_n494), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT111), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n815), .B1(new_n791), .B2(new_n792), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n808), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n809), .A2(new_n810), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n808), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n731), .A2(new_n565), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n788), .A3(new_n714), .ZN(new_n822));
  INV_X1    g621(.A(new_n783), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n787), .A2(new_n788), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n820), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n789), .A2(KEYINPUT51), .A3(new_n790), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n819), .B1(new_n828), .B2(new_n814), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n807), .B1(new_n817), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT110), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n818), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n809), .A2(KEYINPUT110), .A3(new_n810), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n815), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n835), .B1(new_n826), .B2(new_n827), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT53), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n828), .A2(new_n814), .ZN(new_n838));
  INV_X1    g637(.A(new_n819), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n837), .A2(KEYINPUT112), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n830), .A2(new_n841), .ZN(G1339gat));
  NAND3_X1  g641(.A1(new_n665), .A2(new_n671), .A3(new_n668), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n673), .A2(KEYINPUT54), .A3(new_n843), .ZN(new_n844));
  AOI211_X1 g643(.A(KEYINPUT54), .B(new_n671), .C1(new_n665), .C2(new_n668), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n845), .A2(KEYINPUT113), .A3(new_n679), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n669), .A2(new_n848), .A3(new_n672), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n847), .B1(new_n849), .B2(new_n680), .ZN(new_n850));
  OAI211_X1 g649(.A(KEYINPUT55), .B(new_n844), .C1(new_n846), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT114), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT113), .B1(new_n845), .B2(new_n679), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n849), .A2(new_n847), .A3(new_n680), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n855), .A2(new_n856), .A3(KEYINPUT55), .A4(new_n844), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n661), .A2(new_n249), .A3(new_n251), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n230), .A2(new_n233), .ZN(new_n860));
  OAI22_X1  g659(.A1(new_n860), .A2(new_n238), .B1(new_n237), .B2(new_n239), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n247), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n862), .B1(new_n241), .B2(new_n248), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n714), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n855), .A2(new_n844), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT55), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n681), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n858), .A2(new_n859), .A3(new_n864), .A4(new_n867), .ZN(new_n868));
  OR3_X1    g667(.A1(new_n684), .A2(new_n863), .A3(new_n714), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n758), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n685), .A2(new_n252), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n559), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n560), .A3(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n301), .A3(new_n252), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n870), .A2(new_n871), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n495), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n560), .A2(new_n523), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n697), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(G113gat), .B1(new_n881), .B2(new_n253), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n876), .A2(new_n882), .ZN(G1340gat));
  AOI21_X1  g682(.A(G120gat), .B1(new_n875), .B2(new_n759), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n881), .A2(new_n275), .A3(new_n684), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(G1341gat));
  NAND4_X1  g685(.A1(new_n878), .A2(G127gat), .A3(new_n758), .A4(new_n880), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n887), .A2(KEYINPUT115), .ZN(new_n888));
  AOI21_X1  g687(.A(G127gat), .B1(new_n875), .B2(new_n758), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n887), .A2(KEYINPUT115), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(G1342gat));
  NAND2_X1  g690(.A1(new_n714), .A2(new_n288), .ZN(new_n892));
  OR3_X1    g691(.A1(new_n874), .A2(KEYINPUT56), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(G134gat), .B1(new_n881), .B2(new_n661), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT56), .B1(new_n874), .B2(new_n892), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT116), .ZN(G1343gat));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(KEYINPUT58), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n495), .B1(new_n870), .B2(new_n871), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT117), .ZN(new_n904));
  OAI211_X1 g703(.A(KEYINPUT57), .B(new_n495), .C1(new_n870), .C2(new_n871), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n744), .A2(new_n879), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n901), .A2(KEYINPUT117), .A3(new_n902), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n906), .A2(new_n252), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(G141gat), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n898), .A2(KEYINPUT58), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n744), .A2(new_n494), .A3(new_n717), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n872), .A2(new_n560), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n252), .A2(new_n258), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT118), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n911), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n900), .B1(new_n910), .B2(new_n917), .ZN(new_n918));
  AOI211_X1 g717(.A(new_n899), .B(new_n916), .C1(new_n909), .C2(G141gat), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(G1344gat));
  XNOR2_X1  g719(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n921));
  INV_X1    g720(.A(new_n913), .ZN(new_n922));
  AOI211_X1 g721(.A(G148gat), .B(new_n921), .C1(new_n922), .C2(new_n759), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT59), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n925), .B2(new_n684), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n684), .A2(new_n921), .ZN(new_n927));
  INV_X1    g726(.A(new_n903), .ZN(new_n928));
  INV_X1    g727(.A(new_n905), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n907), .B(new_n927), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n923), .B1(new_n931), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g731(.A(G155gat), .B1(new_n925), .B2(new_n705), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n922), .A2(new_n282), .A3(new_n758), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1346gat));
  NOR3_X1   g734(.A1(new_n925), .A2(new_n283), .A3(new_n661), .ZN(new_n936));
  AOI21_X1  g735(.A(G162gat), .B1(new_n922), .B2(new_n714), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(G1347gat));
  NOR2_X1   g737(.A1(new_n560), .A2(new_n523), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n878), .A2(new_n521), .A3(new_n939), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n940), .A2(new_n381), .A3(new_n253), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT121), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n942), .B1(new_n877), .B2(new_n560), .ZN(new_n943));
  OAI211_X1 g742(.A(KEYINPUT121), .B(new_n358), .C1(new_n870), .C2(new_n871), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n523), .A2(new_n495), .A3(new_n697), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n945), .A2(KEYINPUT122), .A3(new_n946), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n949), .A2(new_n252), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n941), .B1(new_n951), .B2(new_n381), .ZN(G1348gat));
  NAND4_X1  g751(.A1(new_n949), .A2(new_n382), .A3(new_n759), .A4(new_n950), .ZN(new_n953));
  OAI21_X1  g752(.A(G176gat), .B1(new_n940), .B2(new_n684), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1349gat));
  OAI22_X1  g754(.A1(new_n940), .A2(new_n705), .B1(new_n363), .B2(new_n362), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n945), .A2(new_n359), .A3(new_n758), .A4(new_n946), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g757(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n958), .B(new_n959), .ZN(G1350gat));
  OAI21_X1  g759(.A(G190gat), .B1(new_n940), .B2(new_n661), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT61), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n949), .A2(new_n360), .A3(new_n714), .A4(new_n950), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1351gat));
  NOR2_X1   g763(.A1(new_n928), .A2(new_n929), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n522), .A2(new_n939), .ZN(new_n966));
  XOR2_X1   g765(.A(new_n966), .B(KEYINPUT125), .Z(new_n967));
  NOR2_X1   g766(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(G197gat), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n253), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n522), .A2(new_n495), .A3(new_n717), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT124), .ZN(new_n972));
  INV_X1    g771(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n945), .A2(new_n252), .A3(new_n973), .ZN(new_n974));
  AOI22_X1  g773(.A1(new_n968), .A2(new_n970), .B1(new_n974), .B2(new_n969), .ZN(G1352gat));
  NAND2_X1  g774(.A1(new_n968), .A2(new_n759), .ZN(new_n976));
  XNOR2_X1  g775(.A(KEYINPUT126), .B(G204gat), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n684), .A2(new_n977), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n945), .A2(new_n973), .A3(new_n979), .ZN(new_n980));
  OR2_X1    g779(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n978), .A2(new_n981), .A3(new_n982), .ZN(G1353gat));
  INV_X1    g782(.A(KEYINPUT63), .ZN(new_n984));
  AOI211_X1 g783(.A(new_n705), .B(new_n967), .C1(new_n903), .C2(new_n905), .ZN(new_n985));
  INV_X1    g784(.A(G211gat), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(new_n967), .ZN(new_n988));
  OAI211_X1 g787(.A(new_n758), .B(new_n988), .C1(new_n928), .C2(new_n929), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n989), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n987), .A2(new_n990), .A3(KEYINPUT127), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n992));
  OAI211_X1 g791(.A(new_n992), .B(new_n984), .C1(new_n985), .C2(new_n986), .ZN(new_n993));
  NAND4_X1  g792(.A1(new_n945), .A2(new_n986), .A3(new_n758), .A4(new_n973), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n991), .A2(new_n993), .A3(new_n994), .ZN(G1354gat));
  INV_X1    g794(.A(G218gat), .ZN(new_n996));
  NAND4_X1  g795(.A1(new_n945), .A2(new_n996), .A3(new_n714), .A4(new_n973), .ZN(new_n997));
  NOR3_X1   g796(.A1(new_n965), .A2(new_n661), .A3(new_n967), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n997), .B1(new_n998), .B2(new_n996), .ZN(G1355gat));
endmodule


