//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT2), .ZN(new_n203));
  INV_X1    g002(.A(G141gat), .ZN(new_n204));
  INV_X1    g003(.A(G148gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n203), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G155gat), .B(G162gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT74), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(G155gat), .B2(G162gat), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n208), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n209), .B1(new_n208), .B2(new_n211), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G211gat), .ZN(new_n215));
  INV_X1    g014(.A(G218gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G211gat), .A2(G218gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT72), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT22), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT22), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT72), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n224), .A3(new_n218), .ZN(new_n225));
  XNOR2_X1  g024(.A(G197gat), .B(G204gat), .ZN(new_n226));
  AND3_X1   g025(.A1(new_n220), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n220), .B1(new_n225), .B2(new_n226), .ZN(new_n228));
  NOR3_X1   g027(.A1(new_n227), .A2(new_n228), .A3(KEYINPUT29), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n214), .B1(new_n229), .B2(KEYINPUT3), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT3), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(new_n212), .B2(new_n213), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT75), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT75), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n234), .B(new_n231), .C1(new_n212), .C2(new_n213), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT29), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n217), .A2(KEYINPUT73), .A3(new_n218), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n225), .A2(new_n237), .A3(new_n226), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n237), .B1(new_n225), .B2(new_n226), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n230), .B1(new_n236), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G228gat), .A2(G233gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT79), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT29), .ZN(new_n246));
  XNOR2_X1  g045(.A(G141gat), .B(G148gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT2), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n248), .B1(G155gat), .B2(G162gat), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n211), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n209), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n208), .A2(new_n209), .A3(new_n211), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n234), .B1(new_n254), .B2(new_n231), .ZN(new_n255));
  AOI211_X1 g054(.A(KEYINPUT75), .B(KEYINPUT3), .C1(new_n252), .C2(new_n253), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n246), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n240), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n246), .B1(new_n238), .B2(new_n239), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(new_n231), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n243), .B1(new_n260), .B2(new_n214), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n245), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n245), .B(new_n261), .C1(new_n236), .C2(new_n241), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n244), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT80), .B1(new_n265), .B2(G22gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(G78gat), .B(G106gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT31), .B(G50gat), .ZN(new_n268));
  XOR2_X1   g067(.A(new_n267), .B(new_n268), .Z(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n261), .B1(new_n236), .B2(new_n241), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT79), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n272), .A2(new_n263), .B1(new_n243), .B2(new_n242), .ZN(new_n273));
  INV_X1    g072(.A(G22gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI221_X4 g074(.A(G22gat), .B1(new_n242), .B2(new_n243), .C1(new_n272), .C2(new_n263), .ZN(new_n276));
  OAI22_X1  g075(.A1(new_n266), .A2(new_n270), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT32), .ZN(new_n278));
  INV_X1    g077(.A(G120gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G113gat), .ZN(new_n280));
  INV_X1    g079(.A(G113gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G120gat), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT1), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G127gat), .B(G134gat), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT68), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n283), .A2(KEYINPUT68), .A3(new_n284), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G127gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G134gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(new_n288), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n283), .A2(new_n292), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n286), .A2(new_n287), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT24), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT24), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n298), .A2(G183gat), .A3(G190gat), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n295), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n301), .B1(KEYINPUT23), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G169gat), .ZN(new_n304));
  INV_X1    g103(.A(G176gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(new_n305), .A3(KEYINPUT23), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT25), .ZN(new_n307));
  NOR3_X1   g106(.A1(new_n300), .A2(new_n303), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT65), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n295), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n299), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT66), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n306), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n301), .A2(KEYINPUT66), .A3(KEYINPUT23), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n303), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n314), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n308), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n304), .A2(new_n305), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT26), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n324), .A3(new_n302), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n301), .A2(KEYINPUT26), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n296), .A3(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT27), .B(G183gat), .ZN(new_n328));
  INV_X1    g127(.A(G190gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT28), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n328), .A2(KEYINPUT28), .A3(new_n329), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n327), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n294), .B1(new_n322), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n290), .A2(KEYINPUT67), .A3(G134gat), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n280), .A2(new_n282), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n289), .B(new_n336), .C1(KEYINPUT1), .C2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n287), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n338), .B1(new_n339), .B2(new_n285), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n332), .A2(new_n333), .ZN(new_n341));
  INV_X1    g140(.A(new_n327), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n303), .B1(new_n312), .B2(new_n313), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT25), .B1(new_n344), .B2(new_n318), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n340), .B(new_n343), .C1(new_n345), .C2(new_n308), .ZN(new_n346));
  NAND2_X1  g145(.A1(G227gat), .A2(G233gat), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n347), .B(KEYINPUT64), .Z(new_n348));
  NAND3_X1  g147(.A1(new_n335), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT69), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n335), .A2(new_n346), .A3(KEYINPUT69), .A4(new_n348), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n278), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  XOR2_X1   g153(.A(KEYINPUT70), .B(KEYINPUT33), .Z(new_n355));
  AOI21_X1  g154(.A(new_n355), .B1(new_n351), .B2(new_n352), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(G15gat), .B(G43gat), .Z(new_n358));
  XNOR2_X1  g157(.A(G71gat), .B(G99gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n354), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n348), .B1(new_n335), .B2(new_n346), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT34), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT71), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n362), .A2(new_n363), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT71), .B1(new_n362), .B2(new_n363), .ZN(new_n368));
  NOR3_X1   g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  AOI221_X4 g168(.A(new_n278), .B1(new_n355), .B2(new_n360), .C1(new_n351), .C2(new_n352), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n361), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  OR3_X1    g171(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n373));
  INV_X1    g172(.A(new_n360), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n353), .A2(new_n356), .A3(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n373), .B1(new_n375), .B2(new_n370), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n265), .A2(G22gat), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n274), .B(new_n244), .C1(new_n262), .C2(new_n264), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n377), .A2(KEYINPUT80), .A3(new_n378), .A4(new_n269), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n277), .A2(new_n372), .A3(new_n376), .A4(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G8gat), .B(G36gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(G64gat), .B(G92gat), .ZN(new_n382));
  XOR2_X1   g181(.A(new_n381), .B(new_n382), .Z(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(G226gat), .A2(G233gat), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n343), .B1(new_n345), .B2(new_n308), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n386), .B1(new_n387), .B2(new_n246), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n320), .A2(new_n321), .ZN(new_n389));
  INV_X1    g188(.A(new_n308), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n334), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(new_n385), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n388), .A2(new_n392), .A3(new_n240), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n385), .B1(new_n391), .B2(KEYINPUT29), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n387), .A2(new_n386), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n241), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n384), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n240), .B1(new_n388), .B2(new_n392), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n394), .A2(new_n241), .A3(new_n395), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n399), .A3(new_n383), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n397), .A2(KEYINPUT30), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT30), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n398), .A2(new_n399), .A3(new_n402), .A4(new_n383), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT4), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n294), .A2(new_n406), .A3(new_n254), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT4), .B1(new_n340), .B2(new_n214), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT78), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n214), .A2(KEYINPUT3), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n340), .B(new_n411), .C1(new_n255), .C2(new_n256), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n286), .A2(new_n287), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n413), .A2(new_n254), .A3(new_n338), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n414), .A2(KEYINPUT78), .A3(KEYINPUT4), .ZN(new_n415));
  NAND2_X1  g214(.A1(G225gat), .A2(G233gat), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n416), .B(KEYINPUT76), .Z(new_n417));
  NOR2_X1   g216(.A1(new_n417), .A2(KEYINPUT5), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n410), .A2(new_n412), .A3(new_n415), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n340), .A2(new_n214), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(new_n414), .A3(KEYINPUT77), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT77), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n340), .A2(new_n422), .A3(new_n214), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n417), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT5), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n407), .A2(new_n408), .ZN(new_n426));
  INV_X1    g225(.A(new_n417), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n412), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n419), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G1gat), .B(G29gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT0), .ZN(new_n431));
  XNOR2_X1  g230(.A(G57gat), .B(G85gat), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n431), .B(new_n432), .Z(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n433), .B(new_n419), .C1(new_n425), .C2(new_n428), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n429), .A2(KEYINPUT6), .A3(new_n434), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n405), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT35), .B1(new_n380), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n379), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT80), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n444), .B1(new_n273), .B2(new_n274), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n445), .A2(new_n269), .B1(new_n377), .B2(new_n378), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT35), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n376), .A2(new_n372), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n404), .B1(new_n439), .B2(new_n438), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n447), .A2(new_n448), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n442), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT82), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT36), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n373), .A2(new_n375), .A3(new_n370), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n369), .B1(new_n361), .B2(new_n371), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n376), .A2(new_n372), .A3(KEYINPUT36), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n410), .A2(new_n412), .A3(new_n415), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n417), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT39), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n421), .A2(new_n423), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n462), .B1(new_n463), .B2(new_n427), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n460), .A2(new_n462), .A3(new_n417), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n433), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT40), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n465), .A2(KEYINPUT40), .A3(new_n433), .A4(new_n466), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n404), .A2(new_n469), .A3(new_n435), .A4(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n400), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT37), .B1(new_n393), .B2(new_n396), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT37), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n398), .A2(new_n399), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n473), .A2(new_n475), .A3(new_n384), .ZN(new_n476));
  XOR2_X1   g275(.A(KEYINPUT81), .B(KEYINPUT38), .Z(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n472), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n473), .A2(new_n477), .A3(new_n475), .A4(new_n384), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n479), .A2(new_n438), .A3(new_n439), .A4(new_n480), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n471), .A2(new_n481), .A3(new_n379), .A4(new_n277), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n277), .A2(new_n379), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n441), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n459), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n452), .A2(new_n453), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n453), .B1(new_n452), .B2(new_n485), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G15gat), .B(G22gat), .ZN(new_n489));
  INV_X1    g288(.A(G1gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT16), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n492), .B1(G1gat), .B2(new_n489), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT84), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n494), .B1(new_n489), .B2(G1gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(G8gat), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G8gat), .ZN(new_n497));
  OAI221_X1 g296(.A(new_n492), .B1(new_n494), .B2(new_n497), .C1(G1gat), .C2(new_n489), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT85), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT15), .ZN(new_n502));
  OR2_X1    g301(.A1(G43gat), .A2(G50gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(G43gat), .A2(G50gat), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(KEYINPUT83), .B(G43gat), .ZN(new_n506));
  INV_X1    g305(.A(G50gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(KEYINPUT14), .B(G29gat), .ZN(new_n511));
  INV_X1    g310(.A(G36gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G29gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n505), .B1(new_n510), .B2(new_n516), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n516), .A2(new_n505), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n496), .A2(new_n498), .A3(KEYINPUT85), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n501), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT17), .B1(new_n517), .B2(new_n518), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT17), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n516), .A2(new_n505), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n513), .A2(new_n515), .B1(new_n508), .B2(new_n509), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n523), .B(new_n524), .C1(new_n525), .C2(new_n505), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n522), .A2(new_n498), .A3(new_n496), .A4(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G229gat), .A2(G233gat), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n521), .A2(new_n527), .A3(KEYINPUT18), .A4(new_n528), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n529), .A2(KEYINPUT88), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n521), .A2(KEYINPUT89), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT89), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n501), .A2(new_n532), .A3(new_n519), .A4(new_n520), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n501), .A2(new_n520), .ZN(new_n534));
  INV_X1    g333(.A(new_n519), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n531), .A2(new_n533), .A3(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n528), .B(KEYINPUT13), .Z(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n529), .A2(KEYINPUT88), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n530), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n521), .A2(new_n527), .A3(new_n528), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT86), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT18), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT86), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n521), .A2(new_n527), .A3(new_n545), .A4(new_n528), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G113gat), .B(G141gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(G197gat), .ZN(new_n549));
  XOR2_X1   g348(.A(KEYINPUT11), .B(G169gat), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n551), .B(KEYINPUT12), .Z(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n541), .B(new_n547), .C1(KEYINPUT87), .C2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n547), .A2(new_n530), .A3(new_n539), .A4(new_n540), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n530), .A2(new_n539), .A3(KEYINPUT87), .A4(new_n540), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(new_n556), .A3(new_n552), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT94), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(G232gat), .A2(G233gat), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT41), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n561), .B(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G85gat), .A2(G92gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT7), .ZN(new_n569));
  NAND2_X1  g368(.A1(G99gat), .A2(G106gat), .ZN(new_n570));
  INV_X1    g369(.A(G85gat), .ZN(new_n571));
  INV_X1    g370(.A(G92gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(KEYINPUT8), .A2(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G99gat), .B(G106gat), .Z(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n575), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n577), .A2(new_n569), .A3(new_n573), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  OAI22_X1  g378(.A1(new_n535), .A2(new_n579), .B1(new_n564), .B2(new_n563), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n522), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n526), .A2(new_n579), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT93), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NOR3_X1   g384(.A1(new_n582), .A2(new_n583), .A3(KEYINPUT93), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n581), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n559), .A2(new_n560), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G134gat), .B(G162gat), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n587), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n591), .B1(new_n587), .B2(new_n589), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n567), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n594), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(new_n566), .A3(new_n592), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT90), .ZN(new_n599));
  INV_X1    g398(.A(G57gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n599), .B1(new_n600), .B2(G64gat), .ZN(new_n601));
  INV_X1    g400(.A(G64gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(KEYINPUT90), .A3(G57gat), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n601), .B(new_n603), .C1(G57gat), .C2(new_n602), .ZN(new_n604));
  NAND2_X1  g403(.A1(G71gat), .A2(G78gat), .ZN(new_n605));
  OR2_X1    g404(.A1(G71gat), .A2(G78gat), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT9), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n600), .A2(G64gat), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n602), .A2(G57gat), .ZN(new_n611));
  OAI21_X1  g410(.A(KEYINPUT9), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n606), .A2(new_n605), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT92), .ZN(new_n616));
  AOI22_X1  g415(.A1(new_n608), .A2(new_n604), .B1(new_n612), .B2(new_n613), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT92), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n616), .A2(new_n619), .A3(KEYINPUT21), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n534), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n617), .A2(KEYINPUT21), .ZN(new_n622));
  XNOR2_X1  g421(.A(G127gat), .B(G155gat), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n622), .B(new_n623), .Z(new_n624));
  XNOR2_X1  g423(.A(new_n621), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G231gat), .A2(G233gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT91), .ZN(new_n627));
  XOR2_X1   g426(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G183gat), .B(G211gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n625), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n575), .A2(KEYINPUT95), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n609), .A2(new_n614), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n579), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT10), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n617), .A2(new_n576), .A3(new_n578), .A4(new_n633), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n576), .A2(new_n578), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n639), .A2(new_n616), .A3(KEYINPUT10), .A4(new_n619), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G230gat), .A2(G233gat), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n635), .A2(new_n637), .ZN(new_n644));
  INV_X1    g443(.A(new_n642), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g446(.A(G120gat), .B(G148gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT96), .ZN(new_n649));
  XNOR2_X1  g448(.A(G176gat), .B(G204gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(KEYINPUT97), .B1(new_n647), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT97), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n643), .A2(new_n654), .A3(new_n646), .A4(new_n651), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n651), .B(KEYINPUT98), .Z(new_n657));
  NAND2_X1  g456(.A1(new_n647), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n598), .A2(new_n632), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n488), .A2(new_n558), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n440), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n662), .A2(KEYINPUT99), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(KEYINPUT99), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(new_n490), .ZN(G1324gat));
  INV_X1    g467(.A(new_n661), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT16), .B(G8gat), .Z(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(new_n404), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(G8gat), .B1(new_n661), .B2(new_n405), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT42), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(G1325gat));
  INV_X1    g476(.A(G15gat), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n669), .A2(new_n678), .A3(new_n449), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n459), .A2(KEYINPUT100), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n681), .B1(new_n457), .B2(new_n458), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(G15gat), .B1(new_n661), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT101), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n679), .A2(KEYINPUT101), .A3(new_n685), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(G1326gat));
  NOR2_X1   g489(.A1(new_n661), .A2(new_n447), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT43), .B(G22gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  INV_X1    g492(.A(new_n598), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(new_n486), .B2(new_n487), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n452), .A2(new_n485), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n598), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(new_n695), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n558), .ZN(new_n702));
  INV_X1    g501(.A(new_n659), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n632), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G29gat), .B1(new_n706), .B2(new_n666), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n694), .A2(new_n704), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n558), .B(new_n708), .C1(new_n486), .C2(new_n487), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(G29gat), .A3(new_n666), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n712), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n707), .A2(new_n713), .A3(new_n714), .ZN(G1328gat));
  OAI21_X1  g514(.A(G36gat), .B1(new_n706), .B2(new_n405), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n709), .A2(G36gat), .A3(new_n405), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n716), .A2(new_n719), .A3(new_n720), .ZN(G1329gat));
  INV_X1    g520(.A(new_n459), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n697), .A2(new_n722), .A3(new_n700), .A4(new_n705), .ZN(new_n723));
  INV_X1    g522(.A(new_n506), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n449), .A2(new_n506), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n725), .B(KEYINPUT47), .C1(new_n709), .C2(new_n726), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n697), .A2(new_n683), .A3(new_n700), .A4(new_n705), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n728), .A2(KEYINPUT103), .A3(new_n724), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT103), .B1(new_n728), .B2(new_n724), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n709), .A2(new_n726), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n727), .B1(new_n732), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g532(.A(new_n709), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n447), .A2(G50gat), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n697), .A2(new_n483), .A3(new_n700), .A4(new_n705), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G50gat), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n734), .A2(KEYINPUT105), .A3(new_n735), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n738), .A2(KEYINPUT48), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n736), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT48), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT104), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI22_X1  g544(.A1(new_n739), .A2(G50gat), .B1(new_n734), .B2(new_n735), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT104), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n746), .A2(new_n747), .A3(KEYINPUT48), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n742), .B1(new_n745), .B2(new_n748), .ZN(G1331gat));
  NOR2_X1   g548(.A1(new_n598), .A2(new_n632), .ZN(new_n750));
  AND4_X1   g549(.A1(new_n702), .A2(new_n698), .A3(new_n750), .A4(new_n659), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n665), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g552(.A(new_n405), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT106), .ZN(new_n756));
  NOR2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1333gat));
  INV_X1    g557(.A(G71gat), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n751), .A2(new_n759), .A3(new_n449), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n751), .A2(new_n683), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n761), .B2(new_n759), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g562(.A1(new_n751), .A2(new_n483), .ZN(new_n764));
  XNOR2_X1  g563(.A(KEYINPUT107), .B(G78gat), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1335gat));
  INV_X1    g565(.A(new_n632), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n558), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n703), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n701), .A2(new_n665), .A3(new_n770), .ZN(new_n771));
  AND2_X1   g570(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n772));
  NOR2_X1   g571(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n698), .A2(new_n598), .A3(new_n768), .A4(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n699), .A2(new_n769), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n777), .B2(new_n772), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n665), .A2(new_n571), .A3(new_n659), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n771), .A2(new_n571), .B1(new_n779), .B2(new_n780), .ZN(G1336gat));
  NAND4_X1  g580(.A1(new_n697), .A2(new_n404), .A3(new_n700), .A4(new_n770), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n404), .A2(new_n572), .A3(new_n659), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n783), .B(KEYINPUT109), .Z(new_n784));
  AOI22_X1  g583(.A1(G92gat), .A2(new_n782), .B1(new_n778), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1337gat));
  NOR2_X1   g586(.A1(new_n703), .A2(G99gat), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n778), .A2(new_n449), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n701), .A2(new_n683), .A3(new_n770), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT110), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G99gat), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n790), .A2(KEYINPUT110), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n789), .B1(new_n792), .B2(new_n793), .ZN(G1338gat));
  NAND4_X1  g593(.A1(new_n697), .A2(new_n483), .A3(new_n700), .A4(new_n770), .ZN(new_n795));
  XOR2_X1   g594(.A(KEYINPUT111), .B(G106gat), .Z(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n447), .A2(G106gat), .A3(new_n703), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n778), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n797), .A2(new_n799), .A3(KEYINPUT112), .ZN(new_n800));
  XNOR2_X1  g599(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n800), .B(new_n801), .ZN(G1339gat));
  OAI21_X1  g601(.A(KEYINPUT114), .B1(new_n641), .B2(new_n642), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n638), .A2(new_n640), .A3(new_n804), .A4(new_n645), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n645), .B1(new_n638), .B2(new_n640), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n651), .B1(new_n807), .B2(new_n808), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(KEYINPUT55), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n656), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT55), .B1(new_n810), .B2(new_n811), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n557), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n555), .B1(new_n556), .B2(new_n552), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n541), .A2(new_n553), .A3(new_n547), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n537), .A2(new_n538), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n528), .B1(new_n521), .B2(new_n527), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n551), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(new_n659), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n598), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n597), .A2(new_n595), .A3(new_n819), .A4(new_n822), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n825), .A2(new_n814), .A3(new_n813), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n632), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n660), .A2(new_n702), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n447), .ZN(new_n830));
  INV_X1    g629(.A(new_n449), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n665), .A2(new_n405), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n281), .B1(new_n833), .B2(new_n558), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT115), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n666), .B1(new_n827), .B2(new_n828), .ZN(new_n836));
  INV_X1    g635(.A(new_n380), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n404), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT116), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n840), .A2(new_n281), .A3(new_n558), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n835), .A2(new_n841), .ZN(G1340gat));
  NAND3_X1  g641(.A1(new_n840), .A2(new_n279), .A3(new_n659), .ZN(new_n843));
  OR3_X1    g642(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n844));
  OAI21_X1  g643(.A(G120gat), .B1(new_n844), .B2(new_n703), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(G1341gat));
  NAND3_X1  g645(.A1(new_n833), .A2(G127gat), .A3(new_n767), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n836), .A2(new_n837), .A3(new_n405), .A4(new_n767), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(KEYINPUT117), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n290), .B1(new_n848), .B2(KEYINPUT117), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n851), .B(new_n852), .ZN(G1342gat));
  OAI21_X1  g652(.A(G134gat), .B1(new_n844), .B2(new_n694), .ZN(new_n854));
  OR3_X1    g653(.A1(new_n694), .A2(G134gat), .A3(new_n404), .ZN(new_n855));
  OR3_X1    g654(.A1(new_n838), .A2(KEYINPUT56), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT56), .B1(new_n838), .B2(new_n855), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n854), .A2(new_n856), .A3(KEYINPUT119), .A4(new_n857), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1343gat));
  OAI21_X1  g661(.A(new_n483), .B1(new_n680), .B2(new_n682), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT121), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n865), .B(new_n483), .C1(new_n680), .C2(new_n682), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n836), .A2(new_n864), .A3(new_n405), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n558), .A2(new_n204), .ZN(new_n868));
  XOR2_X1   g667(.A(new_n868), .B(KEYINPUT122), .Z(new_n869));
  NOR2_X1   g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n832), .A2(new_n722), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT57), .B1(new_n829), .B2(new_n483), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n483), .A2(KEYINPUT57), .ZN(new_n873));
  INV_X1    g672(.A(new_n814), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n874), .A2(KEYINPUT120), .A3(new_n656), .A4(new_n812), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n876), .B1(new_n813), .B2(new_n814), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n558), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n598), .B1(new_n878), .B2(new_n823), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n632), .B1(new_n879), .B2(new_n826), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n873), .B1(new_n880), .B2(new_n828), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n558), .B(new_n871), .C1(new_n872), .C2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n870), .B1(G141gat), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n882), .B2(G141gat), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n883), .A2(new_n885), .A3(KEYINPUT58), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887));
  AOI221_X4 g686(.A(new_n870), .B1(new_n884), .B2(new_n887), .C1(G141gat), .C2(new_n882), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n886), .A2(new_n888), .ZN(G1344gat));
  NAND2_X1  g688(.A1(new_n880), .A2(new_n828), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT57), .B1(new_n890), .B2(new_n483), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n827), .A2(new_n828), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n873), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n871), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n703), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  OAI211_X1 g696(.A(KEYINPUT59), .B(G148gat), .C1(new_n894), .C2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT59), .B1(new_n867), .B2(new_n703), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n205), .ZN(new_n900));
  INV_X1    g699(.A(new_n872), .ZN(new_n901));
  INV_X1    g700(.A(new_n881), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(new_n904), .A3(new_n896), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n898), .A2(new_n900), .A3(new_n905), .ZN(G1345gat));
  NAND2_X1  g705(.A1(new_n903), .A2(new_n871), .ZN(new_n907));
  OAI21_X1  g706(.A(G155gat), .B1(new_n907), .B2(new_n632), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n867), .A2(G155gat), .A3(new_n632), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n908), .A2(KEYINPUT124), .A3(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n912));
  INV_X1    g711(.A(G155gat), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n895), .B1(new_n901), .B2(new_n902), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n767), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n912), .B1(new_n915), .B2(new_n909), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n911), .A2(new_n916), .ZN(G1346gat));
  OAI21_X1  g716(.A(G162gat), .B1(new_n907), .B2(new_n694), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n694), .A2(G162gat), .A3(new_n404), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n836), .A2(new_n864), .A3(new_n866), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1347gat));
  NAND2_X1  g720(.A1(new_n666), .A2(new_n404), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(new_n831), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n447), .A3(new_n829), .ZN(new_n924));
  OAI21_X1  g723(.A(G169gat), .B1(new_n924), .B2(new_n702), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT125), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n892), .A2(new_n665), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n380), .A2(new_n405), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n304), .A3(new_n558), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n926), .A2(new_n931), .ZN(G1348gat));
  OAI21_X1  g731(.A(G176gat), .B1(new_n924), .B2(new_n703), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n659), .A2(new_n305), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n929), .B2(new_n934), .ZN(G1349gat));
  NAND3_X1  g734(.A1(new_n930), .A2(new_n328), .A3(new_n767), .ZN(new_n936));
  OAI21_X1  g735(.A(G183gat), .B1(new_n924), .B2(new_n632), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT60), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT60), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n936), .A2(new_n940), .A3(new_n937), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1350gat));
  OAI21_X1  g741(.A(G190gat), .B1(new_n924), .B2(new_n694), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT61), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n930), .A2(new_n329), .A3(new_n598), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1351gat));
  NOR4_X1   g745(.A1(new_n892), .A2(new_n405), .A3(new_n665), .A4(new_n863), .ZN(new_n947));
  AOI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n558), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n894), .A2(new_n683), .A3(new_n922), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n558), .A2(G197gat), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(G1352gat));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n659), .ZN(new_n952));
  XNOR2_X1  g751(.A(KEYINPUT126), .B(G204gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n703), .A2(new_n953), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n947), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g755(.A(new_n956), .B(KEYINPUT62), .Z(new_n957));
  NAND2_X1  g756(.A1(new_n954), .A2(new_n957), .ZN(G1353gat));
  NAND3_X1  g757(.A1(new_n947), .A2(new_n215), .A3(new_n767), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n922), .A2(new_n683), .ZN(new_n960));
  OAI211_X1 g759(.A(new_n767), .B(new_n960), .C1(new_n891), .C2(new_n893), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n961), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT63), .B1(new_n961), .B2(G211gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(G1354gat));
  OAI21_X1  g763(.A(new_n960), .B1(new_n891), .B2(new_n893), .ZN(new_n965));
  OAI21_X1  g764(.A(G218gat), .B1(new_n965), .B2(new_n694), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n947), .A2(new_n216), .A3(new_n598), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n966), .A2(new_n967), .A3(KEYINPUT127), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(G1355gat));
endmodule


