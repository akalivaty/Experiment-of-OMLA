//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT73), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G125), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G140), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT72), .B1(new_n195), .B2(G146), .ZN(new_n196));
  XNOR2_X1  g010(.A(G125), .B(G140), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT72), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n196), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT16), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(new_n191), .A3(G125), .ZN(new_n203));
  OAI211_X1 g017(.A(G146), .B(new_n203), .C1(new_n195), .C2(new_n202), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT24), .B(G110), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT65), .A2(G128), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(G119), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT68), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT69), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n214), .B1(new_n209), .B2(G119), .ZN(new_n215));
  INV_X1    g029(.A(G119), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT69), .A3(G128), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n212), .A2(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n210), .A2(KEYINPUT68), .A3(G119), .A4(new_n211), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n207), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT71), .ZN(new_n221));
  INV_X1    g035(.A(G110), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT23), .B1(new_n209), .B2(G119), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT70), .B1(new_n216), .B2(G128), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(new_n209), .A3(G119), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n223), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n210), .A2(KEYINPUT23), .A3(G119), .A4(new_n211), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n220), .A2(new_n221), .B1(new_n222), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n212), .A2(new_n213), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n215), .A2(new_n217), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n219), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n206), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT71), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n205), .B1(new_n230), .B2(new_n235), .ZN(new_n236));
  OR2_X1    g050(.A1(new_n229), .A2(new_n222), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n218), .A2(new_n207), .A3(new_n219), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n203), .B1(new_n195), .B2(new_n202), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n199), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(new_n204), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n237), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n190), .B1(new_n236), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n205), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n229), .A2(new_n222), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n246), .B1(new_n234), .B2(KEYINPUT71), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n220), .A2(new_n221), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n245), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(KEYINPUT73), .A3(new_n242), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT22), .B(G137), .ZN(new_n251));
  INV_X1    g065(.A(G953), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n252), .A2(G221), .A3(G234), .ZN(new_n253));
  XOR2_X1   g067(.A(new_n251), .B(new_n253), .Z(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n244), .A2(new_n250), .A3(new_n255), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n190), .B(new_n254), .C1(new_n236), .C2(new_n243), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT25), .B1(new_n258), .B2(new_n188), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT25), .ZN(new_n260));
  AOI211_X1 g074(.A(new_n260), .B(G902), .C1(new_n256), .C2(new_n257), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n189), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n189), .A2(G902), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n199), .A2(G143), .ZN(new_n266));
  INV_X1    g080(.A(G143), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G146), .ZN(new_n268));
  AND2_X1   g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(G143), .B(G146), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT0), .B(G128), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT64), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT11), .ZN(new_n276));
  INV_X1    g090(.A(G134), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(G137), .ZN(new_n278));
  INV_X1    g092(.A(G137), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(KEYINPUT11), .A3(G134), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n277), .A2(G137), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G131), .ZN(new_n283));
  INV_X1    g097(.A(G131), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n278), .A2(new_n280), .A3(new_n284), .A4(new_n281), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n270), .B(KEYINPUT64), .C1(new_n271), .C2(new_n272), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n275), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n266), .A2(new_n268), .ZN(new_n289));
  AND2_X1   g103(.A1(KEYINPUT65), .A2(G128), .ZN(new_n290));
  NOR2_X1   g104(.A1(KEYINPUT65), .A2(G128), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT1), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n293), .B1(G143), .B2(new_n199), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n289), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n271), .A2(new_n293), .A3(G128), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n277), .A2(G137), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n279), .A2(G134), .ZN(new_n299));
  OAI21_X1  g113(.A(G131), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n285), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT30), .B1(new_n288), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n285), .A2(new_n300), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n304), .B1(new_n295), .B2(new_n296), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n273), .B1(new_n285), .B2(new_n283), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT30), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(KEYINPUT2), .A2(G113), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NOR3_X1   g125(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(G116), .B(G119), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n314), .B(new_n309), .C1(new_n311), .C2(new_n312), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n303), .A2(new_n308), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n273), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n297), .A2(new_n301), .B1(new_n286), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n319), .ZN(new_n323));
  INV_X1    g137(.A(G237), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(new_n252), .A3(G210), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(KEYINPUT27), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT26), .B(G101), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n326), .B(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT31), .B1(new_n320), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n288), .A2(new_n302), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n318), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n333), .B1(new_n322), .B2(new_n319), .ZN(new_n334));
  NOR4_X1   g148(.A1(new_n305), .A2(new_n306), .A3(new_n318), .A4(KEYINPUT28), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n332), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n328), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n331), .A2(new_n307), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n322), .A2(KEYINPUT30), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n318), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n286), .A2(new_n321), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n302), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(new_n318), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n344), .A2(new_n337), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT31), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n341), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n330), .A2(new_n338), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(G472), .A2(G902), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT32), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(KEYINPUT67), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n336), .A2(new_n328), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n344), .A2(new_n328), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n341), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(KEYINPUT29), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n343), .A2(new_n318), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n356), .B1(new_n334), .B2(new_n335), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n328), .A2(KEYINPUT29), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n188), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(G472), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n348), .A2(KEYINPUT32), .A3(new_n349), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n265), .B1(new_n351), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n273), .A2(G125), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n364), .B1(new_n297), .B2(G125), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT80), .B(G224), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(G953), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n365), .B(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT78), .ZN(new_n369));
  INV_X1    g183(.A(G104), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT3), .B1(new_n370), .B2(G107), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n372));
  INV_X1    g186(.A(G107), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(G104), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n370), .A2(G107), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G101), .ZN(new_n377));
  INV_X1    g191(.A(G101), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n371), .A2(new_n374), .A3(new_n378), .A4(new_n375), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(KEYINPUT4), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n318), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT76), .ZN(new_n382));
  OR2_X1    g196(.A1(KEYINPUT75), .A2(KEYINPUT4), .ZN(new_n383));
  NAND2_X1  g197(.A1(KEYINPUT75), .A2(KEYINPUT4), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n378), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n376), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n382), .B1(new_n376), .B2(new_n385), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n369), .B1(new_n381), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n387), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n376), .A2(new_n385), .A3(new_n382), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n392), .A2(KEYINPUT78), .A3(new_n318), .A4(new_n380), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n314), .A2(KEYINPUT5), .ZN(new_n394));
  INV_X1    g208(.A(G113), .ZN(new_n395));
  INV_X1    g209(.A(G116), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(G119), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT5), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n395), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n394), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n317), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n370), .A2(G107), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n373), .A2(G104), .ZN(new_n403));
  OAI21_X1  g217(.A(G101), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n379), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(G110), .B(G122), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n389), .A2(new_n393), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n389), .A2(new_n393), .A3(new_n407), .ZN(new_n410));
  INV_X1    g224(.A(new_n408), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT79), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  AOI22_X1  g227(.A1(KEYINPUT6), .A2(new_n409), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n318), .B(new_n380), .C1(new_n386), .C2(new_n387), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n406), .B1(new_n416), .B2(new_n369), .ZN(new_n417));
  AOI211_X1 g231(.A(new_n415), .B(new_n412), .C1(new_n417), .C2(new_n393), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n368), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT7), .B1(new_n366), .B2(G953), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n365), .B(new_n420), .ZN(new_n421));
  XOR2_X1   g235(.A(new_n408), .B(KEYINPUT8), .Z(new_n422));
  INV_X1    g236(.A(new_n401), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n422), .B1(new_n423), .B2(new_n405), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT83), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT82), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n399), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n394), .A2(KEYINPUT81), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT81), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n314), .A2(new_n429), .A3(KEYINPUT5), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n399), .A2(new_n426), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n427), .A2(new_n428), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n432), .A2(new_n317), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n424), .B(new_n425), .C1(new_n433), .C2(new_n405), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n405), .B1(new_n432), .B2(new_n317), .ZN(new_n435));
  INV_X1    g249(.A(new_n422), .ZN(new_n436));
  INV_X1    g250(.A(new_n405), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n436), .B1(new_n401), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT83), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n421), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(G902), .B1(new_n440), .B2(new_n409), .ZN(new_n441));
  OAI21_X1  g255(.A(G210), .B1(G237), .B2(G902), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n419), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT84), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n419), .A2(new_n441), .ZN(new_n445));
  INV_X1    g259(.A(new_n442), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT84), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n419), .A2(new_n441), .A3(new_n448), .A4(new_n442), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n444), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G214), .B1(G237), .B2(G902), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G221), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT9), .B(G234), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n453), .B1(new_n455), .B2(new_n188), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n456), .B(KEYINPUT74), .Z(new_n457));
  INV_X1    g271(.A(G469), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n380), .B(new_n321), .C1(new_n386), .C2(new_n387), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n266), .A2(KEYINPUT1), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n271), .B1(G128), .B2(new_n460), .ZN(new_n461));
  AND4_X1   g275(.A1(new_n293), .A2(new_n266), .A3(new_n268), .A4(G128), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n379), .B(new_n404), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT10), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n283), .A2(new_n285), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n437), .A2(new_n297), .A3(KEYINPUT10), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n459), .A2(new_n465), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT77), .ZN(new_n469));
  XNOR2_X1  g283(.A(G110), .B(G140), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n252), .A2(G227), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n470), .B(new_n471), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n468), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n469), .B1(new_n468), .B2(new_n472), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT12), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n405), .A2(new_n295), .A3(new_n296), .ZN(new_n476));
  AOI211_X1 g290(.A(new_n475), .B(new_n466), .C1(new_n463), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n463), .A2(new_n476), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT12), .B1(new_n478), .B2(new_n286), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n473), .A2(new_n474), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n459), .A2(new_n465), .A3(new_n467), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n286), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n472), .B1(new_n483), .B2(new_n468), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n458), .B(new_n188), .C1(new_n481), .C2(new_n484), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n468), .A2(new_n472), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n468), .B1(new_n477), .B2(new_n479), .ZN(new_n487));
  INV_X1    g301(.A(new_n472), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n483), .A2(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(G469), .B1(new_n489), .B2(G902), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n457), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n324), .A2(new_n252), .A3(G214), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n267), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n324), .A2(new_n252), .A3(G143), .A4(G214), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(G131), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT17), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n494), .A2(new_n284), .A3(new_n495), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT88), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n496), .A2(KEYINPUT17), .A3(G131), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n503), .A2(new_n240), .A3(new_n204), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n497), .A2(KEYINPUT88), .A3(new_n498), .A4(new_n499), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(G113), .B(G122), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT87), .B(G104), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n507), .B(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(KEYINPUT18), .A2(G131), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n510), .B1(new_n494), .B2(new_n495), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n195), .A2(G146), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n511), .B1(new_n201), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n494), .A2(new_n495), .A3(new_n510), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT85), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT85), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n494), .A2(new_n516), .A3(new_n495), .A4(new_n510), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n513), .A2(KEYINPUT86), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT86), .B1(new_n513), .B2(new_n518), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n506), .B(new_n509), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n197), .B(KEYINPUT19), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n199), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n497), .A2(new_n499), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n523), .A2(new_n204), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT86), .ZN(new_n526));
  INV_X1    g340(.A(new_n518), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n198), .B1(new_n197), .B2(new_n199), .ZN(new_n528));
  AND4_X1   g342(.A1(new_n198), .A2(new_n192), .A3(new_n194), .A4(new_n199), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n512), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n511), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n526), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n513), .A2(new_n518), .A3(KEYINPUT86), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n525), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n521), .B1(new_n535), .B2(new_n509), .ZN(new_n536));
  NOR2_X1   g350(.A1(G475), .A2(G902), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT20), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT20), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n536), .A2(new_n540), .A3(new_n537), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n252), .A2(G952), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n543), .B1(G234), .B2(G237), .ZN(new_n544));
  AOI211_X1 g358(.A(new_n188), .B(new_n252), .C1(G234), .C2(G237), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT21), .B(G898), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n506), .B1(new_n519), .B2(new_n520), .ZN(new_n549));
  INV_X1    g363(.A(new_n509), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(G902), .B1(new_n551), .B2(new_n521), .ZN(new_n552));
  INV_X1    g366(.A(G475), .ZN(new_n553));
  OR2_X1    g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n290), .A2(new_n291), .A3(new_n267), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT13), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n556), .B1(new_n209), .B2(G143), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n267), .A2(KEYINPUT13), .A3(G128), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(G134), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n210), .A2(G143), .A3(new_n211), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n267), .A2(G128), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n277), .A3(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n396), .A2(G122), .ZN(new_n564));
  INV_X1    g378(.A(G122), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n565), .A2(G116), .ZN(new_n566));
  OAI21_X1  g380(.A(G107), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(G116), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n396), .A2(G122), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n569), .A3(new_n373), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n560), .A2(new_n563), .A3(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n454), .A2(new_n187), .A3(G953), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n561), .A2(new_n277), .A3(new_n562), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n277), .B1(new_n561), .B2(new_n562), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n373), .B1(new_n568), .B2(KEYINPUT14), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n564), .B2(new_n566), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n568), .B(new_n569), .C1(KEYINPUT14), .C2(new_n373), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n572), .B(new_n573), .C1(new_n576), .C2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT89), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n579), .B(new_n578), .C1(new_n574), .C2(new_n575), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n572), .ZN(new_n585));
  INV_X1    g399(.A(new_n573), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n584), .A2(KEYINPUT89), .A3(new_n572), .A4(new_n573), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n583), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n188), .ZN(new_n590));
  INV_X1    g404(.A(G478), .ZN(new_n591));
  OR2_X1    g405(.A1(new_n591), .A2(KEYINPUT15), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n590), .B(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n542), .A2(new_n548), .A3(new_n554), .A4(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n492), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n363), .A2(new_n452), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(G101), .ZN(G3));
  NAND2_X1  g411(.A1(new_n348), .A2(new_n188), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n598), .A2(G472), .B1(new_n349), .B2(new_n348), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n262), .A2(new_n264), .A3(new_n491), .A4(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n589), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT90), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n589), .A2(KEYINPUT90), .A3(new_n602), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT91), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n584), .A2(new_n607), .A3(new_n572), .A4(new_n573), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n587), .A2(KEYINPUT33), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n581), .A2(KEYINPUT91), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n591), .A2(G902), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n605), .A2(new_n606), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT92), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n590), .A2(new_n591), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n603), .A2(new_n604), .B1(new_n610), .B2(new_n609), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT92), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n616), .A2(new_n617), .A3(new_n606), .A4(new_n612), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n614), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n541), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n540), .B1(new_n536), .B2(new_n537), .ZN(new_n621));
  OAI22_X1  g435(.A1(new_n620), .A2(new_n621), .B1(new_n553), .B2(new_n552), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n419), .A2(new_n441), .A3(new_n442), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n442), .B1(new_n419), .B2(new_n441), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n451), .B(new_n548), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n601), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT34), .B(G104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  INV_X1    g444(.A(new_n593), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n542), .A2(new_n631), .A3(new_n554), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n601), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT35), .B(G107), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  INV_X1    g450(.A(new_n599), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n236), .A2(new_n243), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT93), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n255), .A2(KEYINPUT36), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n263), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n637), .B1(new_n643), .B2(new_n262), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n452), .A2(new_n644), .A3(new_n595), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT37), .B(G110), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT94), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n645), .B(new_n647), .ZN(G12));
  AOI21_X1  g462(.A(new_n492), .B1(new_n351), .B2(new_n362), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT95), .B(G900), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n544), .B1(new_n545), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n632), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n451), .B1(new_n624), .B2(new_n625), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n262), .B2(new_n643), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n649), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G128), .ZN(G30));
  NAND2_X1  g470(.A1(new_n348), .A2(new_n349), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT32), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(KEYINPUT67), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n337), .B1(new_n341), .B2(new_n323), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n353), .A2(new_n356), .ZN(new_n662));
  OAI21_X1  g476(.A(KEYINPUT96), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n188), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n661), .A2(new_n662), .A3(KEYINPUT96), .ZN(new_n665));
  OAI21_X1  g479(.A(G472), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT67), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n350), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n660), .A2(new_n666), .A3(new_n668), .A4(new_n361), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n451), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n622), .A2(new_n631), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n651), .B(KEYINPUT39), .Z(new_n674));
  NAND2_X1  g488(.A1(new_n491), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(KEYINPUT40), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n450), .B(KEYINPUT38), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n643), .A2(new_n262), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n673), .A2(new_n676), .A3(new_n677), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G143), .ZN(G45));
  INV_X1    g495(.A(new_n651), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n619), .A2(new_n622), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n649), .A2(new_n654), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT97), .B(G146), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G48));
  NAND3_X1  g500(.A1(new_n362), .A2(new_n660), .A3(new_n668), .ZN(new_n687));
  INV_X1    g501(.A(new_n264), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n258), .A2(new_n188), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n260), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n258), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n688), .B1(new_n692), .B2(new_n189), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n474), .A2(new_n480), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n468), .A2(new_n469), .A3(new_n472), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n484), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI211_X1 g510(.A(KEYINPUT98), .B(G469), .C1(new_n696), .C2(G902), .ZN(new_n697));
  INV_X1    g511(.A(new_n474), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n478), .A2(new_n286), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n475), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n478), .A2(KEYINPUT12), .A3(new_n286), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n698), .A2(new_n702), .A3(new_n695), .ZN(new_n703));
  INV_X1    g517(.A(new_n484), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(KEYINPUT98), .A2(G469), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n188), .A3(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n456), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n697), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n627), .A2(new_n687), .A3(new_n693), .A4(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT41), .B(G113), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT99), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n711), .B(new_n713), .ZN(G15));
  NAND4_X1  g528(.A1(new_n633), .A2(new_n687), .A3(new_n693), .A4(new_n710), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G116), .ZN(G18));
  NOR2_X1   g530(.A1(new_n653), .A2(new_n709), .ZN(new_n717));
  INV_X1    g531(.A(new_n594), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n717), .A2(new_n678), .A3(new_n687), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  NAND2_X1  g534(.A1(new_n357), .A2(new_n337), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n330), .A2(new_n721), .A3(new_n347), .ZN(new_n722));
  XOR2_X1   g536(.A(new_n349), .B(KEYINPUT100), .Z(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT101), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT101), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n722), .A2(new_n726), .A3(new_n723), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT102), .B1(new_n598), .B2(G472), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT102), .ZN(new_n730));
  INV_X1    g544(.A(G472), .ZN(new_n731));
  AOI211_X1 g545(.A(new_n730), .B(new_n731), .C1(new_n348), .C2(new_n188), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n728), .A2(new_n729), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n672), .A2(new_n709), .ZN(new_n734));
  INV_X1    g548(.A(new_n626), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n733), .A2(new_n693), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G122), .ZN(G24));
  NAND4_X1  g551(.A1(new_n717), .A2(new_n733), .A3(new_n683), .A4(new_n678), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  AOI21_X1  g553(.A(new_n671), .B1(new_n445), .B2(new_n446), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n740), .A2(new_n444), .A3(new_n449), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n456), .B1(new_n485), .B2(new_n490), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n683), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT103), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n348), .A2(KEYINPUT32), .A3(new_n349), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n744), .B1(new_n745), .B2(new_n350), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n659), .A2(KEYINPUT103), .A3(new_n361), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n747), .A3(new_n360), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n693), .ZN(new_n749));
  OAI21_X1  g563(.A(KEYINPUT42), .B1(new_n743), .B2(new_n749), .ZN(new_n750));
  AND4_X1   g564(.A1(new_n444), .A2(new_n740), .A3(new_n742), .A4(new_n449), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n623), .A2(KEYINPUT42), .A3(new_n651), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n363), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n284), .ZN(G33));
  NAND4_X1  g569(.A1(new_n751), .A2(new_n687), .A3(new_n693), .A4(new_n652), .ZN(new_n756));
  XNOR2_X1  g570(.A(KEYINPUT104), .B(G134), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(G36));
  INV_X1    g572(.A(new_n622), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT105), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT43), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n619), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n759), .B(new_n619), .C1(new_n760), .C2(KEYINPUT43), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(new_n637), .A3(new_n678), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n486), .A2(new_n483), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n472), .B1(new_n702), .B2(new_n468), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n489), .A2(KEYINPUT45), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n773), .A3(G469), .ZN(new_n774));
  NAND2_X1  g588(.A1(G469), .A2(G902), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT46), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n485), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n774), .A2(KEYINPUT46), .A3(new_n775), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n780), .A2(new_n708), .A3(new_n674), .A4(new_n741), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n781), .B1(new_n766), .B2(new_n767), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n768), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  AOI21_X1  g598(.A(KEYINPUT47), .B1(new_n780), .B2(new_n708), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n786));
  AOI211_X1 g600(.A(new_n786), .B(new_n456), .C1(new_n778), .C2(new_n779), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n683), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n740), .A2(new_n444), .A3(new_n449), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n789), .A2(new_n687), .A3(new_n693), .A4(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n788), .A2(KEYINPUT106), .A3(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT106), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n785), .A2(new_n787), .ZN(new_n794));
  INV_X1    g608(.A(new_n791), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  INV_X1    g612(.A(new_n457), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n693), .A2(new_n451), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT107), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n697), .A2(new_n707), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n762), .B1(KEYINPUT49), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT108), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n670), .B1(KEYINPUT49), .B2(new_n802), .ZN(new_n806));
  OR3_X1    g620(.A1(new_n805), .A2(new_n677), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(G952), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n252), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT50), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n697), .A2(new_n707), .A3(new_n671), .A4(new_n708), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(KEYINPUT112), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n677), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n544), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n763), .B2(new_n764), .ZN(new_n816));
  OR3_X1    g630(.A1(new_n728), .A2(new_n729), .A3(new_n732), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n265), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n810), .B1(new_n814), .B2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n813), .A2(new_n816), .A3(KEYINPUT50), .A4(new_n818), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n819), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n802), .A2(new_n799), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n741), .B(new_n823), .C1(new_n788), .C2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n817), .A2(new_n679), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n790), .A2(new_n709), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n816), .A2(KEYINPUT113), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT113), .B1(new_n816), .B2(new_n827), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n826), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n693), .A2(new_n670), .A3(new_n827), .A4(new_n544), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n619), .A2(new_n622), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n822), .A2(new_n825), .A3(new_n830), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT51), .ZN(new_n835));
  INV_X1    g649(.A(new_n824), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n790), .B1(new_n794), .B2(new_n836), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n837), .A2(new_n823), .B1(new_n831), .B2(new_n832), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n838), .A2(new_n839), .A3(new_n822), .A4(new_n830), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n717), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT114), .B1(new_n819), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n816), .A2(new_n844), .A3(new_n717), .A4(new_n818), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n623), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n543), .B1(new_n831), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT115), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n846), .A2(KEYINPUT115), .A3(new_n848), .ZN(new_n852));
  INV_X1    g666(.A(new_n749), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n853), .B1(new_n828), .B2(new_n829), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT48), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT48), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n856), .B(new_n853), .C1(new_n828), .C2(new_n829), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n851), .A2(new_n852), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n841), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n653), .A2(new_n672), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n742), .A2(new_n682), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n679), .A2(new_n860), .A3(new_n669), .A4(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n655), .A2(new_n684), .A3(new_n738), .A4(new_n862), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT52), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n693), .A2(new_n687), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n595), .A2(new_n451), .A3(new_n450), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n736), .B(new_n719), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n450), .A2(new_n451), .A3(new_n548), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n600), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n623), .A2(KEYINPUT109), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT109), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n619), .A2(new_n871), .A3(new_n622), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n632), .A3(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n750), .A2(new_n753), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n711), .A2(new_n645), .A3(new_n715), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n751), .A2(new_n733), .A3(new_n683), .A4(new_n678), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n542), .A2(new_n593), .A3(new_n554), .A4(new_n682), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n880), .B1(new_n262), .B2(new_n643), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(new_n687), .A3(new_n491), .A4(new_n741), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n756), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n875), .A2(new_n876), .A3(new_n878), .A4(new_n884), .ZN(new_n885));
  XNOR2_X1  g699(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n864), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n869), .A2(new_n873), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n888), .A2(new_n596), .A3(new_n719), .A4(new_n736), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n889), .A2(new_n754), .A3(new_n877), .A4(new_n883), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n684), .A2(new_n862), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n891), .A2(KEYINPUT52), .A3(new_n655), .A4(new_n738), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT52), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n863), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT53), .B1(new_n890), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT54), .B1(new_n887), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n886), .B1(new_n864), .B2(new_n885), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT54), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n890), .A2(new_n895), .A3(KEYINPUT53), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n897), .A2(KEYINPUT111), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT111), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n898), .A2(new_n900), .A3(new_n903), .A4(new_n899), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n859), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT116), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n809), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI211_X1 g721(.A(KEYINPUT116), .B(new_n859), .C1(new_n902), .C2(new_n904), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n807), .B1(new_n907), .B2(new_n908), .ZN(G75));
  AOI21_X1  g723(.A(new_n188), .B1(new_n898), .B2(new_n900), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(G210), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT56), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n414), .A2(new_n418), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n368), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT55), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n911), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n915), .B1(new_n911), .B2(new_n912), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n808), .A2(G953), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT117), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n916), .A2(new_n917), .A3(new_n920), .ZN(G51));
  NAND2_X1  g735(.A1(new_n901), .A2(KEYINPUT118), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT118), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n898), .A2(new_n900), .A3(new_n923), .A4(new_n899), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n898), .A2(new_n900), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n922), .B(new_n924), .C1(new_n899), .C2(new_n925), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n775), .B(KEYINPUT57), .Z(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n705), .ZN(new_n929));
  INV_X1    g743(.A(new_n774), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n910), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n920), .B1(new_n929), .B2(new_n931), .ZN(G54));
  AND2_X1   g746(.A1(KEYINPUT58), .A2(G475), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n910), .A2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n536), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n919), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT119), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n934), .B2(new_n935), .ZN(new_n938));
  AOI211_X1 g752(.A(KEYINPUT119), .B(new_n536), .C1(new_n910), .C2(new_n933), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(G60));
  AND2_X1   g754(.A1(new_n616), .A2(new_n606), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n902), .A2(new_n904), .ZN(new_n943));
  NAND2_X1  g757(.A1(G478), .A2(G902), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT59), .Z(new_n945));
  OAI21_X1  g759(.A(new_n942), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n942), .A2(new_n945), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n920), .B1(new_n926), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n946), .A2(new_n948), .ZN(G63));
  NAND2_X1  g763(.A1(G217), .A2(G902), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT60), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n898), .B2(new_n900), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n641), .A2(new_n642), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(KEYINPUT120), .ZN(new_n955));
  OR2_X1    g769(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n919), .B(new_n956), .C1(new_n952), .C2(new_n258), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT120), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n952), .A2(new_n958), .A3(new_n953), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n955), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n952), .A2(new_n258), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n919), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT121), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n961), .A2(new_n919), .A3(new_n954), .A4(new_n956), .ZN(new_n965));
  AOI22_X1  g779(.A1(new_n960), .A2(new_n964), .B1(KEYINPUT61), .B2(new_n965), .ZN(G66));
  OAI21_X1  g780(.A(G953), .B1(new_n366), .B2(new_n546), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n889), .A2(new_n877), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n968), .B2(G953), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n913), .B1(G898), .B2(new_n252), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G69));
  AOI21_X1  g785(.A(new_n252), .B1(G227), .B2(G900), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n790), .A2(new_n675), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n873), .A2(new_n363), .A3(new_n973), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT123), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n797), .A2(new_n783), .A3(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n655), .A2(new_n684), .A3(new_n738), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n680), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT62), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n978), .A2(new_n981), .A3(new_n680), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n252), .B1(new_n976), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n303), .A2(new_n308), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT122), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(new_n522), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n984), .A2(KEYINPUT124), .A3(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(KEYINPUT124), .B1(new_n984), .B2(new_n987), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI22_X1  g805(.A1(new_n792), .A2(new_n796), .B1(new_n768), .B2(new_n782), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n853), .A2(new_n860), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n780), .A2(new_n708), .A3(new_n674), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n756), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n995), .A2(new_n754), .A3(new_n977), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n252), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT125), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n252), .A2(G900), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(G953), .B1(new_n992), .B2(new_n996), .ZN(new_n1003));
  OAI21_X1  g817(.A(KEYINPUT125), .B1(new_n1003), .B2(new_n1000), .ZN(new_n1004));
  INV_X1    g818(.A(new_n987), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n972), .B1(new_n991), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n990), .ZN(new_n1008));
  AND4_X1   g822(.A1(new_n1006), .A2(new_n1008), .A3(new_n988), .A4(new_n972), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1007), .A2(new_n1009), .ZN(G72));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT63), .Z(new_n1012));
  INV_X1    g826(.A(new_n968), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1012), .B1(new_n997), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n354), .B(KEYINPUT127), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1012), .ZN(new_n1017));
  AOI211_X1 g831(.A(new_n1017), .B(new_n661), .C1(new_n341), .C2(new_n353), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1018), .B1(new_n887), .B2(new_n896), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1016), .A2(new_n919), .A3(new_n1019), .ZN(new_n1020));
  NOR3_X1   g834(.A1(new_n976), .A2(new_n983), .A3(new_n1013), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n661), .B1(new_n1021), .B2(new_n1017), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT126), .ZN(new_n1023));
  OR2_X1    g837(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1020), .B1(new_n1024), .B2(new_n1025), .ZN(G57));
endmodule


