//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G140), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT77), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G227), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n189), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT1), .B1(new_n193), .B2(G146), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(G146), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  OAI211_X1 g011(.A(G128), .B(new_n194), .C1(new_n195), .C2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n193), .A2(G146), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n199), .B(new_n200), .C1(KEYINPUT1), .C2(new_n201), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n198), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT3), .B1(new_n204), .B2(G107), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  INV_X1    g020(.A(G107), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G104), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT79), .B1(new_n207), .B2(G104), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT79), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(new_n204), .A3(G107), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n209), .A2(new_n210), .A3(new_n211), .A4(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n204), .A2(G107), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n207), .A2(G104), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n210), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n203), .A2(new_n214), .A3(KEYINPUT10), .A4(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT10), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n211), .A2(new_n205), .A3(new_n213), .A4(new_n208), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n218), .B1(new_n221), .B2(G101), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n198), .A2(new_n202), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n220), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n221), .A2(G101), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT4), .B1(new_n221), .B2(G101), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT4), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n221), .A2(new_n228), .A3(G101), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT0), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(new_n201), .ZN(new_n231));
  NOR2_X1   g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  OAI22_X1  g046(.A1(new_n195), .A2(new_n197), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n199), .B(new_n200), .C1(new_n230), .C2(new_n201), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n229), .A2(new_n235), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n219), .B(new_n224), .C1(new_n227), .C2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT11), .ZN(new_n238));
  INV_X1    g052(.A(G134), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n238), .B1(new_n239), .B2(G137), .ZN(new_n240));
  INV_X1    g054(.A(G137), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(KEYINPUT11), .A3(G134), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(G137), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G131), .ZN(new_n245));
  INV_X1    g059(.A(G131), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n240), .A2(new_n242), .A3(new_n246), .A4(new_n243), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n237), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n221), .A2(G101), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n214), .A2(KEYINPUT4), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(new_n235), .A3(new_n229), .ZN(new_n252));
  INV_X1    g066(.A(new_n248), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n252), .A2(new_n253), .A3(new_n219), .A4(new_n224), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n192), .B1(new_n249), .B2(new_n254), .ZN(new_n255));
  OR2_X1    g069(.A1(new_n255), .A2(KEYINPUT82), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n192), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT81), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n254), .A2(KEYINPUT81), .A3(new_n192), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n222), .B(new_n223), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n248), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT12), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n261), .A2(KEYINPUT12), .A3(new_n248), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n259), .A2(new_n260), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n255), .A2(KEYINPUT82), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n256), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G469), .ZN(new_n270));
  INV_X1    g084(.A(G902), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n249), .A2(new_n254), .A3(new_n192), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n266), .A2(KEYINPUT80), .A3(new_n254), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n192), .B(KEYINPUT78), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT80), .B1(new_n266), .B2(new_n254), .ZN(new_n277));
  OAI211_X1 g091(.A(G469), .B(new_n273), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(G469), .A2(G902), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n272), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT9), .B(G234), .ZN(new_n281));
  OAI21_X1  g095(.A(G221), .B1(new_n281), .B2(G902), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G140), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G125), .ZN(new_n285));
  INV_X1    g099(.A(G125), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G140), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n196), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(G146), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(KEYINPUT88), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G237), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n190), .A3(G214), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n294), .B(new_n193), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT18), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(new_n246), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n291), .A2(KEYINPUT88), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n292), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n294), .B(G143), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n301), .B(KEYINPUT89), .C1(new_n296), .C2(new_n246), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT89), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n303), .B1(new_n295), .B2(new_n297), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n285), .A2(new_n287), .A3(KEYINPUT16), .ZN(new_n307));
  OR3_X1    g121(.A1(new_n286), .A2(KEYINPUT16), .A3(G140), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n307), .A2(G146), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(G146), .B1(new_n307), .B2(new_n308), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n295), .A2(KEYINPUT17), .A3(G131), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n295), .A2(G131), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n301), .A2(new_n246), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n311), .B(new_n312), .C1(new_n315), .C2(KEYINPUT17), .ZN(new_n316));
  XNOR2_X1  g130(.A(G113), .B(G122), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(new_n204), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n306), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n318), .B1(new_n306), .B2(new_n316), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n271), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G475), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n289), .A2(KEYINPUT90), .A3(KEYINPUT19), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n324), .B1(new_n289), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n309), .B1(new_n326), .B2(new_n196), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n315), .A2(new_n327), .B1(new_n300), .B2(new_n305), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n319), .B1(new_n328), .B2(new_n318), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT20), .ZN(new_n330));
  NOR2_X1   g144(.A1(G475), .A2(G902), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n330), .B1(new_n329), .B2(new_n331), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n323), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G478), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(KEYINPUT15), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n193), .A2(G128), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n201), .A2(G143), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(new_n239), .ZN(new_n342));
  INV_X1    g156(.A(G116), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G122), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(G122), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n344), .B1(new_n345), .B2(KEYINPUT14), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(KEYINPUT14), .B2(new_n344), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G107), .ZN(new_n348));
  XNOR2_X1  g162(.A(G116), .B(G122), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n207), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n342), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n339), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(KEYINPUT13), .B2(new_n340), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n352), .A2(KEYINPUT13), .ZN(new_n354));
  OAI21_X1  g168(.A(G134), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n341), .A2(new_n239), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n349), .B(new_n207), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n351), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n281), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(G217), .A3(new_n190), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n361), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n351), .A2(new_n358), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n338), .B1(new_n365), .B2(new_n271), .ZN(new_n366));
  AOI211_X1 g180(.A(G902), .B(new_n337), .C1(new_n362), .C2(new_n364), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G952), .ZN(new_n370));
  AOI211_X1 g184(.A(G953), .B(new_n370), .C1(G234), .C2(G237), .ZN(new_n371));
  AOI211_X1 g185(.A(new_n271), .B(new_n190), .C1(G234), .C2(G237), .ZN(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT21), .B(G898), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n335), .A2(new_n369), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n283), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(G110), .B(G122), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(G116), .B(G119), .ZN(new_n379));
  NAND2_X1  g193(.A1(KEYINPUT2), .A2(G113), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT66), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT66), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(KEYINPUT2), .A3(G113), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  OR2_X1    g198(.A1(KEYINPUT2), .A2(G113), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n379), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT67), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n381), .A2(new_n383), .ZN(new_n388));
  INV_X1    g202(.A(G119), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G116), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n343), .A2(G119), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n385), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n387), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n384), .A2(KEYINPUT67), .A3(new_n379), .A4(new_n385), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n386), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n229), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n227), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT5), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(new_n389), .A3(G116), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G113), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n400), .B1(KEYINPUT5), .B2(new_n379), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n401), .B1(new_n393), .B2(new_n394), .ZN(new_n402));
  INV_X1    g216(.A(new_n222), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n378), .B1(new_n397), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n395), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(new_n251), .A3(new_n229), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n404), .A3(new_n377), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n406), .A2(KEYINPUT6), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G224), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(G953), .ZN(new_n412));
  AOI21_X1  g226(.A(G125), .B1(new_n198), .B2(new_n202), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT83), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n233), .A2(G125), .A3(new_n234), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n233), .A2(KEYINPUT83), .A3(G125), .A4(new_n234), .ZN(new_n417));
  AOI21_X1  g231(.A(KEYINPUT84), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n414), .ZN(new_n419));
  INV_X1    g233(.A(new_n413), .ZN(new_n420));
  AND4_X1   g234(.A1(KEYINPUT84), .A2(new_n419), .A3(new_n420), .A4(new_n417), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n412), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n419), .A2(new_n420), .A3(new_n417), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT84), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n416), .A2(KEYINPUT84), .A3(new_n417), .ZN(new_n426));
  INV_X1    g240(.A(new_n412), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT6), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n430), .B(new_n378), .C1(new_n397), .C2(new_n405), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n410), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n427), .A2(KEYINPUT7), .ZN(new_n433));
  INV_X1    g247(.A(new_n415), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n433), .B1(new_n434), .B2(new_n413), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n435), .B1(new_n423), .B2(new_n433), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n395), .A2(new_n396), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n437), .A2(new_n251), .B1(new_n403), .B2(new_n402), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n436), .B1(new_n438), .B2(new_n377), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n377), .B(KEYINPUT8), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT85), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n402), .B2(new_n403), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n404), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n402), .A2(new_n403), .A3(new_n441), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n440), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(G902), .B1(new_n439), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n432), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G210), .B1(G237), .B2(G902), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT86), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n448), .B1(new_n432), .B2(new_n446), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT86), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n432), .A2(new_n446), .A3(new_n448), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT87), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT87), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n432), .A2(new_n446), .A3(new_n457), .A4(new_n448), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n452), .A2(new_n454), .A3(new_n456), .A4(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(G214), .B1(G237), .B2(G902), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n187), .B1(new_n376), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G234), .ZN(new_n463));
  OAI21_X1  g277(.A(G217), .B1(new_n463), .B2(G902), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(KEYINPUT71), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT25), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT23), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n468), .B1(new_n389), .B2(G128), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n389), .A2(G128), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(G119), .B(G128), .ZN(new_n473));
  INV_X1    g287(.A(G110), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT24), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT24), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(G110), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n472), .A2(G110), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n479), .B1(new_n309), .B2(new_n310), .ZN(new_n480));
  OAI22_X1  g294(.A1(new_n472), .A2(G110), .B1(new_n473), .B2(new_n478), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n307), .A2(new_n308), .A3(G146), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n482), .A3(new_n290), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT73), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(KEYINPUT22), .B(G137), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT72), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n489), .B(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n480), .A2(new_n483), .A3(KEYINPUT73), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n486), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n489), .B(new_n490), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n485), .A3(new_n484), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT74), .B1(new_n497), .B2(new_n271), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT74), .ZN(new_n499));
  AOI211_X1 g313(.A(new_n499), .B(G902), .C1(new_n494), .C2(new_n496), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n467), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(KEYINPUT25), .A3(new_n271), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT75), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n503), .B(new_n467), .C1(new_n498), .C2(new_n500), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n466), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n466), .A2(new_n271), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT76), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n497), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT32), .ZN(new_n514));
  NOR2_X1   g328(.A1(G472), .A2(G902), .ZN(new_n515));
  XOR2_X1   g329(.A(new_n515), .B(KEYINPUT70), .Z(new_n516));
  INV_X1    g330(.A(G210), .ZN(new_n517));
  NOR3_X1   g331(.A1(new_n517), .A2(G237), .A3(G953), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT27), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT26), .B(G101), .ZN(new_n520));
  XOR2_X1   g334(.A(new_n519), .B(new_n520), .Z(new_n521));
  NOR2_X1   g335(.A1(new_n239), .A2(G137), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n241), .A2(G134), .ZN(new_n523));
  OAI21_X1  g337(.A(G131), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT68), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n247), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n525), .B1(new_n247), .B2(new_n524), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n203), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n248), .A2(new_n235), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n395), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n245), .A2(new_n247), .B1(new_n233), .B2(new_n234), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT64), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n247), .A2(new_n524), .ZN(new_n534));
  OAI22_X1  g348(.A1(new_n532), .A2(new_n533), .B1(new_n223), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n529), .A2(KEYINPUT64), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n407), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT28), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT28), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n531), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n521), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n528), .A2(new_n529), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT30), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT69), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT69), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n528), .A2(new_n546), .A3(KEYINPUT30), .A4(new_n529), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n544), .B1(new_n535), .B2(new_n536), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT65), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT65), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n551), .B(new_n544), .C1(new_n535), .C2(new_n536), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n548), .A2(new_n550), .A3(new_n407), .A4(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(new_n531), .A3(new_n521), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n542), .B1(new_n554), .B2(KEYINPUT31), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT31), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n553), .A2(new_n556), .A3(new_n531), .A4(new_n521), .ZN(new_n557));
  AOI211_X1 g371(.A(new_n514), .B(new_n516), .C1(new_n555), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(KEYINPUT31), .ZN(new_n559));
  INV_X1    g373(.A(new_n542), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n516), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT32), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n543), .A2(new_n407), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n543), .A2(new_n407), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT28), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n568), .A2(new_n541), .ZN(new_n569));
  INV_X1    g383(.A(new_n521), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT29), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(G902), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n539), .A2(new_n521), .A3(new_n541), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n571), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n521), .B1(new_n553), .B2(new_n531), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n573), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(G472), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n513), .B1(new_n564), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n461), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n580), .A2(KEYINPUT91), .A3(new_n375), .A4(new_n283), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n462), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(G101), .ZN(G3));
  NAND2_X1  g397(.A1(new_n561), .A2(new_n562), .ZN(new_n584));
  AOI21_X1  g398(.A(G902), .B1(new_n555), .B2(new_n557), .ZN(new_n585));
  INV_X1    g399(.A(G472), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n280), .A2(new_n282), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n513), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n460), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n450), .B2(new_n455), .ZN(new_n591));
  INV_X1    g405(.A(new_n374), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n365), .A2(new_n271), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(G478), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT33), .B1(new_n363), .B2(KEYINPUT92), .ZN(new_n596));
  OR2_X1    g410(.A1(new_n365), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n365), .A2(new_n596), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n597), .A2(new_n271), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n595), .B1(new_n599), .B2(G478), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n335), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n593), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n589), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT34), .B(G104), .Z(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G6));
  OAI211_X1 g419(.A(new_n369), .B(new_n323), .C1(new_n334), .C2(new_n333), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n593), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n589), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT35), .B(G107), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G9));
  NOR2_X1   g424(.A1(new_n492), .A2(KEYINPUT36), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT94), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n484), .B(KEYINPUT93), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n510), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n507), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n587), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n462), .A2(new_n581), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT37), .B(G110), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G12));
  NAND2_X1  g434(.A1(new_n584), .A2(new_n514), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n516), .B1(new_n555), .B2(new_n557), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(KEYINPUT32), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(new_n623), .A3(new_n578), .ZN(new_n624));
  INV_X1    g438(.A(new_n591), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n616), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT95), .ZN(new_n628));
  INV_X1    g442(.A(G900), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n372), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n371), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n628), .B1(new_n606), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n334), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n635), .A2(new_n332), .B1(G475), .B2(new_n322), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n636), .A2(KEYINPUT95), .A3(new_n369), .A4(new_n632), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n638), .A2(new_n283), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n627), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G128), .ZN(G30));
  XOR2_X1   g455(.A(new_n459), .B(KEYINPUT38), .Z(new_n642));
  NOR2_X1   g456(.A1(new_n636), .A2(new_n368), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n616), .A2(new_n460), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n570), .B1(new_n566), .B2(new_n567), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n554), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n586), .B1(new_n647), .B2(new_n271), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n564), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n632), .B(KEYINPUT39), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n283), .A2(new_n651), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n645), .A2(new_n650), .A3(new_n653), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G143), .ZN(G45));
  NOR2_X1   g470(.A1(new_n601), .A2(new_n633), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n588), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n627), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G146), .ZN(G48));
  AOI21_X1  g475(.A(new_n507), .B1(new_n497), .B2(new_n511), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n269), .A2(new_n271), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(KEYINPUT96), .A3(G469), .ZN(new_n664));
  NAND2_X1  g478(.A1(KEYINPUT96), .A2(G469), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n269), .A2(new_n271), .A3(new_n665), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n664), .A2(new_n282), .A3(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n624), .A2(new_n662), .A3(new_n602), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT41), .B(G113), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G15));
  NAND4_X1  g484(.A1(new_n624), .A2(new_n607), .A3(new_n662), .A4(new_n667), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G116), .ZN(G18));
  NAND4_X1  g486(.A1(new_n624), .A2(new_n626), .A3(new_n375), .A4(new_n667), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G119), .ZN(G21));
  AND4_X1   g488(.A1(new_n592), .A2(new_n664), .A3(new_n282), .A4(new_n666), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n561), .A2(new_n271), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT98), .B(G472), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n568), .A2(KEYINPUT97), .A3(new_n541), .ZN(new_n679));
  AOI21_X1  g493(.A(KEYINPUT97), .B1(new_n568), .B2(new_n541), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n570), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n559), .A3(new_n557), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n676), .A2(new_n678), .B1(new_n562), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n643), .A2(new_n591), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n675), .A2(new_n662), .A3(new_n683), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G122), .ZN(G24));
  OR2_X1    g501(.A1(new_n507), .A2(new_n615), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n683), .A2(new_n688), .A3(new_n657), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n667), .A2(new_n591), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT99), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G125), .ZN(G27));
  OAI21_X1  g508(.A(KEYINPUT101), .B1(new_n459), .B2(new_n590), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n266), .A2(new_n254), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT80), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n274), .A3(new_n275), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n273), .B(KEYINPUT100), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n272), .B(new_n279), .C1(new_n701), .C2(new_n270), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n453), .B(new_n451), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n456), .A2(new_n458), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT101), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n703), .A2(new_n704), .A3(new_n705), .A4(new_n460), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n695), .A2(new_n282), .A3(new_n702), .A4(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n578), .B1(new_n622), .B2(KEYINPUT32), .ZN(new_n709));
  AOI21_X1  g523(.A(KEYINPUT102), .B1(new_n622), .B2(KEYINPUT32), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n558), .A2(KEYINPUT102), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n513), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n708), .A2(new_n713), .A3(new_n657), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT42), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n624), .A2(new_n662), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n707), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(new_n718), .A3(new_n657), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n246), .ZN(G33));
  AND3_X1   g535(.A1(new_n695), .A2(new_n282), .A3(new_n706), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n722), .A2(new_n579), .A3(new_n638), .A4(new_n702), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G134), .ZN(G36));
  NAND2_X1  g538(.A1(new_n699), .A2(new_n273), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n270), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT103), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n699), .A2(new_n700), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n728), .B1(new_n729), .B2(KEYINPUT45), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n701), .A2(KEYINPUT103), .A3(new_n726), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n727), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(KEYINPUT46), .A3(new_n279), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n272), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT46), .B1(new_n732), .B2(new_n279), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n282), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n636), .A2(new_n600), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n738), .A2(KEYINPUT43), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(KEYINPUT43), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n587), .A2(new_n688), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(KEYINPUT44), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n695), .A2(new_n706), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n737), .A2(new_n651), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT104), .B(G137), .Z(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G39));
  INV_X1    g560(.A(KEYINPUT47), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n736), .A2(new_n747), .ZN(new_n748));
  OAI211_X1 g562(.A(KEYINPUT47), .B(new_n282), .C1(new_n734), .C2(new_n735), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n743), .ZN(new_n751));
  NOR4_X1   g565(.A1(new_n751), .A2(new_n662), .A3(new_n624), .A4(new_n658), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G140), .ZN(G42));
  INV_X1    g568(.A(KEYINPUT54), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n756));
  INV_X1    g570(.A(new_n366), .ZN(new_n757));
  INV_X1    g571(.A(new_n367), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT106), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g574(.A(KEYINPUT106), .B1(new_n366), .B2(new_n367), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n761), .A3(new_n632), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n335), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n763), .B1(new_n507), .B2(new_n615), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n588), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n743), .A2(new_n756), .A3(new_n624), .A4(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n765), .A2(new_n624), .A3(new_n706), .A4(new_n695), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT108), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n682), .A2(new_n562), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n770), .B1(new_n585), .B2(new_n677), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n771), .A2(new_n658), .A3(new_n616), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n708), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n723), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT109), .B1(new_n769), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n707), .A2(new_n658), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n718), .B1(new_n776), .B2(new_n713), .ZN(new_n777));
  NOR4_X1   g591(.A1(new_n707), .A2(new_n716), .A3(KEYINPUT42), .A4(new_n658), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n668), .A2(new_n673), .A3(new_n671), .A4(new_n686), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n766), .A2(new_n768), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT109), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n781), .A2(new_n782), .A3(new_n723), .A4(new_n773), .ZN(new_n783));
  XOR2_X1   g597(.A(new_n601), .B(KEYINPUT105), .Z(new_n784));
  NAND2_X1  g598(.A1(new_n760), .A2(new_n761), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n636), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT107), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n374), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n580), .A3(new_n589), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n582), .A2(new_n618), .A3(new_n789), .ZN(new_n790));
  AND4_X1   g604(.A1(new_n775), .A2(new_n780), .A3(new_n783), .A4(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n282), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n633), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n616), .A2(new_n702), .A3(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n616), .A2(KEYINPUT110), .A3(new_n702), .A4(new_n793), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n684), .B1(new_n564), .B2(new_n649), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n627), .B1(new_n639), .B2(new_n659), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n693), .A2(KEYINPUT52), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n690), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n692), .B1(new_n803), .B2(new_n772), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n689), .A2(new_n690), .A3(KEYINPUT99), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n801), .B(new_n800), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n802), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n791), .A2(KEYINPUT53), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n775), .A2(new_n780), .A3(new_n783), .A4(new_n790), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n806), .B(KEYINPUT52), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n755), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT111), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n783), .A2(new_n790), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n717), .A2(new_n638), .B1(new_n708), .B2(new_n772), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n782), .B1(new_n818), .B2(new_n781), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n816), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n775), .A2(KEYINPUT111), .A3(new_n783), .A4(new_n790), .ZN(new_n821));
  AND4_X1   g635(.A1(new_n668), .A2(new_n673), .A3(new_n671), .A4(new_n686), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n715), .A2(KEYINPUT53), .A3(new_n719), .A4(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n808), .B2(new_n802), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n820), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  XOR2_X1   g639(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n826));
  AND3_X1   g640(.A1(new_n825), .A2(new_n814), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n815), .B1(new_n827), .B2(KEYINPUT113), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT114), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n825), .A2(new_n814), .A3(new_n826), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT113), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n739), .A2(new_n371), .A3(new_n740), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n771), .A2(new_n513), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n663), .B(new_n665), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n837), .A2(new_n792), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n743), .B(new_n836), .C1(new_n750), .C2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n667), .A2(new_n590), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n836), .A2(KEYINPUT50), .A3(new_n642), .A4(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT50), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n642), .A2(new_n840), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n842), .B1(new_n843), .B2(new_n835), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n722), .A2(new_n837), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(new_n688), .A3(new_n683), .A4(new_n833), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n650), .A2(new_n513), .A3(new_n631), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n335), .A2(new_n600), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n846), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n845), .A2(new_n847), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n839), .A2(KEYINPUT51), .A3(new_n851), .ZN(new_n852));
  AOI211_X1 g666(.A(new_n370), .B(G953), .C1(new_n836), .C2(new_n803), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n846), .A2(new_n848), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(new_n854), .B2(new_n601), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n846), .A2(new_n713), .A3(new_n833), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n856), .A2(KEYINPUT48), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(KEYINPUT48), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT51), .B1(new_n839), .B2(new_n851), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n828), .A2(new_n829), .A3(new_n832), .A4(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n825), .A2(new_n814), .A3(KEYINPUT113), .A4(new_n826), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT53), .B1(new_n791), .B2(new_n809), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n812), .A2(new_n813), .A3(new_n811), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT54), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n832), .A2(new_n864), .A3(new_n867), .A4(new_n862), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT114), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n370), .A2(new_n190), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n863), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n837), .B(KEYINPUT49), .ZN(new_n872));
  INV_X1    g686(.A(new_n650), .ZN(new_n873));
  NOR4_X1   g687(.A1(new_n513), .A2(new_n590), .A3(new_n792), .A4(new_n738), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n642), .A2(new_n872), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n871), .A2(new_n875), .ZN(G75));
  INV_X1    g690(.A(KEYINPUT56), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n271), .B1(new_n825), .B2(new_n814), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n877), .B1(new_n879), .B2(new_n517), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n410), .A2(new_n431), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(new_n429), .Z(new_n882));
  XOR2_X1   g696(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n883));
  XNOR2_X1  g697(.A(new_n882), .B(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n880), .A2(new_n885), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n190), .A2(G952), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(G51));
  NAND2_X1  g703(.A1(new_n830), .A2(KEYINPUT116), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT116), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n825), .A2(new_n814), .A3(new_n891), .A4(new_n826), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n825), .A2(new_n814), .ZN(new_n893));
  INV_X1    g707(.A(new_n826), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n890), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n279), .B(KEYINPUT57), .Z(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n269), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n732), .B(KEYINPUT117), .Z(new_n900));
  NAND2_X1  g714(.A1(new_n878), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n888), .B1(new_n899), .B2(new_n901), .ZN(G54));
  INV_X1    g716(.A(new_n329), .ZN(new_n903));
  NAND2_X1  g717(.A1(KEYINPUT58), .A2(G475), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n903), .B1(new_n879), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n888), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n878), .A2(KEYINPUT58), .A3(G475), .A4(new_n329), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT118), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT118), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n905), .A2(new_n910), .A3(new_n906), .A4(new_n907), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n909), .A2(new_n911), .ZN(G60));
  AND2_X1   g726(.A1(new_n597), .A2(new_n598), .ZN(new_n913));
  NAND2_X1  g727(.A1(G478), .A2(G902), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT59), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n896), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n832), .A2(new_n864), .A3(new_n867), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n913), .B1(new_n917), .B2(new_n915), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n916), .A2(new_n918), .A3(new_n888), .ZN(G63));
  NAND2_X1  g733(.A1(G217), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT60), .Z(new_n921));
  NAND2_X1  g735(.A1(new_n893), .A2(new_n921), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n614), .B(KEYINPUT120), .Z(new_n923));
  OAI21_X1  g737(.A(new_n906), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n497), .B(KEYINPUT121), .Z(new_n927));
  AOI21_X1  g741(.A(KEYINPUT122), .B1(new_n922), .B2(new_n927), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n922), .A2(KEYINPUT122), .A3(new_n927), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  XOR2_X1   g744(.A(KEYINPUT119), .B(KEYINPUT61), .Z(new_n931));
  AND2_X1   g745(.A1(new_n922), .A2(new_n927), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n931), .B1(new_n932), .B2(new_n924), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n930), .A2(new_n933), .ZN(G66));
  NOR3_X1   g748(.A1(new_n373), .A2(new_n411), .A3(new_n190), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n790), .A2(new_n822), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(new_n190), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n881), .B1(G898), .B2(new_n190), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G69));
  NAND3_X1  g753(.A1(new_n548), .A2(new_n550), .A3(new_n552), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(new_n326), .Z(new_n941));
  OR2_X1    g755(.A1(new_n941), .A2(G953), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT123), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n652), .B1(new_n784), .B2(new_n787), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n579), .A3(new_n743), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n744), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n944), .B1(new_n744), .B2(new_n946), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n753), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n693), .A2(new_n655), .A3(new_n801), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT62), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n943), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n949), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n947), .ZN(new_n955));
  INV_X1    g769(.A(new_n952), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n955), .A2(new_n956), .A3(KEYINPUT124), .A4(new_n753), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n942), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n941), .B1(G900), .B2(new_n190), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n744), .A2(new_n723), .ZN(new_n960));
  INV_X1    g774(.A(new_n651), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n713), .A2(new_n685), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n736), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(new_n750), .B2(new_n752), .ZN(new_n964));
  AND4_X1   g778(.A1(new_n693), .A2(new_n715), .A3(new_n719), .A4(new_n801), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n960), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n959), .B1(new_n966), .B2(new_n190), .ZN(new_n967));
  OAI21_X1  g781(.A(KEYINPUT126), .B1(new_n958), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(G227), .ZN(new_n969));
  OAI21_X1  g783(.A(G953), .B1(new_n969), .B2(new_n629), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT125), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n971), .ZN(new_n973));
  OAI211_X1 g787(.A(KEYINPUT126), .B(new_n973), .C1(new_n958), .C2(new_n967), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(G72));
  NAND2_X1  g789(.A1(new_n553), .A2(new_n531), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n521), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n953), .A2(new_n936), .A3(new_n957), .ZN(new_n978));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  AOI21_X1  g794(.A(new_n977), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n976), .A2(new_n521), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n960), .A2(new_n936), .A3(new_n964), .A4(new_n965), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT127), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n983), .A2(new_n984), .A3(new_n980), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n984), .B1(new_n983), .B2(new_n980), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n982), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n906), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n976), .A2(new_n570), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n980), .B1(new_n989), .B2(new_n576), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n990), .B1(new_n810), .B2(new_n814), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n981), .A2(new_n988), .A3(new_n991), .ZN(G57));
endmodule


