

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594;

  NOR2_X1 U325 ( .A1(n471), .A2(n566), .ZN(n593) );
  NOR2_X1 U326 ( .A1(n585), .A2(n526), .ZN(n335) );
  NAND2_X1 U327 ( .A1(n548), .A2(n551), .ZN(n486) );
  XNOR2_X2 U328 ( .A(n333), .B(n332), .ZN(n589) );
  XNOR2_X1 U329 ( .A(n464), .B(KEYINPUT123), .ZN(n581) );
  XNOR2_X1 U330 ( .A(n336), .B(KEYINPUT81), .ZN(n389) );
  XNOR2_X1 U331 ( .A(G36GAT), .B(G190GAT), .ZN(n336) );
  XNOR2_X1 U332 ( .A(G176GAT), .B(G204GAT), .ZN(n315) );
  XOR2_X1 U333 ( .A(n580), .B(KEYINPUT36), .Z(n492) );
  INV_X1 U334 ( .A(KEYINPUT37), .ZN(n493) );
  XOR2_X1 U335 ( .A(n352), .B(n351), .Z(n580) );
  XOR2_X1 U336 ( .A(n399), .B(n398), .Z(n540) );
  OR2_X1 U337 ( .A1(n371), .A2(n370), .ZN(n372) );
  INV_X1 U338 ( .A(KEYINPUT101), .ZN(n386) );
  XNOR2_X1 U339 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U340 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U341 ( .A(n340), .B(n339), .ZN(n342) );
  XNOR2_X1 U342 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U343 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U344 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U345 ( .A(n316), .B(n315), .ZN(n383) );
  XNOR2_X1 U346 ( .A(n327), .B(n326), .ZN(n333) );
  XNOR2_X1 U347 ( .A(n496), .B(n495), .ZN(n537) );
  INV_X1 U348 ( .A(G218GAT), .ZN(n472) );
  XNOR2_X1 U349 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U350 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U351 ( .A(n500), .B(G29GAT), .ZN(n501) );
  XNOR2_X1 U352 ( .A(n475), .B(n474), .ZN(G1355GAT) );
  XNOR2_X1 U353 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  XOR2_X1 U354 ( .A(KEYINPUT68), .B(G8GAT), .Z(n294) );
  XNOR2_X1 U355 ( .A(G169GAT), .B(G15GAT), .ZN(n293) );
  XNOR2_X1 U356 ( .A(n294), .B(n293), .ZN(n310) );
  XOR2_X1 U357 ( .A(G113GAT), .B(G141GAT), .Z(n296) );
  XNOR2_X1 U358 ( .A(G197GAT), .B(G22GAT), .ZN(n295) );
  XNOR2_X1 U359 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U360 ( .A(n297), .B(G50GAT), .Z(n299) );
  XOR2_X1 U361 ( .A(G1GAT), .B(KEYINPUT70), .Z(n354) );
  XNOR2_X1 U362 ( .A(n354), .B(G36GAT), .ZN(n298) );
  XNOR2_X1 U363 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U364 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n301) );
  NAND2_X1 U365 ( .A1(G229GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U366 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U367 ( .A(n303), .B(n302), .Z(n308) );
  XOR2_X1 U368 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n305) );
  XNOR2_X1 U369 ( .A(G43GAT), .B(G29GAT), .ZN(n304) );
  XNOR2_X1 U370 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U371 ( .A(KEYINPUT7), .B(n306), .Z(n350) );
  XNOR2_X1 U372 ( .A(n350), .B(KEYINPUT29), .ZN(n307) );
  XNOR2_X1 U373 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U374 ( .A(n310), .B(n309), .ZN(n585) );
  INV_X1 U375 ( .A(G64GAT), .ZN(n311) );
  NAND2_X1 U376 ( .A1(n311), .A2(KEYINPUT74), .ZN(n314) );
  INV_X1 U377 ( .A(KEYINPUT74), .ZN(n312) );
  NAND2_X1 U378 ( .A1(G64GAT), .A2(n312), .ZN(n313) );
  NAND2_X1 U379 ( .A1(n314), .A2(n313), .ZN(n316) );
  XOR2_X1 U380 ( .A(G120GAT), .B(G71GAT), .Z(n446) );
  XNOR2_X1 U381 ( .A(n383), .B(n446), .ZN(n318) );
  AND2_X1 U382 ( .A1(G230GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U383 ( .A(n318), .B(n317), .ZN(n319) );
  NAND2_X1 U384 ( .A1(n319), .A2(KEYINPUT75), .ZN(n321) );
  OR2_X1 U385 ( .A1(n319), .A2(KEYINPUT75), .ZN(n320) );
  NAND2_X1 U386 ( .A1(n321), .A2(n320), .ZN(n327) );
  XOR2_X1 U387 ( .A(G57GAT), .B(KEYINPUT13), .Z(n353) );
  XOR2_X1 U388 ( .A(n353), .B(KEYINPUT33), .Z(n325) );
  XOR2_X1 U389 ( .A(KEYINPUT73), .B(KEYINPUT31), .Z(n323) );
  XNOR2_X1 U390 ( .A(KEYINPUT76), .B(KEYINPUT32), .ZN(n322) );
  XOR2_X1 U391 ( .A(n323), .B(n322), .Z(n324) );
  XOR2_X1 U392 ( .A(G78GAT), .B(G148GAT), .Z(n329) );
  XNOR2_X1 U393 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n328) );
  XNOR2_X1 U394 ( .A(n329), .B(n328), .ZN(n429) );
  XOR2_X1 U395 ( .A(G92GAT), .B(KEYINPUT72), .Z(n331) );
  XNOR2_X1 U396 ( .A(G99GAT), .B(G85GAT), .ZN(n330) );
  XNOR2_X1 U397 ( .A(n331), .B(n330), .ZN(n338) );
  XNOR2_X1 U398 ( .A(n429), .B(n338), .ZN(n332) );
  XOR2_X1 U399 ( .A(KEYINPUT41), .B(n589), .Z(n569) );
  INV_X1 U400 ( .A(n569), .ZN(n526) );
  XNOR2_X1 U401 ( .A(KEYINPUT46), .B(KEYINPUT116), .ZN(n334) );
  XNOR2_X1 U402 ( .A(n335), .B(n334), .ZN(n371) );
  XOR2_X1 U403 ( .A(G106GAT), .B(n389), .Z(n340) );
  NAND2_X1 U404 ( .A1(G232GAT), .A2(G233GAT), .ZN(n337) );
  XOR2_X1 U405 ( .A(G50GAT), .B(G162GAT), .Z(n437) );
  XOR2_X1 U406 ( .A(G134GAT), .B(KEYINPUT79), .Z(n410) );
  XOR2_X1 U407 ( .A(n437), .B(n410), .Z(n341) );
  XNOR2_X1 U408 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U409 ( .A(KEYINPUT10), .B(KEYINPUT82), .Z(n344) );
  XNOR2_X1 U410 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n343) );
  XOR2_X1 U411 ( .A(n344), .B(n343), .Z(n345) );
  XNOR2_X1 U412 ( .A(n346), .B(n345), .ZN(n352) );
  XOR2_X1 U413 ( .A(KEYINPUT66), .B(KEYINPUT80), .Z(n348) );
  XNOR2_X1 U414 ( .A(KEYINPUT78), .B(KEYINPUT11), .ZN(n347) );
  XNOR2_X1 U415 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U416 ( .A(n350), .B(n349), .ZN(n351) );
  INV_X1 U417 ( .A(n580), .ZN(n562) );
  XOR2_X1 U418 ( .A(G22GAT), .B(G155GAT), .Z(n436) );
  XOR2_X1 U419 ( .A(n353), .B(n436), .Z(n356) );
  XOR2_X1 U420 ( .A(G15GAT), .B(G127GAT), .Z(n447) );
  XNOR2_X1 U421 ( .A(n354), .B(n447), .ZN(n355) );
  XNOR2_X1 U422 ( .A(n356), .B(n355), .ZN(n361) );
  XNOR2_X1 U423 ( .A(G8GAT), .B(G183GAT), .ZN(n357) );
  XNOR2_X1 U424 ( .A(n357), .B(KEYINPUT83), .ZN(n394) );
  XOR2_X1 U425 ( .A(KEYINPUT85), .B(n394), .Z(n359) );
  NAND2_X1 U426 ( .A1(G231GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U427 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U428 ( .A(n361), .B(n360), .Z(n369) );
  XOR2_X1 U429 ( .A(G64GAT), .B(G78GAT), .Z(n363) );
  XNOR2_X1 U430 ( .A(G71GAT), .B(G211GAT), .ZN(n362) );
  XNOR2_X1 U431 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U432 ( .A(KEYINPUT84), .B(KEYINPUT14), .Z(n365) );
  XNOR2_X1 U433 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n364) );
  XNOR2_X1 U434 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U435 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U436 ( .A(n369), .B(n368), .Z(n558) );
  NAND2_X1 U437 ( .A1(n562), .A2(n558), .ZN(n370) );
  XNOR2_X1 U438 ( .A(KEYINPUT117), .B(n372), .ZN(n373) );
  XNOR2_X1 U439 ( .A(n373), .B(KEYINPUT47), .ZN(n378) );
  NOR2_X1 U440 ( .A1(n558), .A2(n492), .ZN(n374) );
  XOR2_X1 U441 ( .A(KEYINPUT45), .B(n374), .Z(n375) );
  NOR2_X1 U442 ( .A1(n589), .A2(n375), .ZN(n376) );
  NAND2_X1 U443 ( .A1(n376), .A2(n585), .ZN(n377) );
  NAND2_X1 U444 ( .A1(n378), .A2(n377), .ZN(n380) );
  XNOR2_X1 U445 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n379) );
  XNOR2_X1 U446 ( .A(n380), .B(n379), .ZN(n547) );
  XOR2_X1 U447 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n382) );
  XNOR2_X1 U448 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n381) );
  XNOR2_X1 U449 ( .A(n382), .B(n381), .ZN(n452) );
  XNOR2_X1 U450 ( .A(n383), .B(n452), .ZN(n399) );
  XOR2_X1 U451 ( .A(KEYINPUT98), .B(KEYINPUT100), .Z(n385) );
  XNOR2_X1 U452 ( .A(G92GAT), .B(KEYINPUT99), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n385), .B(n384), .ZN(n391) );
  NAND2_X1 U454 ( .A1(G226GAT), .A2(G233GAT), .ZN(n387) );
  XOR2_X1 U455 ( .A(n391), .B(n390), .Z(n397) );
  XOR2_X1 U456 ( .A(KEYINPUT93), .B(G218GAT), .Z(n393) );
  XNOR2_X1 U457 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n392) );
  XNOR2_X1 U458 ( .A(n393), .B(n392), .ZN(n440) );
  XNOR2_X1 U459 ( .A(G197GAT), .B(n440), .ZN(n395) );
  XOR2_X1 U460 ( .A(n395), .B(n394), .Z(n396) );
  XNOR2_X1 U461 ( .A(n397), .B(n396), .ZN(n398) );
  INV_X1 U462 ( .A(n540), .ZN(n477) );
  NAND2_X1 U463 ( .A1(n547), .A2(n477), .ZN(n401) );
  XOR2_X1 U464 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n400) );
  XNOR2_X1 U465 ( .A(n401), .B(n400), .ZN(n423) );
  XOR2_X1 U466 ( .A(KEYINPUT6), .B(KEYINPUT95), .Z(n403) );
  XNOR2_X1 U467 ( .A(G1GAT), .B(G120GAT), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U469 ( .A(G155GAT), .B(G148GAT), .Z(n405) );
  XNOR2_X1 U470 ( .A(G29GAT), .B(G127GAT), .ZN(n404) );
  XNOR2_X1 U471 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n407), .B(n406), .ZN(n422) );
  XOR2_X1 U473 ( .A(KEYINPUT96), .B(KEYINPUT1), .Z(n409) );
  XNOR2_X1 U474 ( .A(KEYINPUT97), .B(KEYINPUT4), .ZN(n408) );
  XNOR2_X1 U475 ( .A(n409), .B(n408), .ZN(n414) );
  XOR2_X1 U476 ( .A(G85GAT), .B(n410), .Z(n412) );
  XOR2_X1 U477 ( .A(G113GAT), .B(KEYINPUT0), .Z(n450) );
  XNOR2_X1 U478 ( .A(n450), .B(G162GAT), .ZN(n411) );
  XNOR2_X1 U479 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U480 ( .A(n414), .B(n413), .Z(n416) );
  NAND2_X1 U481 ( .A1(G225GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U482 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U483 ( .A(n417), .B(G57GAT), .Z(n420) );
  XNOR2_X1 U484 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n418) );
  XNOR2_X1 U485 ( .A(n418), .B(KEYINPUT2), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n428), .B(KEYINPUT5), .ZN(n419) );
  XNOR2_X1 U487 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U488 ( .A(n422), .B(n421), .ZN(n538) );
  NAND2_X1 U489 ( .A1(n423), .A2(n538), .ZN(n424) );
  XNOR2_X1 U490 ( .A(n424), .B(KEYINPUT65), .ZN(n469) );
  XOR2_X1 U491 ( .A(KEYINPUT91), .B(KEYINPUT22), .Z(n426) );
  NAND2_X1 U492 ( .A1(G228GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U493 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U494 ( .A(n427), .B(KEYINPUT24), .Z(n431) );
  XNOR2_X1 U495 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U496 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U497 ( .A(G204GAT), .B(KEYINPUT23), .Z(n433) );
  XNOR2_X1 U498 ( .A(KEYINPUT92), .B(KEYINPUT94), .ZN(n432) );
  XNOR2_X1 U499 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U500 ( .A(n435), .B(n434), .Z(n439) );
  XNOR2_X1 U501 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U502 ( .A(n439), .B(n438), .ZN(n442) );
  XOR2_X1 U503 ( .A(G197GAT), .B(n440), .Z(n441) );
  XOR2_X1 U504 ( .A(n442), .B(n441), .Z(n485) );
  NAND2_X1 U505 ( .A1(n469), .A2(n485), .ZN(n443) );
  XNOR2_X1 U506 ( .A(n443), .B(KEYINPUT55), .ZN(n463) );
  XOR2_X1 U507 ( .A(KEYINPUT90), .B(G176GAT), .Z(n445) );
  XNOR2_X1 U508 ( .A(G43GAT), .B(G99GAT), .ZN(n444) );
  XNOR2_X1 U509 ( .A(n445), .B(n444), .ZN(n462) );
  XOR2_X1 U510 ( .A(G190GAT), .B(G134GAT), .Z(n449) );
  XNOR2_X1 U511 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U512 ( .A(n449), .B(n448), .ZN(n451) );
  XOR2_X1 U513 ( .A(n451), .B(n450), .Z(n460) );
  XNOR2_X1 U514 ( .A(n452), .B(G183GAT), .ZN(n454) );
  AND2_X1 U515 ( .A1(G227GAT), .A2(G233GAT), .ZN(n453) );
  XNOR2_X1 U516 ( .A(n454), .B(n453), .ZN(n458) );
  XOR2_X1 U517 ( .A(KEYINPUT87), .B(KEYINPUT20), .Z(n456) );
  XNOR2_X1 U518 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n455) );
  XNOR2_X1 U519 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U520 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U521 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U522 ( .A(n462), .B(n461), .ZN(n513) );
  NAND2_X1 U523 ( .A1(n463), .A2(n513), .ZN(n464) );
  NAND2_X1 U524 ( .A1(n581), .A2(n569), .ZN(n468) );
  XOR2_X1 U525 ( .A(G176GAT), .B(KEYINPUT56), .Z(n466) );
  XNOR2_X1 U526 ( .A(KEYINPUT124), .B(KEYINPUT57), .ZN(n465) );
  XNOR2_X1 U527 ( .A(n468), .B(n467), .ZN(G1349GAT) );
  INV_X1 U528 ( .A(n469), .ZN(n471) );
  NOR2_X1 U529 ( .A1(n513), .A2(n485), .ZN(n470) );
  XOR2_X1 U530 ( .A(n470), .B(KEYINPUT26), .Z(n566) );
  INV_X1 U531 ( .A(n593), .ZN(n584) );
  NOR2_X1 U532 ( .A1(n492), .A2(n584), .ZN(n475) );
  XNOR2_X1 U533 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n473) );
  NOR2_X1 U534 ( .A1(n589), .A2(n585), .ZN(n476) );
  XOR2_X1 U535 ( .A(KEYINPUT77), .B(n476), .Z(n507) );
  XNOR2_X1 U536 ( .A(n540), .B(KEYINPUT27), .ZN(n484) );
  OR2_X1 U537 ( .A1(n566), .A2(n484), .ZN(n481) );
  NAND2_X1 U538 ( .A1(n477), .A2(n513), .ZN(n478) );
  NAND2_X1 U539 ( .A1(n485), .A2(n478), .ZN(n479) );
  XOR2_X1 U540 ( .A(KEYINPUT25), .B(n479), .Z(n480) );
  NAND2_X1 U541 ( .A1(n481), .A2(n480), .ZN(n482) );
  NAND2_X1 U542 ( .A1(n482), .A2(n538), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n483), .B(KEYINPUT103), .ZN(n489) );
  NOR2_X1 U544 ( .A1(n538), .A2(n484), .ZN(n548) );
  XNOR2_X1 U545 ( .A(n485), .B(KEYINPUT28), .ZN(n551) );
  NOR2_X1 U546 ( .A1(n513), .A2(n486), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n487), .B(KEYINPUT102), .ZN(n488) );
  NOR2_X1 U548 ( .A1(n489), .A2(n488), .ZN(n506) );
  INV_X1 U549 ( .A(n558), .ZN(n592) );
  NOR2_X1 U550 ( .A1(n506), .A2(n592), .ZN(n490) );
  XOR2_X1 U551 ( .A(n490), .B(KEYINPUT106), .Z(n491) );
  NOR2_X1 U552 ( .A1(n492), .A2(n491), .ZN(n496) );
  INV_X1 U553 ( .A(KEYINPUT107), .ZN(n494) );
  NAND2_X1 U554 ( .A1(n507), .A2(n537), .ZN(n498) );
  XOR2_X1 U555 ( .A(KEYINPUT38), .B(KEYINPUT108), .Z(n497) );
  XNOR2_X1 U556 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U557 ( .A(KEYINPUT109), .B(n499), .ZN(n524) );
  NOR2_X1 U558 ( .A1(n538), .A2(n524), .ZN(n502) );
  XNOR2_X1 U559 ( .A(KEYINPUT110), .B(KEYINPUT39), .ZN(n500) );
  XNOR2_X1 U560 ( .A(KEYINPUT34), .B(KEYINPUT105), .ZN(n510) );
  NAND2_X1 U561 ( .A1(n592), .A2(n562), .ZN(n503) );
  XNOR2_X1 U562 ( .A(n503), .B(KEYINPUT16), .ZN(n504) );
  XNOR2_X1 U563 ( .A(n504), .B(KEYINPUT86), .ZN(n505) );
  NOR2_X1 U564 ( .A1(n506), .A2(n505), .ZN(n527) );
  NAND2_X1 U565 ( .A1(n527), .A2(n507), .ZN(n508) );
  XNOR2_X1 U566 ( .A(n508), .B(KEYINPUT104), .ZN(n516) );
  NOR2_X1 U567 ( .A1(n538), .A2(n516), .ZN(n509) );
  XNOR2_X1 U568 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U569 ( .A(G1GAT), .B(n511), .ZN(G1324GAT) );
  NOR2_X1 U570 ( .A1(n516), .A2(n540), .ZN(n512) );
  XOR2_X1 U571 ( .A(G8GAT), .B(n512), .Z(G1325GAT) );
  XNOR2_X1 U572 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n515) );
  INV_X1 U573 ( .A(n513), .ZN(n549) );
  NOR2_X1 U574 ( .A1(n549), .A2(n516), .ZN(n514) );
  XNOR2_X1 U575 ( .A(n515), .B(n514), .ZN(G1326GAT) );
  NOR2_X1 U576 ( .A1(n516), .A2(n551), .ZN(n517) );
  XOR2_X1 U577 ( .A(G22GAT), .B(n517), .Z(G1327GAT) );
  NOR2_X1 U578 ( .A1(n540), .A2(n524), .ZN(n519) );
  XNOR2_X1 U579 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n518) );
  XNOR2_X1 U580 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U581 ( .A(n520), .B(G36GAT), .ZN(G1329GAT) );
  NOR2_X1 U582 ( .A1(n524), .A2(n549), .ZN(n522) );
  XNOR2_X1 U583 ( .A(KEYINPUT40), .B(KEYINPUT113), .ZN(n521) );
  XNOR2_X1 U584 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U585 ( .A(n523), .B(G43GAT), .ZN(G1330GAT) );
  NOR2_X1 U586 ( .A1(n551), .A2(n524), .ZN(n525) );
  XOR2_X1 U587 ( .A(G50GAT), .B(n525), .Z(G1331GAT) );
  INV_X1 U588 ( .A(n585), .ZN(n576) );
  NOR2_X1 U589 ( .A1(n576), .A2(n526), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n536), .A2(n527), .ZN(n533) );
  NOR2_X1 U591 ( .A1(n538), .A2(n533), .ZN(n528) );
  XOR2_X1 U592 ( .A(G57GAT), .B(n528), .Z(n529) );
  XNOR2_X1 U593 ( .A(KEYINPUT42), .B(n529), .ZN(G1332GAT) );
  NOR2_X1 U594 ( .A1(n540), .A2(n533), .ZN(n530) );
  XOR2_X1 U595 ( .A(KEYINPUT114), .B(n530), .Z(n531) );
  XNOR2_X1 U596 ( .A(G64GAT), .B(n531), .ZN(G1333GAT) );
  NOR2_X1 U597 ( .A1(n549), .A2(n533), .ZN(n532) );
  XOR2_X1 U598 ( .A(G71GAT), .B(n532), .Z(G1334GAT) );
  NOR2_X1 U599 ( .A1(n551), .A2(n533), .ZN(n535) );
  XNOR2_X1 U600 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(G1335GAT) );
  NAND2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n544) );
  NOR2_X1 U603 ( .A1(n538), .A2(n544), .ZN(n539) );
  XOR2_X1 U604 ( .A(G85GAT), .B(n539), .Z(G1336GAT) );
  NOR2_X1 U605 ( .A1(n540), .A2(n544), .ZN(n542) );
  XNOR2_X1 U606 ( .A(G92GAT), .B(KEYINPUT115), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(G1337GAT) );
  NOR2_X1 U608 ( .A1(n549), .A2(n544), .ZN(n543) );
  XOR2_X1 U609 ( .A(G99GAT), .B(n543), .Z(G1338GAT) );
  NOR2_X1 U610 ( .A1(n551), .A2(n544), .ZN(n545) );
  XOR2_X1 U611 ( .A(KEYINPUT44), .B(n545), .Z(n546) );
  XNOR2_X1 U612 ( .A(G106GAT), .B(n546), .ZN(G1339GAT) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n565) );
  NOR2_X1 U614 ( .A1(n549), .A2(n565), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n550), .B(KEYINPUT118), .ZN(n552) );
  NAND2_X1 U616 ( .A1(n552), .A2(n551), .ZN(n561) );
  NOR2_X1 U617 ( .A1(n585), .A2(n561), .ZN(n553) );
  XOR2_X1 U618 ( .A(G113GAT), .B(n553), .Z(G1340GAT) );
  NOR2_X1 U619 ( .A1(n561), .A2(n526), .ZN(n557) );
  XOR2_X1 U620 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n555) );
  XNOR2_X1 U621 ( .A(G120GAT), .B(KEYINPUT120), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1341GAT) );
  NOR2_X1 U624 ( .A1(n558), .A2(n561), .ZN(n559) );
  XOR2_X1 U625 ( .A(KEYINPUT50), .B(n559), .Z(n560) );
  XNOR2_X1 U626 ( .A(G127GAT), .B(n560), .ZN(G1342GAT) );
  NOR2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n564) );
  XNOR2_X1 U628 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(G1343GAT) );
  XOR2_X1 U630 ( .A(G141GAT), .B(KEYINPUT121), .Z(n568) );
  NOR2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n574) );
  NAND2_X1 U632 ( .A1(n574), .A2(n576), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G1344GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n571) );
  NAND2_X1 U635 ( .A1(n574), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G148GAT), .B(n572), .ZN(G1345GAT) );
  NAND2_X1 U638 ( .A1(n574), .A2(n592), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U640 ( .A1(n580), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U642 ( .A1(n576), .A2(n581), .ZN(n577) );
  XNOR2_X1 U643 ( .A(G169GAT), .B(n577), .ZN(G1348GAT) );
  XOR2_X1 U644 ( .A(G183GAT), .B(KEYINPUT125), .Z(n579) );
  NAND2_X1 U645 ( .A1(n581), .A2(n592), .ZN(n578) );
  XNOR2_X1 U646 ( .A(n579), .B(n578), .ZN(G1350GAT) );
  XNOR2_X1 U647 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n583) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(G1351GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n587) );
  XNOR2_X1 U651 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(G197GAT), .B(n588), .ZN(G1352GAT) );
  XOR2_X1 U654 ( .A(G204GAT), .B(KEYINPUT61), .Z(n591) );
  NAND2_X1 U655 ( .A1(n593), .A2(n589), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n591), .B(n590), .ZN(G1353GAT) );
  NAND2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(n594), .B(G211GAT), .ZN(G1354GAT) );
endmodule

