//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n635, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926;
  NOR2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT77), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G141gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT76), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G141gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G148gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n208), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n211), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n204), .A2(KEYINPUT2), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n203), .A2(KEYINPUT77), .A3(new_n204), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n207), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(KEYINPUT74), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT74), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n220), .A3(KEYINPUT2), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n213), .A2(new_n209), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT73), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n204), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(KEYINPUT73), .A2(G155gat), .A3(G162gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n202), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n223), .A2(KEYINPUT75), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT75), .B1(new_n223), .B2(new_n227), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n218), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT3), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n232), .B(new_n218), .C1(new_n228), .C2(new_n229), .ZN(new_n233));
  XOR2_X1   g032(.A(G127gat), .B(G134gat), .Z(new_n234));
  NOR2_X1   g033(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n235));
  INV_X1    g034(.A(G120gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT68), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G120gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n239), .A3(G113gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n236), .A2(G113gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT69), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n243), .B1(new_n236), .B2(G113gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT1), .ZN(new_n246));
  INV_X1    g045(.A(G113gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n247), .A2(G120gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n246), .B1(new_n241), .B2(new_n248), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n235), .A2(new_n245), .B1(new_n249), .B2(new_n234), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n231), .A2(new_n233), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G225gat), .A2(G233gat), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n218), .B(new_n250), .C1(new_n228), .C2(new_n229), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n229), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n223), .A2(KEYINPUT75), .A3(new_n227), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n259), .A2(KEYINPUT4), .A3(new_n218), .A4(new_n250), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n252), .A2(new_n253), .A3(new_n256), .A4(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT5), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n230), .A2(new_n251), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n254), .ZN(new_n264));
  INV_X1    g063(.A(new_n253), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n262), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n260), .A2(new_n256), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n268), .A2(new_n262), .A3(new_n253), .A4(new_n252), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G1gat), .B(G29gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT0), .ZN(new_n272));
  XNOR2_X1  g071(.A(G57gat), .B(G85gat), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n272), .B(new_n273), .Z(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n267), .A2(new_n274), .A3(new_n269), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n270), .A2(KEYINPUT6), .A3(new_n275), .ZN(new_n280));
  NAND2_X1  g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281));
  INV_X1    g080(.A(G169gat), .ZN(new_n282));
  INV_X1    g081(.A(G176gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT26), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n281), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT26), .B1(new_n282), .B2(new_n283), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT27), .B(G183gat), .ZN(new_n290));
  INV_X1    g089(.A(G190gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n292), .A2(new_n293), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n289), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT23), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT23), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(G169gat), .B2(G176gat), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n297), .A2(new_n299), .A3(new_n287), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(new_n281), .ZN(new_n302));
  NAND3_X1  g101(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n300), .A2(KEYINPUT25), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT65), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n306), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n303), .A2(KEYINPUT65), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n302), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT25), .B1(new_n300), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT66), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n305), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AOI211_X1 g111(.A(KEYINPUT66), .B(KEYINPUT25), .C1(new_n300), .C2(new_n309), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n296), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n315));
  INV_X1    g114(.A(G226gat), .ZN(new_n316));
  INV_X1    g115(.A(G233gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n314), .A2(new_n315), .A3(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G197gat), .B(G204gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT22), .ZN(new_n322));
  INV_X1    g121(.A(G211gat), .ZN(new_n323));
  INV_X1    g122(.A(G218gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G211gat), .B(G218gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n321), .A3(new_n325), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n329), .A2(KEYINPUT72), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT72), .B1(new_n329), .B2(new_n330), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n318), .B(new_n296), .C1(new_n312), .C2(new_n313), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n334), .B1(new_n320), .B2(new_n335), .ZN(new_n338));
  XNOR2_X1  g137(.A(G8gat), .B(G36gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(G64gat), .B(G92gat), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n339), .B(new_n340), .Z(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  OR4_X1    g141(.A1(KEYINPUT30), .A2(new_n337), .A3(new_n338), .A4(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n342), .B1(new_n337), .B2(new_n338), .ZN(new_n344));
  INV_X1    g143(.A(new_n338), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n345), .A2(new_n336), .A3(new_n341), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n346), .A3(KEYINPUT30), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n279), .A2(new_n280), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT87), .B(KEYINPUT35), .ZN(new_n349));
  XOR2_X1   g148(.A(G78gat), .B(G106gat), .Z(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(KEYINPUT79), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n351), .B(G50gat), .Z(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT78), .B(KEYINPUT31), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT29), .B1(new_n329), .B2(new_n330), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n230), .B1(KEYINPUT3), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT82), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n233), .A2(new_n315), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n334), .ZN(new_n361));
  NAND2_X1  g160(.A1(G228gat), .A2(G233gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n230), .B(KEYINPUT82), .C1(KEYINPUT3), .C2(new_n356), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n359), .A2(new_n361), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n362), .B(KEYINPUT80), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n329), .A2(KEYINPUT81), .A3(new_n330), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n367), .B(new_n315), .C1(KEYINPUT81), .C2(new_n329), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n368), .A2(new_n232), .B1(new_n259), .B2(new_n218), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n333), .B1(new_n233), .B2(new_n315), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n366), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G22gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n365), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n372), .B1(new_n365), .B2(new_n371), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n355), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n365), .A2(new_n371), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G22gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n378), .A2(new_n373), .A3(new_n354), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n349), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n314), .A2(new_n250), .ZN(new_n381));
  NAND2_X1  g180(.A1(G227gat), .A2(G233gat), .ZN(new_n382));
  XOR2_X1   g181(.A(new_n382), .B(KEYINPUT64), .Z(new_n383));
  OAI211_X1 g182(.A(new_n251), .B(new_n296), .C1(new_n312), .C2(new_n313), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n381), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT32), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT33), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  XOR2_X1   g187(.A(G15gat), .B(G43gat), .Z(new_n389));
  XNOR2_X1  g188(.A(G71gat), .B(G99gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n386), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n391), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n385), .B(KEYINPUT32), .C1(new_n387), .C2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n381), .A2(new_n384), .ZN(new_n397));
  OAI211_X1 g196(.A(KEYINPUT70), .B(new_n396), .C1(new_n397), .C2(new_n383), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n383), .B1(new_n381), .B2(new_n384), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT70), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n395), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AND4_X1   g200(.A1(new_n392), .A2(new_n394), .A3(new_n398), .A4(new_n401), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n392), .A2(new_n394), .B1(new_n398), .B2(new_n401), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT86), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n392), .A2(new_n394), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n398), .A2(new_n401), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n392), .A2(new_n394), .A3(new_n398), .A4(new_n401), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT86), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n348), .B(new_n380), .C1(new_n405), .C2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT88), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n279), .A2(new_n280), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n402), .A2(new_n403), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n376), .A2(new_n379), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n343), .A2(new_n347), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n411), .A2(new_n412), .B1(KEYINPUT35), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n404), .B1(new_n402), .B2(new_n403), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n408), .A2(KEYINPUT86), .A3(new_n409), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n421), .A2(KEYINPUT88), .A3(new_n348), .A4(new_n380), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n343), .A2(new_n347), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n268), .A2(new_n252), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n265), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n274), .B1(new_n425), .B2(KEYINPUT39), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT40), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n427), .A2(KEYINPUT83), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT39), .B1(new_n264), .B2(new_n265), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n429), .B1(new_n424), .B2(new_n265), .ZN(new_n430));
  OR3_X1    g229(.A1(new_n426), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  OAI211_X1 g230(.A(KEYINPUT83), .B(new_n427), .C1(new_n426), .C2(new_n430), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n423), .A2(new_n431), .A3(new_n276), .A4(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n342), .A2(KEYINPUT37), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT38), .B1(new_n344), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT37), .B1(new_n337), .B2(new_n338), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT84), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT84), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n438), .B(KEYINPUT37), .C1(new_n337), .C2(new_n338), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n435), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT85), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n435), .A2(new_n442), .A3(new_n437), .A4(new_n439), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n341), .B1(new_n345), .B2(new_n336), .ZN(new_n445));
  INV_X1    g244(.A(new_n434), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n436), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT38), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n448), .A2(new_n279), .A3(new_n280), .A4(new_n346), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n415), .B(new_n433), .C1(new_n444), .C2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n415), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n413), .A2(new_n416), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n414), .A2(KEYINPUT36), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT36), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n454), .B1(new_n402), .B2(new_n403), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n451), .A2(new_n452), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n418), .A2(new_n422), .B1(new_n450), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G43gat), .B(G50gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT15), .ZN(new_n459));
  NAND2_X1  g258(.A1(G29gat), .A2(G36gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NOR3_X1   g262(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n464));
  OAI22_X1  g263(.A1(new_n458), .A2(KEYINPUT15), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT89), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n464), .B1(new_n468), .B2(new_n462), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n469), .B1(new_n468), .B2(new_n462), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n470), .A2(new_n460), .ZN(new_n471));
  OAI211_X1 g270(.A(KEYINPUT90), .B(new_n467), .C1(new_n471), .C2(new_n459), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT90), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n459), .B1(new_n470), .B2(new_n460), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n473), .B1(new_n474), .B2(new_n466), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G15gat), .B(G22gat), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT91), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n480), .A2(G1gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(new_n479), .A3(G1gat), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT16), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(G8gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n477), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(G8gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n485), .B(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n476), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(G229gat), .A2(G233gat), .ZN(new_n492));
  XOR2_X1   g291(.A(new_n492), .B(KEYINPUT13), .Z(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT92), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT17), .B1(new_n472), .B2(new_n475), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n467), .B1(new_n471), .B2(new_n459), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n498), .A2(KEYINPUT17), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n489), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n500), .A2(new_n487), .A3(KEYINPUT18), .A4(new_n492), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n491), .A2(KEYINPUT92), .A3(new_n493), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n496), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n500), .A2(new_n492), .A3(new_n487), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT18), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G113gat), .B(G141gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(G197gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT11), .B(G169gat), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n509), .B(new_n510), .Z(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT12), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n506), .B(KEYINPUT93), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n496), .A2(new_n501), .A3(new_n502), .A4(new_n512), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n507), .A2(new_n513), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n457), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G71gat), .A2(G78gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT9), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT97), .ZN(new_n522));
  XNOR2_X1  g321(.A(G57gat), .B(G64gat), .ZN(new_n523));
  OR2_X1    g322(.A1(G71gat), .A2(G78gat), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n523), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT98), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT98), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n522), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(G57gat), .B(G64gat), .Z(new_n531));
  INV_X1    g330(.A(KEYINPUT95), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n523), .A2(KEYINPUT95), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(new_n521), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n524), .B1(KEYINPUT94), .B2(new_n519), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n536), .B1(KEYINPUT94), .B2(new_n519), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n535), .A2(KEYINPUT96), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT96), .B1(new_n535), .B2(new_n537), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n530), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT21), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G127gat), .B(G155gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n489), .B1(new_n541), .B2(new_n542), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G231gat), .A2(G233gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT99), .ZN(new_n549));
  XOR2_X1   g348(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G183gat), .B(G211gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n547), .A2(new_n553), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT100), .B(KEYINPUT7), .ZN(new_n558));
  INV_X1    g357(.A(G85gat), .ZN(new_n559));
  INV_X1    g358(.A(G92gat), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n558), .B(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT101), .B1(G99gat), .B2(G106gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT8), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(KEYINPUT101), .A2(G99gat), .A3(G106gat), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n565), .A2(new_n566), .B1(new_n559), .B2(new_n560), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G99gat), .B(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n562), .A2(new_n569), .A3(new_n567), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(KEYINPUT102), .A3(new_n572), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n572), .A2(KEYINPUT102), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AND2_X1   g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n477), .A2(new_n575), .B1(KEYINPUT41), .B2(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n574), .B(new_n573), .C1(new_n497), .C2(new_n499), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G190gat), .B(G218gat), .Z(new_n580));
  AND2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n579), .A2(new_n580), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n576), .A2(KEYINPUT41), .ZN(new_n583));
  XNOR2_X1  g382(.A(G134gat), .B(G162gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  OR3_X1    g385(.A1(new_n581), .A2(new_n582), .A3(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n586), .B1(new_n581), .B2(new_n582), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n557), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G230gat), .A2(G233gat), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT103), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n535), .A2(new_n537), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT96), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n596), .A2(new_n538), .B1(new_n527), .B2(new_n529), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n593), .B1(new_n575), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(new_n572), .A3(new_n571), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n541), .A2(KEYINPUT103), .A3(new_n574), .A4(new_n573), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n592), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n592), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT104), .B(KEYINPUT10), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n598), .A2(new_n601), .A3(new_n599), .A4(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n575), .A2(KEYINPUT10), .A3(new_n597), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G120gat), .B(G148gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(G176gat), .B(G204gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  OR3_X1    g410(.A1(new_n602), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n611), .B1(new_n602), .B2(new_n607), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n591), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n518), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n618), .A2(new_n413), .ZN(new_n619));
  XOR2_X1   g418(.A(KEYINPUT105), .B(G1gat), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(G1324gat));
  INV_X1    g420(.A(new_n618), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n488), .B1(new_n622), .B2(new_n423), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT16), .B(G8gat), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n618), .A2(new_n416), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(KEYINPUT42), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(KEYINPUT42), .B2(new_n625), .ZN(G1325gat));
  NAND2_X1  g426(.A1(new_n453), .A2(new_n455), .ZN(new_n628));
  OAI21_X1  g427(.A(G15gat), .B1(new_n618), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n405), .A2(new_n410), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n630), .A2(G15gat), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n629), .B1(new_n618), .B2(new_n631), .ZN(G1326gat));
  NAND2_X1  g431(.A1(new_n518), .A2(new_n451), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n633), .A2(new_n616), .ZN(new_n634));
  XOR2_X1   g433(.A(KEYINPUT43), .B(G22gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(G1327gat));
  NAND3_X1  g435(.A1(new_n413), .A2(new_n380), .A3(new_n416), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n412), .B1(new_n630), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n417), .A2(KEYINPUT35), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(new_n422), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n450), .A2(new_n456), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n556), .A2(new_n614), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(new_n517), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n642), .A2(new_n590), .A3(new_n645), .ZN(new_n646));
  NOR3_X1   g445(.A1(new_n646), .A2(G29gat), .A3(new_n413), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n647), .B(KEYINPUT45), .Z(new_n648));
  INV_X1    g447(.A(KEYINPUT106), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n650), .B1(new_n457), .B2(new_n589), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n642), .A2(KEYINPUT44), .A3(new_n590), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n645), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n649), .B1(new_n654), .B2(new_n413), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(G29gat), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n654), .A2(new_n649), .A3(new_n413), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n648), .B1(new_n656), .B2(new_n657), .ZN(G1328gat));
  OAI21_X1  g457(.A(G36gat), .B1(new_n654), .B2(new_n416), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n646), .A2(G36gat), .A3(new_n416), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT46), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(G1329gat));
  INV_X1    g461(.A(new_n628), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(G43gat), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n646), .A2(new_n630), .ZN(new_n665));
  OAI22_X1  g464(.A1(new_n654), .A2(new_n664), .B1(G43gat), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g466(.A(G50gat), .B1(new_n654), .B2(new_n415), .ZN(new_n668));
  OR3_X1    g467(.A1(new_n644), .A2(G50gat), .A3(new_n589), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n668), .B1(new_n633), .B2(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1331gat));
  AND4_X1   g471(.A1(new_n517), .A2(new_n642), .A3(new_n591), .A4(new_n614), .ZN(new_n673));
  INV_X1    g472(.A(new_n413), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G57gat), .ZN(G1332gat));
  INV_X1    g475(.A(KEYINPUT49), .ZN(new_n677));
  INV_X1    g476(.A(G64gat), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n423), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT108), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n673), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n677), .A2(new_n678), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1333gat));
  XNOR2_X1  g482(.A(new_n421), .B(KEYINPUT109), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(G71gat), .B1(new_n673), .B2(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n663), .A2(G71gat), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n686), .B1(new_n673), .B2(new_n687), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n451), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G78gat), .ZN(G1335gat));
  OAI21_X1  g490(.A(new_n513), .B1(new_n503), .B2(new_n506), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n504), .A2(new_n505), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT93), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n694), .B2(new_n515), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n695), .A2(new_n615), .A3(new_n556), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n651), .A2(new_n652), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT110), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT110), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n651), .A2(new_n699), .A3(new_n652), .A4(new_n696), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n698), .A2(new_n674), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n559), .B1(new_n701), .B2(KEYINPUT111), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(KEYINPUT111), .B2(new_n701), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n695), .A2(new_n556), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n642), .A2(new_n590), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT51), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n642), .A2(KEYINPUT51), .A3(new_n590), .A4(new_n704), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n614), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n711), .A2(new_n559), .A3(new_n674), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n703), .A2(new_n712), .ZN(G1336gat));
  OAI21_X1  g512(.A(G92gat), .B1(new_n697), .B2(new_n416), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT52), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n416), .A2(G92gat), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n714), .B(new_n715), .C1(new_n710), .C2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT114), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n698), .A2(new_n423), .A3(new_n700), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n707), .A2(KEYINPUT112), .A3(new_n708), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT112), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n705), .A2(new_n722), .A3(new_n706), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n615), .A2(new_n717), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n721), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n720), .A2(G92gat), .B1(new_n725), .B2(KEYINPUT113), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT113), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n721), .A2(new_n727), .A3(new_n723), .A4(new_n724), .ZN(new_n728));
  AOI211_X1 g527(.A(new_n719), .B(new_n715), .C1(new_n726), .C2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n720), .A2(G92gat), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n725), .A2(KEYINPUT113), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT114), .B1(new_n732), .B2(KEYINPUT52), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n718), .B1(new_n729), .B2(new_n733), .ZN(G1337gat));
  NAND3_X1  g533(.A1(new_n698), .A2(new_n663), .A3(new_n700), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G99gat), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n630), .A2(G99gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n710), .B2(new_n737), .ZN(G1338gat));
  NOR2_X1   g537(.A1(new_n415), .A2(G106gat), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT53), .B1(new_n711), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT115), .ZN(new_n741));
  OAI21_X1  g540(.A(G106gat), .B1(new_n697), .B2(new_n415), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n741), .B1(new_n740), .B2(new_n742), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT53), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n698), .A2(new_n451), .A3(new_n700), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n721), .A2(new_n723), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n614), .A2(new_n739), .ZN(new_n748));
  AOI22_X1  g547(.A1(G106gat), .A2(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI22_X1  g548(.A1(new_n743), .A2(new_n744), .B1(new_n745), .B2(new_n749), .ZN(G1339gat));
  NAND2_X1  g549(.A1(new_n605), .A2(new_n606), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n592), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT54), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n606), .A2(new_n603), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n753), .B1(new_n605), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n610), .B1(new_n607), .B2(new_n753), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n758), .A2(KEYINPUT55), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT117), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n756), .A2(new_n757), .A3(KEYINPUT116), .A4(KEYINPUT55), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n612), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT55), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n752), .B2(new_n755), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT116), .B1(new_n764), .B2(new_n757), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n760), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n757), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT116), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n769), .A2(KEYINPUT117), .A3(new_n612), .A4(new_n761), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n759), .B1(new_n766), .B2(new_n770), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n500), .A2(new_n487), .ZN(new_n772));
  OAI22_X1  g571(.A1(new_n772), .A2(new_n492), .B1(new_n491), .B2(new_n493), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n511), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n694), .B2(new_n515), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n771), .A2(new_n590), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(KEYINPUT118), .A3(new_n614), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n615), .B2(new_n775), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n771), .B2(new_n695), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n777), .B1(new_n782), .B2(new_n590), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n557), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n616), .A2(new_n695), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n413), .A2(new_n423), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n787), .A2(new_n415), .A3(new_n421), .A4(new_n788), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n789), .A2(new_n247), .A3(new_n517), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n785), .B1(new_n783), .B2(new_n557), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n414), .A2(new_n415), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n791), .A2(new_n413), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n416), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n695), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n790), .B1(new_n796), .B2(new_n247), .ZN(G1340gat));
  OAI21_X1  g596(.A(G120gat), .B1(new_n789), .B2(new_n615), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n614), .A2(new_n237), .A3(new_n239), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n794), .B2(new_n799), .ZN(G1341gat));
  OAI21_X1  g599(.A(G127gat), .B1(new_n789), .B2(new_n557), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n557), .A2(G127gat), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n794), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n801), .B(KEYINPUT119), .C1(new_n794), .C2(new_n802), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(G1342gat));
  INV_X1    g606(.A(new_n793), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n589), .A2(new_n423), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n810), .A2(G134gat), .ZN(new_n811));
  OR3_X1    g610(.A1(new_n808), .A2(KEYINPUT56), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(G134gat), .B1(new_n789), .B2(new_n589), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT56), .B1(new_n808), .B2(new_n811), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(G1343gat));
  NAND2_X1  g614(.A1(new_n628), .A2(new_n788), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n695), .B1(KEYINPUT55), .B2(new_n758), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n769), .A2(new_n612), .A3(new_n761), .ZN(new_n818));
  OAI22_X1  g617(.A1(new_n817), .A2(new_n818), .B1(new_n615), .B2(new_n775), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n589), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n556), .B1(new_n777), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n451), .B1(new_n821), .B2(new_n785), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n816), .B1(new_n822), .B2(KEYINPUT57), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824));
  AOI211_X1 g623(.A(new_n517), .B(new_n759), .C1(new_n766), .C2(new_n770), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n589), .B1(new_n825), .B2(new_n781), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n556), .B1(new_n826), .B2(new_n777), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n824), .B(new_n451), .C1(new_n827), .C2(new_n785), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n823), .A2(new_n828), .A3(new_n695), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(G141gat), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n413), .B1(new_n784), .B2(new_n786), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n663), .A2(new_n415), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n517), .A2(G141gat), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n831), .A2(new_n416), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n832), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n791), .A2(new_n413), .A3(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n838), .A2(KEYINPUT120), .A3(new_n416), .A4(new_n833), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n830), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT58), .ZN(new_n841));
  NOR2_X1   g640(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n842));
  AND2_X1   g641(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n830), .B(new_n834), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(new_n844), .ZN(G1344gat));
  INV_X1    g644(.A(new_n838), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n423), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n208), .A3(new_n614), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n823), .A2(new_n828), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(new_n615), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n850), .A2(KEYINPUT59), .A3(new_n208), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT57), .B1(new_n791), .B2(new_n415), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n785), .B(KEYINPUT122), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n824), .B(new_n451), .C1(new_n854), .C2(new_n821), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n816), .A2(new_n615), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n852), .B1(new_n857), .B2(G148gat), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n848), .B1(new_n851), .B2(new_n858), .ZN(G1345gat));
  INV_X1    g658(.A(G155gat), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n847), .A2(new_n860), .A3(new_n556), .ZN(new_n861));
  OAI21_X1  g660(.A(G155gat), .B1(new_n849), .B2(new_n557), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1346gat));
  NAND3_X1  g662(.A1(new_n823), .A2(new_n828), .A3(new_n590), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(G162gat), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n810), .A2(G162gat), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n865), .B1(new_n846), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT123), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT123), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n865), .B(new_n869), .C1(new_n846), .C2(new_n866), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(G1347gat));
  NOR2_X1   g670(.A1(new_n674), .A2(new_n416), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n684), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n787), .A2(new_n415), .A3(new_n874), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(new_n282), .A3(new_n517), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n791), .A2(new_n792), .A3(new_n873), .ZN(new_n877));
  AOI21_X1  g676(.A(G169gat), .B1(new_n877), .B2(new_n695), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n876), .A2(new_n878), .ZN(G1348gat));
  OAI21_X1  g678(.A(G176gat), .B1(new_n875), .B2(new_n615), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n877), .A2(new_n283), .A3(new_n614), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1349gat));
  OAI21_X1  g681(.A(G183gat), .B1(new_n875), .B2(new_n557), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n877), .A2(new_n290), .A3(new_n556), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g685(.A1(new_n877), .A2(new_n291), .A3(new_n590), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n875), .A2(new_n589), .ZN(new_n888));
  NOR2_X1   g687(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n291), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n889), .B1(new_n888), .B2(new_n890), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n887), .B1(new_n891), .B2(new_n892), .ZN(G1351gat));
  NOR2_X1   g692(.A1(new_n873), .A2(new_n663), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n853), .A2(new_n695), .A3(new_n855), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(G197gat), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n787), .A2(KEYINPUT125), .A3(new_n832), .A4(new_n872), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT125), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n832), .A2(new_n872), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n791), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n517), .A2(G197gat), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n897), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n896), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT126), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT126), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n896), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1352gat));
  AND2_X1   g706(.A1(new_n853), .A2(new_n855), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n614), .A3(new_n894), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(G204gat), .ZN(new_n910));
  NOR4_X1   g709(.A1(new_n791), .A2(G204gat), .A3(new_n615), .A4(new_n899), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n910), .A2(new_n913), .A3(new_n914), .ZN(G1353gat));
  INV_X1    g714(.A(KEYINPUT127), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n853), .A2(new_n556), .A3(new_n855), .A4(new_n894), .ZN(new_n917));
  AND4_X1   g716(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT63), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n323), .B1(KEYINPUT127), .B2(new_n919), .ZN(new_n920));
  AOI22_X1  g719(.A1(new_n917), .A2(new_n920), .B1(new_n916), .B2(KEYINPUT63), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n897), .A2(new_n900), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n556), .A2(new_n323), .ZN(new_n923));
  OAI22_X1  g722(.A1(new_n918), .A2(new_n921), .B1(new_n922), .B2(new_n923), .ZN(G1354gat));
  AND3_X1   g723(.A1(new_n908), .A2(new_n590), .A3(new_n894), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n590), .A2(new_n324), .ZN(new_n926));
  OAI22_X1  g725(.A1(new_n925), .A2(new_n324), .B1(new_n922), .B2(new_n926), .ZN(G1355gat));
endmodule


