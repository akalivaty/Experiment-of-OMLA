//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980, new_n981;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  NAND2_X1  g005(.A1(G229gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT16), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(new_n210), .B2(G1gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G1gat), .B2(new_n209), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(G8gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT90), .B(G36gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G29gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n217), .A2(KEYINPUT14), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(KEYINPUT14), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT15), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n216), .A2(KEYINPUT15), .A3(new_n218), .A4(new_n219), .ZN(new_n223));
  XNOR2_X1  g022(.A(G43gat), .B(G50gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT17), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n223), .A2(new_n224), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n226), .B1(new_n225), .B2(new_n227), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n214), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n225), .A2(new_n227), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT91), .B1(new_n232), .B2(new_n213), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  OAI211_X1 g033(.A(KEYINPUT91), .B(new_n214), .C1(new_n229), .C2(new_n230), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n208), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT18), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n232), .B(new_n213), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n240), .B(new_n208), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n242), .B1(new_n236), .B2(KEYINPUT18), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n206), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n236), .A2(KEYINPUT18), .ZN(new_n245));
  INV_X1    g044(.A(new_n206), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n245), .A2(new_n246), .A3(new_n237), .A4(new_n242), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT93), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT93), .B1(new_n244), .B2(new_n247), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G8gat), .B(G36gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(G64gat), .B(G92gat), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n253), .B(new_n254), .Z(new_n255));
  NAND2_X1  g054(.A1(G226gat), .A2(G233gat), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n256), .B(KEYINPUT72), .Z(new_n257));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT24), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n259), .A2(G183gat), .A3(G190gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(G183gat), .B(G190gat), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n260), .B1(new_n261), .B2(new_n259), .ZN(new_n262));
  INV_X1    g061(.A(G169gat), .ZN(new_n263));
  INV_X1    g062(.A(G176gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n264), .A3(KEYINPUT23), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT23), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n266), .B1(G169gat), .B2(G176gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(G169gat), .A2(G176gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n258), .B1(new_n262), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT65), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n265), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G190gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(G183gat), .ZN(new_n276));
  INV_X1    g075(.A(G183gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n277), .A2(G190gat), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT24), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n258), .B1(new_n280), .B2(new_n266), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n274), .A2(new_n279), .A3(new_n260), .A4(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n270), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n268), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n284), .B1(new_n280), .B2(KEYINPUT26), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT26), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n286), .A2(new_n263), .A3(new_n264), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n285), .A2(new_n287), .B1(G183gat), .B2(G190gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n277), .A2(KEYINPUT27), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT27), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G183gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(new_n291), .A3(new_n275), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT66), .ZN(new_n293));
  XNOR2_X1  g092(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n294), .B1(new_n292), .B2(new_n293), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n288), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n283), .A2(KEYINPUT74), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT74), .B1(new_n283), .B2(new_n297), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n257), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT29), .B1(new_n283), .B2(new_n297), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT73), .B1(new_n301), .B2(new_n257), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n303));
  INV_X1    g102(.A(new_n257), .ZN(new_n304));
  INV_X1    g103(.A(new_n296), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n307), .A2(new_n288), .B1(new_n270), .B2(new_n282), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n303), .B(new_n304), .C1(new_n308), .C2(KEYINPUT29), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n300), .A2(new_n302), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G211gat), .A2(G218gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT22), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(G197gat), .A2(G204gat), .ZN(new_n316));
  AND2_X1   g115(.A1(G197gat), .A2(G204gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n311), .B(new_n315), .C1(new_n316), .C2(new_n317), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n310), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n257), .A2(KEYINPUT29), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n324), .B1(new_n298), .B2(new_n299), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n283), .A2(new_n297), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(new_n304), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n321), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n255), .B1(new_n323), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT30), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n323), .A2(new_n330), .A3(new_n255), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n323), .A2(new_n330), .ZN(new_n337));
  INV_X1    g136(.A(new_n255), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n337), .A2(KEYINPUT30), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G1gat), .B(G29gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT0), .ZN(new_n343));
  XNOR2_X1  g142(.A(G57gat), .B(G85gat), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n343), .B(new_n344), .Z(new_n345));
  NAND2_X1  g144(.A1(G225gat), .A2(G233gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n346), .B(KEYINPUT79), .Z(new_n347));
  INV_X1    g146(.A(KEYINPUT78), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n349));
  AND2_X1   g148(.A1(G155gat), .A2(G162gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G155gat), .ZN(new_n353));
  INV_X1    g152(.A(G162gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(KEYINPUT75), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G141gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(G148gat), .ZN(new_n360));
  INV_X1    g159(.A(G148gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(G141gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT76), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n360), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT2), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(G155gat), .B2(G162gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n360), .A2(new_n362), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n366), .B1(new_n367), .B2(KEYINPUT76), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n358), .B1(new_n364), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n362), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n361), .A2(KEYINPUT77), .A3(G141gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(new_n360), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n356), .B1(new_n355), .B2(KEYINPUT2), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n348), .B1(new_n369), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n367), .A2(KEYINPUT76), .ZN(new_n378));
  INV_X1    g177(.A(new_n366), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(new_n364), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n358), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(KEYINPUT78), .A3(new_n375), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n377), .A2(new_n383), .A3(KEYINPUT3), .ZN(new_n384));
  XOR2_X1   g183(.A(G113gat), .B(G120gat), .Z(new_n385));
  INV_X1    g184(.A(KEYINPUT69), .ZN(new_n386));
  OR2_X1    g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G127gat), .B(G134gat), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT1), .ZN(new_n389));
  INV_X1    g188(.A(G120gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n390), .A3(G113gat), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT68), .ZN(new_n393));
  INV_X1    g192(.A(G127gat), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n393), .A2(new_n394), .A3(G134gat), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n395), .B1(new_n393), .B2(new_n388), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n385), .A2(new_n389), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n387), .A2(new_n392), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n380), .A2(new_n381), .B1(new_n373), .B2(new_n374), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n347), .B1(new_n384), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n399), .A2(new_n398), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT4), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT80), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n405), .B1(new_n369), .B2(new_n376), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n360), .A2(new_n362), .A3(new_n363), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n363), .B1(new_n360), .B2(new_n362), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n407), .A2(new_n408), .A3(new_n366), .ZN(new_n409));
  OAI211_X1 g208(.A(KEYINPUT80), .B(new_n375), .C1(new_n409), .C2(new_n358), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n406), .A2(new_n398), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n404), .B1(new_n411), .B2(KEYINPUT4), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT5), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n402), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n411), .A2(KEYINPUT4), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n398), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT81), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT81), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n399), .A2(new_n398), .A3(new_n419), .A4(new_n416), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n402), .B1(new_n415), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT82), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT5), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n387), .A2(new_n392), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n396), .A2(new_n397), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n377), .A2(new_n383), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n403), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT83), .B1(new_n429), .B2(new_n347), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT83), .ZN(new_n431));
  INV_X1    g230(.A(new_n347), .ZN(new_n432));
  AOI211_X1 g231(.A(new_n431), .B(new_n432), .C1(new_n428), .C2(new_n403), .ZN(new_n433));
  OAI22_X1  g232(.A1(new_n422), .A2(KEYINPUT82), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n345), .B(new_n414), .C1(new_n424), .C2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n430), .A2(new_n433), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n413), .B1(new_n422), .B2(KEYINPUT82), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n411), .A2(KEYINPUT4), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(new_n418), .A3(new_n420), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT82), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n443), .A3(new_n402), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n439), .A2(new_n440), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n345), .B1(new_n445), .B2(new_n414), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n437), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n414), .B1(new_n424), .B2(new_n434), .ZN(new_n448));
  INV_X1    g247(.A(new_n345), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(KEYINPUT6), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n341), .B1(new_n447), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT84), .B1(new_n322), .B2(KEYINPUT29), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT29), .B1(new_n319), .B2(new_n320), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT84), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n453), .A2(new_n400), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT85), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n457), .A2(new_n458), .A3(new_n377), .A4(new_n383), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n400), .B1(new_n454), .B2(new_n455), .ZN(new_n460));
  AOI211_X1 g259(.A(KEYINPUT84), .B(KEYINPUT29), .C1(new_n319), .C2(new_n320), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n377), .B(new_n383), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT85), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  AND2_X1   g263(.A1(G228gat), .A2(G233gat), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n382), .A2(new_n400), .A3(new_n375), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT29), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT86), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n321), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT29), .B1(new_n399), .B2(new_n400), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT86), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n466), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n406), .A2(new_n410), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n454), .A2(KEYINPUT3), .ZN(new_n476));
  OAI22_X1  g275(.A1(new_n475), .A2(new_n476), .B1(new_n321), .B2(new_n472), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n464), .A2(new_n474), .B1(new_n466), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G22gat), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT87), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n474), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n477), .A2(new_n466), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(G22gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G78gat), .B(G106gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT31), .B(G50gat), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n486), .B(new_n487), .Z(new_n488));
  NAND3_X1  g287(.A1(new_n483), .A2(KEYINPUT87), .A3(G22gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n484), .A2(KEYINPUT88), .ZN(new_n491));
  OR3_X1    g290(.A1(new_n478), .A2(KEYINPUT88), .A3(new_n479), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n488), .B1(new_n478), .B2(new_n479), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n308), .A2(new_n427), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n326), .A2(new_n398), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(G227gat), .A2(G233gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n499), .B(KEYINPUT64), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n503), .A2(KEYINPUT34), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT71), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n498), .A2(KEYINPUT71), .A3(new_n504), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n496), .A2(new_n497), .A3(new_n503), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT32), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT33), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(G15gat), .B(G43gat), .Z(new_n515));
  XNOR2_X1  g314(.A(G71gat), .B(G99gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n512), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n517), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n511), .B(KEYINPUT32), .C1(new_n513), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n510), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n508), .A2(new_n520), .A3(new_n518), .A4(new_n509), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n495), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT35), .B1(new_n452), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n448), .A2(new_n449), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n528), .A2(new_n436), .A3(new_n435), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n450), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n524), .B1(new_n490), .B2(new_n494), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT35), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .A4(new_n341), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n338), .B1(new_n337), .B2(KEYINPUT37), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT38), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n308), .A2(KEYINPUT74), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT74), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n326), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n327), .B1(new_n540), .B2(new_n324), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT37), .B1(new_n541), .B2(new_n321), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n310), .A2(new_n321), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n536), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n335), .B1(new_n535), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n322), .B1(new_n325), .B2(new_n328), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n546), .B1(new_n322), .B2(new_n310), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT37), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n255), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n337), .A2(KEYINPUT37), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n536), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n545), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(new_n529), .A3(new_n450), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT89), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n384), .A2(new_n401), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n432), .B1(new_n412), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT39), .B1(new_n429), .B2(new_n347), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT39), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n558), .A2(KEYINPUT40), .A3(new_n345), .A4(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT40), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n345), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n556), .A2(new_n557), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n414), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n442), .A2(new_n443), .A3(new_n402), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n567), .A2(new_n438), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n566), .B1(new_n568), .B2(new_n440), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n561), .B(new_n565), .C1(new_n569), .C2(new_n345), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n554), .B1(new_n570), .B2(new_n341), .ZN(new_n571));
  NOR3_X1   g370(.A1(new_n334), .A2(new_n331), .A3(new_n332), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(new_n339), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n558), .A2(new_n345), .A3(new_n560), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n448), .A2(new_n449), .B1(new_n574), .B2(new_n562), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n573), .A2(new_n575), .A3(KEYINPUT89), .A4(new_n561), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n553), .A2(new_n571), .A3(new_n495), .A4(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n495), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n452), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n524), .B(KEYINPUT36), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n577), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n252), .B1(new_n534), .B2(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G57gat), .B(G64gat), .Z(new_n584));
  INV_X1    g383(.A(KEYINPUT9), .ZN(new_n585));
  INV_X1    g384(.A(G71gat), .ZN(new_n586));
  INV_X1    g385(.A(G78gat), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G71gat), .B(G78gat), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n584), .A2(new_n590), .A3(new_n588), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT21), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(new_n394), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n592), .A2(new_n593), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT94), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT21), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(new_n214), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n599), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(G155gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(G183gat), .B(G211gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n604), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G99gat), .A2(G106gat), .ZN(new_n610));
  INV_X1    g409(.A(G85gat), .ZN(new_n611));
  INV_X1    g410(.A(G92gat), .ZN(new_n612));
  AOI22_X1  g411(.A1(KEYINPUT8), .A2(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT7), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(new_n611), .B2(new_n612), .ZN(new_n615));
  NAND3_X1  g414(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n613), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G99gat), .B(G106gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n617), .A2(new_n619), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n623), .B1(new_n229), .B2(new_n230), .ZN(new_n624));
  AND2_X1   g423(.A1(G232gat), .A2(G233gat), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n232), .A2(new_n622), .B1(KEYINPUT41), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(G190gat), .B(G218gat), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n625), .A2(KEYINPUT41), .ZN(new_n630));
  XNOR2_X1  g429(.A(G134gat), .B(G162gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n628), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n624), .A2(new_n633), .A3(new_n626), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n629), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n632), .B1(new_n629), .B2(new_n634), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n609), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT95), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n609), .A2(KEYINPUT95), .A3(new_n638), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n601), .A2(KEYINPUT10), .A3(new_n622), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n617), .A2(KEYINPUT96), .A3(new_n618), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n600), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n618), .B1(new_n617), .B2(KEYINPUT96), .ZN(new_n648));
  OAI22_X1  g447(.A1(new_n623), .A2(new_n600), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT98), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT97), .B(KEYINPUT10), .Z(new_n651));
  AND3_X1   g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n650), .B1(new_n649), .B2(new_n651), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n645), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(G230gat), .A2(G233gat), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n649), .A2(new_n655), .ZN(new_n659));
  XNOR2_X1  g458(.A(G120gat), .B(G148gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(G176gat), .B(G204gat), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n660), .B(new_n661), .Z(new_n662));
  NAND3_X1  g461(.A1(new_n654), .A2(KEYINPUT99), .A3(new_n655), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n658), .A2(new_n659), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n662), .ZN(new_n665));
  INV_X1    g464(.A(new_n645), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n649), .A2(new_n651), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT98), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n666), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n655), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n659), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n665), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n664), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n644), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n583), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n530), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g480(.A1(new_n678), .A2(new_n573), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT16), .B(G8gat), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT42), .Z(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(G8gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT100), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(G1325gat));
  OAI21_X1  g487(.A(G15gat), .B1(new_n677), .B2(new_n581), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n524), .A2(G15gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n689), .B1(new_n677), .B2(new_n690), .ZN(G1326gat));
  NOR2_X1   g490(.A1(new_n677), .A2(new_n495), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT43), .B(G22gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  INV_X1    g493(.A(new_n675), .ZN(new_n695));
  INV_X1    g494(.A(new_n609), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(new_n638), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n583), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n700), .A2(G29gat), .A3(new_n530), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT45), .Z(new_n702));
  NAND4_X1  g501(.A1(new_n577), .A2(new_n579), .A3(KEYINPUT101), .A4(new_n581), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n534), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n580), .B1(new_n452), .B2(new_n578), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT101), .B1(new_n705), .B2(new_n577), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n637), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n534), .A2(new_n582), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(KEYINPUT44), .A3(new_n637), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n248), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(G29gat), .B1(new_n715), .B2(new_n530), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n702), .A2(new_n716), .ZN(G1328gat));
  NOR3_X1   g516(.A1(new_n700), .A2(new_n341), .A3(new_n215), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT46), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n215), .B1(new_n715), .B2(new_n341), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(G1329gat));
  OAI21_X1  g520(.A(G43gat), .B1(new_n715), .B2(new_n581), .ZN(new_n722));
  NOR2_X1   g521(.A1(KEYINPUT103), .A2(KEYINPUT47), .ZN(new_n723));
  INV_X1    g522(.A(G43gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n699), .A2(new_n724), .A3(new_n525), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n725), .A2(KEYINPUT102), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(KEYINPUT102), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n723), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n722), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(KEYINPUT103), .A2(KEYINPUT47), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1330gat));
  NAND2_X1  g530(.A1(new_n578), .A2(G50gat), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n700), .A2(new_n495), .ZN(new_n733));
  OAI22_X1  g532(.A1(new_n715), .A2(new_n732), .B1(G50gat), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g534(.A(KEYINPUT101), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n582), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n737), .A2(new_n534), .A3(new_n703), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n644), .A2(new_n248), .A3(new_n695), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n679), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n573), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT49), .B(G64gat), .Z(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n744), .B2(new_n746), .ZN(G1333gat));
  NAND3_X1  g546(.A1(new_n741), .A2(G71gat), .A3(new_n580), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT104), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(new_n740), .B2(new_n524), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n586), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n740), .A2(new_n749), .A3(new_n524), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n748), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g553(.A1(new_n741), .A2(new_n578), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g555(.A1(new_n248), .A2(new_n609), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n675), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT105), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n712), .A2(new_n679), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n611), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n761), .B2(new_n760), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n637), .B(new_n757), .C1(new_n704), .C2(new_n706), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n738), .A2(KEYINPUT51), .A3(new_n637), .A4(new_n757), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n768), .A2(new_n611), .A3(new_n679), .A4(new_n675), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n763), .A2(new_n769), .ZN(G1336gat));
  NAND3_X1  g569(.A1(new_n712), .A2(new_n573), .A3(new_n759), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G92gat), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n695), .A2(G92gat), .A3(new_n341), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT52), .B1(new_n768), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n773), .B(KEYINPUT107), .ZN(new_n776));
  AOI22_X1  g575(.A1(new_n771), .A2(G92gat), .B1(new_n768), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(G1337gat));
  NAND3_X1  g578(.A1(new_n712), .A2(new_n580), .A3(new_n759), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G99gat), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n695), .A2(G99gat), .A3(new_n524), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT108), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n781), .A2(new_n784), .ZN(G1338gat));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787));
  OR3_X1    g586(.A1(new_n695), .A2(new_n495), .A3(G106gat), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT109), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n768), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n709), .A2(new_n578), .A3(new_n711), .A4(new_n759), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n790), .A2(KEYINPUT110), .B1(G106gat), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n789), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(new_n766), .B2(new_n767), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT110), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n787), .B1(new_n792), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n788), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT53), .B1(new_n768), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n791), .A2(G106gat), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n786), .B1(new_n797), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n800), .B1(new_n795), .B2(new_n794), .ZN(new_n804));
  INV_X1    g603(.A(new_n796), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT53), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n806), .A2(KEYINPUT111), .A3(new_n801), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n803), .A2(new_n807), .ZN(G1339gat));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n670), .A2(new_n657), .A3(new_n671), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT99), .B1(new_n654), .B2(new_n655), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n671), .B(new_n645), .C1(new_n652), .C2(new_n653), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT54), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n665), .B1(new_n656), .B2(KEYINPUT54), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n809), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n670), .B2(new_n671), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n658), .A2(new_n663), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n662), .B1(new_n672), .B2(new_n817), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(new_n820), .A3(KEYINPUT55), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n816), .A2(new_n248), .A3(new_n664), .A4(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n234), .A2(new_n208), .A3(new_n235), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n239), .B2(new_n241), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n205), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n675), .A2(new_n247), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n637), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n821), .A2(new_n664), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT55), .B1(new_n819), .B2(new_n820), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n247), .A2(new_n637), .A3(new_n825), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n696), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n643), .A2(new_n713), .A3(new_n695), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n526), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n834), .A2(new_n679), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n341), .ZN(new_n836));
  INV_X1    g635(.A(G113gat), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n836), .A2(new_n837), .A3(new_n252), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n835), .A2(KEYINPUT112), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n834), .A2(new_n679), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT112), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(new_n341), .A3(new_n248), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n838), .B1(new_n844), .B2(new_n837), .ZN(G1340gat));
  NOR3_X1   g644(.A1(new_n836), .A2(new_n390), .A3(new_n695), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n843), .A2(new_n341), .A3(new_n675), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(new_n390), .ZN(G1341gat));
  NAND4_X1  g647(.A1(new_n835), .A2(G127gat), .A3(new_n341), .A4(new_n609), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT113), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n843), .A2(new_n341), .A3(new_n609), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n394), .B2(new_n851), .ZN(G1342gat));
  NAND2_X1  g651(.A1(new_n341), .A2(new_n637), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT114), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(G134gat), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n839), .A2(new_n842), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT56), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT115), .ZN(new_n858));
  OAI21_X1  g657(.A(G134gat), .B1(new_n836), .B2(new_n638), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT56), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n839), .A2(new_n860), .A3(new_n842), .A4(new_n855), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n856), .A2(new_n863), .A3(KEYINPUT56), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n858), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n858), .A2(new_n862), .A3(KEYINPUT116), .A4(new_n864), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1343gat));
  NOR2_X1   g668(.A1(new_n580), .A2(new_n530), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n341), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n578), .A2(KEYINPUT57), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n821), .A2(new_n664), .ZN(new_n874));
  XNOR2_X1  g673(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n875), .B1(new_n814), .B2(new_n815), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n874), .B(new_n876), .C1(new_n250), .C2(new_n251), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n637), .B1(new_n877), .B2(new_n826), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n696), .B1(new_n878), .B2(new_n831), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n873), .B1(new_n879), .B2(new_n833), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n832), .A2(new_n833), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT57), .B1(new_n881), .B2(new_n578), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n872), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(G141gat), .B1(new_n883), .B2(new_n713), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n884), .A2(KEYINPUT118), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n884), .A2(KEYINPUT118), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n881), .A2(new_n578), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n887), .A2(new_n871), .ZN(new_n888));
  INV_X1    g687(.A(new_n252), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n359), .A3(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n885), .A2(new_n886), .A3(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT58), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n883), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n889), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n894), .B1(new_n896), .B2(G141gat), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI211_X1 g698(.A(KEYINPUT119), .B(new_n894), .C1(new_n896), .C2(G141gat), .ZN(new_n900));
  OAI22_X1  g699(.A1(new_n892), .A2(new_n893), .B1(new_n899), .B2(new_n900), .ZN(G1344gat));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n877), .A2(new_n826), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n638), .ZN(new_n906));
  INV_X1    g705(.A(new_n831), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n609), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n644), .A2(new_n889), .A3(new_n675), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n904), .B(new_n578), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n887), .A2(KEYINPUT57), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n675), .B1(new_n872), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n913), .B1(new_n912), .B2(new_n872), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n903), .B1(new_n915), .B2(G148gat), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n675), .B(new_n872), .C1(new_n880), .C2(new_n882), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n361), .A2(KEYINPUT59), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT120), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT120), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n917), .A2(new_n921), .A3(new_n918), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n916), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n888), .A2(new_n361), .A3(new_n675), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n902), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(new_n922), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n921), .B1(new_n917), .B2(new_n918), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g728(.A(KEYINPUT122), .B(new_n924), .C1(new_n929), .C2(new_n916), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n926), .A2(new_n930), .ZN(G1345gat));
  AOI21_X1  g730(.A(G155gat), .B1(new_n888), .B2(new_n609), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n609), .A2(G155gat), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT123), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n932), .B1(new_n895), .B2(new_n934), .ZN(G1346gat));
  OAI21_X1  g734(.A(G162gat), .B1(new_n883), .B2(new_n638), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n854), .A2(G162gat), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n870), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n936), .B1(new_n887), .B2(new_n938), .ZN(G1347gat));
  NOR2_X1   g738(.A1(new_n679), .A2(new_n341), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n834), .A2(new_n940), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n941), .A2(G169gat), .A3(new_n713), .ZN(new_n942));
  INV_X1    g741(.A(new_n941), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n889), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n942), .B1(G169gat), .B2(new_n944), .ZN(new_n945));
  XOR2_X1   g744(.A(new_n945), .B(KEYINPUT124), .Z(G1348gat));
  NOR2_X1   g745(.A1(new_n941), .A2(new_n695), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(new_n264), .ZN(G1349gat));
  NAND2_X1  g747(.A1(new_n943), .A2(new_n609), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(new_n277), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n289), .A2(new_n291), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(new_n951), .B2(new_n949), .ZN(new_n952));
  XOR2_X1   g751(.A(new_n952), .B(KEYINPUT60), .Z(G1350gat));
  NOR2_X1   g752(.A1(new_n941), .A2(new_n638), .ZN(new_n954));
  NAND2_X1  g753(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g755(.A(KEYINPUT61), .B(G190gat), .Z(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n954), .B2(new_n957), .ZN(G1351gat));
  NAND2_X1  g757(.A1(new_n940), .A2(new_n581), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n887), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g759(.A(KEYINPUT125), .B(G197gat), .Z(new_n961));
  NAND3_X1  g760(.A1(new_n960), .A2(new_n248), .A3(new_n961), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n910), .A2(new_n911), .ZN(new_n963));
  XOR2_X1   g762(.A(new_n959), .B(KEYINPUT126), .Z(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n965), .A2(new_n252), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n962), .B1(new_n966), .B2(new_n961), .ZN(G1352gat));
  OAI21_X1  g766(.A(G204gat), .B1(new_n965), .B2(new_n695), .ZN(new_n968));
  NOR4_X1   g767(.A1(new_n887), .A2(G204gat), .A3(new_n695), .A4(new_n959), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT62), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n968), .A2(new_n970), .ZN(G1353gat));
  INV_X1    g770(.A(G211gat), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n959), .A2(new_n696), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n972), .B1(new_n963), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT63), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n972), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n887), .B2(new_n976), .ZN(G1354gat));
  AOI21_X1  g776(.A(G218gat), .B1(new_n960), .B2(new_n637), .ZN(new_n978));
  INV_X1    g777(.A(new_n965), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n637), .A2(G218gat), .ZN(new_n980));
  XOR2_X1   g779(.A(new_n980), .B(KEYINPUT127), .Z(new_n981));
  AOI21_X1  g780(.A(new_n978), .B1(new_n979), .B2(new_n981), .ZN(G1355gat));
endmodule


