//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 0 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n539, new_n540, new_n541, new_n542, new_n543, new_n545,
    new_n547, new_n548, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n588,
    new_n589, new_n592, new_n594, new_n595, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT64), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT65), .Z(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  XNOR2_X1  g046(.A(new_n471), .B(KEYINPUT67), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT66), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n463), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n462), .A2(KEYINPUT66), .A3(KEYINPUT3), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n475), .A2(G137), .A3(new_n470), .A4(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n469), .A2(new_n473), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NAND3_X1  g054(.A1(new_n475), .A2(G2105), .A3(new_n476), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n475), .A2(new_n470), .A3(new_n476), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n490), .A2(new_n470), .A3(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n466), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n475), .A2(G138), .A3(new_n470), .A4(new_n476), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n475), .A2(G126), .A3(G2105), .A4(new_n476), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT68), .B(G114), .ZN(new_n497));
  OAI211_X1 g072(.A(G2104), .B(new_n496), .C1(new_n497), .C2(new_n470), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n494), .A2(new_n499), .ZN(G164));
  NAND2_X1  g075(.A1(G75), .A2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G62), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n501), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n511));
  XNOR2_X1  g086(.A(new_n511), .B(KEYINPUT69), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(G543), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n503), .A2(new_n505), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n512), .A2(new_n513), .A3(new_n517), .ZN(new_n518));
  OAI221_X1 g093(.A(new_n509), .B1(new_n514), .B2(new_n515), .C1(new_n516), .C2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND3_X1  g095(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n521));
  INV_X1    g096(.A(new_n514), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G51), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n512), .A2(G89), .A3(new_n513), .A4(new_n517), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n524), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n525), .B1(new_n524), .B2(new_n527), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n521), .B(new_n523), .C1(new_n528), .C2(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  INV_X1    g106(.A(new_n518), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G90), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n522), .A2(G52), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n510), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AOI22_X1  g113(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT71), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  AOI22_X1  g116(.A1(G43), .A2(new_n522), .B1(new_n532), .B2(G81), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  AND3_X1   g119(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G36), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n545), .A2(new_n548), .ZN(G188));
  INV_X1    g124(.A(G53), .ZN(new_n550));
  XOR2_X1   g125(.A(KEYINPUT72), .B(KEYINPUT9), .Z(new_n551));
  NOR3_X1   g126(.A1(new_n514), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT73), .ZN(new_n553));
  OAI21_X1  g128(.A(KEYINPUT9), .B1(new_n514), .B2(new_n550), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n506), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n532), .A2(G91), .B1(G651), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n555), .A2(new_n559), .ZN(G299));
  OAI21_X1  g135(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n561));
  INV_X1    g136(.A(G49), .ZN(new_n562));
  INV_X1    g137(.A(G87), .ZN(new_n563));
  OAI221_X1 g138(.A(new_n561), .B1(new_n514), .B2(new_n562), .C1(new_n563), .C2(new_n518), .ZN(G288));
  NAND2_X1  g139(.A1(G73), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G61), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n506), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  INV_X1    g143(.A(G48), .ZN(new_n569));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  OAI221_X1 g145(.A(new_n568), .B1(new_n514), .B2(new_n569), .C1(new_n570), .C2(new_n518), .ZN(G305));
  XOR2_X1   g146(.A(KEYINPUT75), .B(G47), .Z(new_n572));
  AOI22_X1  g147(.A1(G85), .A2(new_n532), .B1(new_n522), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT74), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n573), .B1(new_n510), .B2(new_n575), .ZN(G290));
  NAND2_X1  g151(.A1(G301), .A2(G868), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n532), .A2(G92), .ZN(new_n578));
  XOR2_X1   g153(.A(new_n578), .B(KEYINPUT10), .Z(new_n579));
  AOI22_X1  g154(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n580));
  XOR2_X1   g155(.A(new_n580), .B(KEYINPUT76), .Z(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n522), .A2(G54), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n579), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n577), .B1(new_n585), .B2(G868), .ZN(G284));
  OAI21_X1  g161(.A(new_n577), .B1(new_n585), .B2(G868), .ZN(G321));
  NAND2_X1  g162(.A1(G286), .A2(G868), .ZN(new_n588));
  INV_X1    g163(.A(G299), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n589), .B2(G868), .ZN(G297));
  OAI21_X1  g165(.A(new_n588), .B1(new_n589), .B2(G868), .ZN(G280));
  XOR2_X1   g166(.A(KEYINPUT77), .B(G559), .Z(new_n592));
  OAI21_X1  g167(.A(new_n585), .B1(G860), .B2(new_n592), .ZN(G148));
  NAND2_X1  g168(.A1(new_n585), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G868), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(G868), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g171(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g172(.A1(new_n481), .A2(G123), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n484), .A2(G135), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n470), .A2(G111), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n462), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI221_X1 g177(.A(new_n602), .B1(new_n601), .B2(new_n600), .C1(G99), .C2(G2105), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n598), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(G2096), .Z(new_n605));
  NAND3_X1  g180(.A1(new_n472), .A2(new_n463), .A3(new_n465), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  XOR2_X1   g182(.A(KEYINPUT78), .B(G2100), .Z(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT13), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n607), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n605), .A2(new_n610), .ZN(G156));
  XNOR2_X1  g186(.A(KEYINPUT15), .B(G2430), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2435), .ZN(new_n613));
  XOR2_X1   g188(.A(G2427), .B(G2438), .Z(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(KEYINPUT14), .ZN(new_n616));
  XNOR2_X1  g191(.A(G2451), .B(G2454), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT80), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT16), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n616), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(G2443), .B(G2446), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(G1341), .B(G1348), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n622), .B(new_n623), .Z(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G14), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(G401));
  XOR2_X1   g201(.A(G2084), .B(G2090), .Z(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(G2067), .B(G2678), .Z(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n630), .A2(new_n631), .A3(KEYINPUT17), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT18), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G2072), .B(G2078), .Z(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n630), .B2(KEYINPUT18), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n634), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2096), .B(G2100), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(G227));
  XNOR2_X1  g214(.A(G1971), .B(G1976), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT19), .ZN(new_n641));
  XOR2_X1   g216(.A(G1956), .B(G2474), .Z(new_n642));
  XOR2_X1   g217(.A(G1961), .B(G1966), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n641), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n642), .A2(new_n643), .ZN(new_n647));
  AOI22_X1  g222(.A1(new_n645), .A2(KEYINPUT20), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n649), .A2(new_n641), .A3(new_n644), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n648), .B(new_n650), .C1(KEYINPUT20), .C2(new_n645), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT81), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n651), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1991), .B(G1996), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1981), .B(G1986), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n656), .B(new_n657), .Z(G229));
  OAI21_X1  g233(.A(KEYINPUT90), .B1(G29), .B2(G33), .ZN(new_n659));
  OR3_X1    g234(.A1(KEYINPUT90), .A2(G29), .A3(G33), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n484), .A2(G139), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT25), .Z(new_n663));
  NAND2_X1  g238(.A1(G115), .A2(G2104), .ZN(new_n664));
  INV_X1    g239(.A(G127), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n664), .B1(new_n466), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT91), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n661), .B(new_n663), .C1(new_n667), .C2(new_n470), .ZN(new_n668));
  INV_X1    g243(.A(G29), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n659), .B(new_n660), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT92), .B(G2072), .Z(new_n671));
  XOR2_X1   g246(.A(new_n670), .B(new_n671), .Z(new_n672));
  INV_X1    g247(.A(G16), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n585), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(G4), .B2(new_n673), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT88), .B(G1348), .Z(new_n676));
  OR2_X1    g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n673), .A2(G19), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(new_n543), .B2(new_n673), .ZN(new_n679));
  AOI22_X1  g254(.A1(new_n675), .A2(new_n676), .B1(G1341), .B2(new_n679), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(G1341), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n669), .A2(G26), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n481), .A2(G128), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n484), .A2(G140), .ZN(new_n684));
  OR2_X1    g259(.A1(G104), .A2(G2105), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n685), .B(G2104), .C1(G116), .C2(new_n470), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n683), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n682), .B1(new_n688), .B2(new_n669), .ZN(new_n689));
  MUX2_X1   g264(.A(new_n682), .B(new_n689), .S(KEYINPUT28), .Z(new_n690));
  INV_X1    g265(.A(G2067), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NAND4_X1  g267(.A1(new_n677), .A2(new_n680), .A3(new_n681), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT89), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n673), .A2(G20), .ZN(new_n695));
  OAI211_X1 g270(.A(KEYINPUT23), .B(new_n695), .C1(new_n589), .C2(new_n673), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(KEYINPUT23), .B2(new_n695), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT98), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(G1956), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(G1956), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n669), .A2(G35), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G162), .B2(new_n669), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT97), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT29), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(G2090), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n673), .A2(G5), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G171), .B2(new_n673), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT96), .Z(new_n708));
  INV_X1    g283(.A(G1961), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n704), .A2(G2090), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n705), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n708), .A2(new_n709), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n669), .A2(G32), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n481), .A2(G129), .B1(G105), .B2(new_n472), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT26), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n484), .A2(G141), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n715), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT95), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n714), .B1(new_n724), .B2(new_n669), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT27), .B(G1996), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT31), .B(G11), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT24), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n669), .B1(new_n729), .B2(G34), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT93), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(G34), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(KEYINPUT93), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n478), .B2(new_n669), .ZN(new_n735));
  INV_X1    g310(.A(G2084), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT94), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n669), .A2(G27), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G164), .B2(new_n669), .ZN(new_n740));
  INV_X1    g315(.A(G2078), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G28), .ZN(new_n743));
  AOI21_X1  g318(.A(G29), .B1(new_n743), .B2(KEYINPUT30), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(KEYINPUT30), .B2(new_n743), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n604), .B2(new_n669), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n736), .B2(new_n735), .ZN(new_n747));
  AND4_X1   g322(.A1(new_n728), .A2(new_n738), .A3(new_n742), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n673), .A2(G21), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G168), .B2(new_n673), .ZN(new_n750));
  INV_X1    g325(.A(G1966), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n727), .A2(new_n748), .A3(new_n752), .ZN(new_n753));
  NOR3_X1   g328(.A1(new_n712), .A2(new_n713), .A3(new_n753), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n694), .A2(new_n699), .A3(new_n700), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n673), .A2(G22), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G166), .B2(new_n673), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1971), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n673), .A2(G23), .ZN(new_n759));
  INV_X1    g334(.A(G288), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(new_n673), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT33), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n758), .B1(G1976), .B2(new_n763), .ZN(new_n764));
  MUX2_X1   g339(.A(G6), .B(G305), .S(G16), .Z(new_n765));
  XOR2_X1   g340(.A(KEYINPUT32), .B(G1981), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT85), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n765), .B(new_n767), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n764), .B(new_n768), .C1(G1976), .C2(new_n763), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT86), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT84), .B(KEYINPUT34), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n669), .A2(G25), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n484), .A2(G131), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(KEYINPUT82), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(KEYINPUT82), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n776), .A2(new_n777), .B1(G119), .B2(new_n481), .ZN(new_n778));
  OR2_X1    g353(.A1(G95), .A2(G2105), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n779), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n774), .B1(new_n781), .B2(new_n669), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT83), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT35), .B(G1991), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n771), .A2(new_n772), .ZN(new_n786));
  MUX2_X1   g361(.A(G24), .B(G290), .S(G16), .Z(new_n787));
  INV_X1    g362(.A(G1986), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n773), .A2(new_n785), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n790), .A2(KEYINPUT87), .A3(KEYINPUT36), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n786), .A2(new_n789), .ZN(new_n792));
  NAND2_X1  g367(.A1(KEYINPUT87), .A2(KEYINPUT36), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n792), .A2(new_n793), .A3(new_n785), .A4(new_n773), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n672), .B(new_n755), .C1(new_n791), .C2(new_n794), .ZN(G311));
  AOI21_X1  g370(.A(new_n755), .B1(new_n791), .B2(new_n794), .ZN(new_n796));
  INV_X1    g371(.A(new_n672), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(G150));
  NAND2_X1  g373(.A1(new_n532), .A2(G93), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n522), .A2(G55), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n799), .B(new_n800), .C1(new_n510), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(G860), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT37), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n585), .A2(G559), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT38), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n543), .A2(new_n802), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n543), .A2(new_n802), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT39), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n806), .B(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n804), .B1(new_n811), .B2(G860), .ZN(G145));
  XNOR2_X1  g387(.A(new_n723), .B(new_n668), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(new_n687), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n815));
  INV_X1    g390(.A(new_n492), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT99), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n499), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n495), .A2(new_n498), .A3(KEYINPUT99), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n813), .A2(new_n687), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n814), .A2(new_n817), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  AND3_X1   g398(.A1(new_n495), .A2(KEYINPUT99), .A3(new_n498), .ZN(new_n824));
  AOI21_X1  g399(.A(KEYINPUT99), .B1(new_n495), .B2(new_n498), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n817), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n813), .A2(new_n687), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n813), .A2(new_n687), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n823), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n781), .A2(new_n607), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n481), .A2(G130), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n484), .A2(G142), .ZN(new_n833));
  OR2_X1    g408(.A1(G106), .A2(G2105), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n834), .B(G2104), .C1(G118), .C2(new_n470), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n832), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n778), .A2(new_n780), .ZN(new_n838));
  INV_X1    g413(.A(new_n607), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AND3_X1   g415(.A1(new_n831), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n837), .B1(new_n831), .B2(new_n840), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(KEYINPUT100), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n841), .B2(new_n842), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n830), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n823), .A2(new_n829), .ZN(new_n849));
  INV_X1    g424(.A(new_n847), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT101), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT101), .ZN(new_n852));
  NOR3_X1   g427(.A1(new_n830), .A2(new_n847), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n848), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n604), .B(new_n478), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n488), .ZN(new_n856));
  AOI21_X1  g431(.A(G37), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(KEYINPUT102), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(new_n830), .B2(new_n843), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(KEYINPUT102), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n859), .B(new_n860), .C1(new_n851), .C2(new_n853), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g438(.A(G299), .B(new_n584), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT103), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n594), .B(new_n809), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OR3_X1    g442(.A1(new_n864), .A2(KEYINPUT104), .A3(KEYINPUT41), .ZN(new_n868));
  XOR2_X1   g443(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n864), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(KEYINPUT104), .B1(new_n864), .B2(KEYINPUT41), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n867), .B1(new_n872), .B2(new_n866), .ZN(new_n873));
  XNOR2_X1  g448(.A(G290), .B(new_n760), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n874), .A2(KEYINPUT106), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(KEYINPUT106), .ZN(new_n876));
  XOR2_X1   g451(.A(G303), .B(G305), .Z(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(KEYINPUT42), .Z(new_n881));
  OR2_X1    g456(.A1(new_n873), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n873), .A2(new_n881), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n883), .A3(G868), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT107), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(G868), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n802), .A2(new_n887), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n886), .B1(new_n889), .B2(new_n885), .ZN(G295));
  OAI21_X1  g465(.A(new_n886), .B1(new_n889), .B2(new_n885), .ZN(G331));
  NAND3_X1  g466(.A1(new_n807), .A2(G301), .A3(new_n808), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(G301), .B1(new_n807), .B2(new_n808), .ZN(new_n894));
  OAI21_X1  g469(.A(G286), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n894), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(G168), .A3(new_n892), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n868), .A2(new_n898), .A3(new_n870), .A4(new_n871), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n895), .A2(new_n897), .A3(new_n864), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n880), .ZN(new_n902));
  AOI21_X1  g477(.A(G37), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n864), .A2(KEYINPUT41), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n898), .B(new_n904), .C1(new_n864), .C2(new_n869), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n905), .B(new_n880), .C1(new_n865), .C2(new_n898), .ZN(new_n906));
  XOR2_X1   g481(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n903), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT109), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n899), .A2(new_n880), .A3(new_n900), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n903), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n907), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n903), .A2(KEYINPUT109), .A3(new_n906), .A4(new_n908), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n911), .A2(new_n914), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n913), .A2(new_n907), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n919), .B1(new_n903), .B2(new_n906), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT44), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n917), .A2(new_n921), .ZN(G397));
  INV_X1    g497(.A(G1384), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n826), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n469), .A2(new_n473), .A3(G40), .A4(new_n477), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n928), .A2(G1996), .A3(new_n723), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT110), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n687), .B(new_n691), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n723), .B2(G1996), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n930), .B1(new_n928), .B2(new_n932), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n838), .A2(new_n784), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n838), .A2(new_n784), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n928), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n928), .ZN(new_n937));
  XNOR2_X1  g512(.A(G290), .B(new_n788), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n933), .B(new_n936), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G8), .ZN(new_n940));
  INV_X1    g515(.A(new_n927), .ZN(new_n941));
  OAI211_X1 g516(.A(KEYINPUT45), .B(new_n923), .C1(new_n494), .C2(new_n499), .ZN(new_n942));
  AOI21_X1  g517(.A(G1384), .B1(new_n821), .B2(new_n817), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n941), .B(new_n942), .C1(new_n943), .C2(KEYINPUT45), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n751), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT50), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n826), .A2(new_n946), .A3(new_n923), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n923), .B1(new_n494), .B2(new_n499), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT50), .ZN(new_n949));
  XNOR2_X1  g524(.A(KEYINPUT116), .B(G2084), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n947), .A2(new_n941), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n940), .B1(new_n945), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(KEYINPUT113), .B(G8), .ZN(new_n953));
  NAND2_X1  g528(.A1(G286), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT51), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT51), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n947), .A2(new_n941), .A3(new_n949), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n960), .A2(new_n950), .B1(new_n944), .B2(new_n751), .ZN(new_n961));
  INV_X1    g536(.A(new_n953), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n956), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n961), .A2(new_n954), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT121), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT121), .ZN(new_n968));
  AOI211_X1 g543(.A(new_n968), .B(new_n965), .C1(new_n956), .C2(new_n963), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT62), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT45), .B1(new_n826), .B2(new_n923), .ZN(new_n971));
  INV_X1    g546(.A(new_n942), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n971), .A2(new_n927), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n951), .B1(new_n973), .B2(G1966), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n958), .B1(new_n974), .B2(new_n953), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n954), .B1(new_n961), .B2(new_n940), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n975), .B1(new_n976), .B2(KEYINPUT51), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n968), .B1(new_n977), .B2(new_n965), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT62), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n964), .A2(KEYINPUT121), .A3(new_n966), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n826), .A2(KEYINPUT45), .A3(new_n923), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n927), .B1(new_n948), .B2(new_n925), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1971), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G2090), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n960), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n984), .A2(KEYINPUT111), .A3(new_n985), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n988), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(G303), .A2(G8), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT55), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n992), .A2(G8), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT112), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n992), .A2(new_n998), .A3(G8), .A4(new_n995), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n943), .A2(new_n941), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1002), .A2(new_n962), .ZN(new_n1003));
  NAND2_X1  g578(.A1(G305), .A2(G1981), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n568), .B1(new_n518), .B2(new_n570), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n514), .A2(new_n569), .ZN(new_n1006));
  OR3_X1    g581(.A1(new_n1005), .A2(new_n1006), .A3(G1981), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1004), .A2(new_n1007), .A3(KEYINPUT49), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1012));
  OAI221_X1 g587(.A(new_n1003), .B1(KEYINPUT49), .B2(new_n1008), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1976), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1003), .B1(new_n1014), .B2(G288), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT52), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT52), .B1(G288), .B2(new_n1014), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1003), .B(new_n1017), .C1(new_n1014), .C2(G288), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1013), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(KEYINPUT115), .B(new_n941), .C1(new_n943), .C2(new_n946), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n946), .B1(new_n826), .B2(new_n923), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1021), .B1(new_n1022), .B2(new_n927), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1020), .B(new_n1023), .C1(KEYINPUT50), .C2(new_n948), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n986), .B1(new_n1024), .B2(G2090), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n953), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n994), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1000), .A2(new_n1019), .A3(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n982), .A2(new_n983), .A3(new_n741), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(G1961), .B2(new_n960), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n926), .A2(KEYINPUT53), .A3(new_n741), .A4(new_n941), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1033), .A2(new_n972), .ZN(new_n1034));
  OAI21_X1  g609(.A(G171), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n970), .A2(new_n981), .A3(new_n1028), .A4(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1000), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1013), .A2(new_n1014), .A3(new_n760), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n1007), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1038), .A2(new_n1019), .B1(new_n1040), .B2(new_n1003), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n961), .A2(G286), .A3(new_n962), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1000), .A2(new_n1019), .A3(new_n1027), .A4(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT63), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n992), .A2(G8), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1044), .B1(new_n1046), .B2(new_n994), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1000), .A2(new_n1019), .A3(new_n1042), .A4(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1037), .A2(new_n1041), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT124), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n947), .A2(new_n941), .A3(new_n949), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1030), .A2(new_n1029), .B1(new_n1052), .B2(new_n709), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1053), .B(G301), .C1(new_n972), .C2(new_n1033), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT123), .ZN(new_n1055));
  INV_X1    g630(.A(new_n982), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1055), .B1(new_n1033), .B2(new_n1056), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n971), .A2(new_n1030), .A3(new_n927), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1058), .A2(KEYINPUT123), .A3(new_n741), .A4(new_n982), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1057), .A2(new_n1053), .A3(new_n1059), .ZN(new_n1060));
  OAI211_X1 g635(.A(KEYINPUT54), .B(new_n1054), .C1(new_n1060), .C2(G301), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n967), .B2(new_n969), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1057), .A2(new_n1059), .A3(new_n1053), .A4(G301), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n1035), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1000), .A2(new_n1066), .A3(new_n1027), .A4(new_n1019), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1051), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1068));
  XOR2_X1   g643(.A(G299), .B(KEYINPUT57), .Z(new_n1069));
  INV_X1    g644(.A(G1956), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1024), .A2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT56), .B(G2072), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n982), .A2(new_n983), .A3(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1069), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1348), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1002), .A2(new_n691), .B1(new_n1052), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(new_n584), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1079), .A2(new_n1069), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1074), .A2(KEYINPUT61), .ZN(new_n1081));
  XOR2_X1   g656(.A(KEYINPUT58), .B(G1341), .Z(new_n1082));
  NAND2_X1  g657(.A1(new_n1001), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT117), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n984), .A2(G1996), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1001), .A2(new_n1086), .A3(new_n1082), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n1090));
  NAND4_X1  g665(.A1(new_n1088), .A2(new_n1089), .A3(new_n543), .A4(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT60), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1076), .A2(new_n585), .A3(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1088), .A2(new_n543), .A3(new_n1090), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1088), .A2(new_n543), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n1097));
  OAI211_X1 g672(.A(KEYINPUT119), .B(new_n1095), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1076), .A2(new_n584), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT60), .B1(new_n1099), .B2(new_n1077), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1081), .A2(new_n1094), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT61), .B1(new_n1074), .B2(KEYINPUT120), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1078), .B(new_n1080), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  AND4_X1   g678(.A1(new_n1000), .A2(new_n1066), .A3(new_n1027), .A4(new_n1019), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n978), .A2(new_n980), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1104), .A2(KEYINPUT124), .A3(new_n1105), .A4(new_n1061), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1068), .A2(new_n1103), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n939), .B1(new_n1050), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n937), .A2(G1996), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1109), .B(KEYINPUT46), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n937), .B1(new_n724), .B2(new_n931), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1112), .B(KEYINPUT47), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n933), .A2(new_n935), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n688), .A2(new_n691), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n937), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n937), .A2(G290), .A3(G1986), .ZN(new_n1117));
  XOR2_X1   g692(.A(new_n1117), .B(KEYINPUT48), .Z(new_n1118));
  AND3_X1   g693(.A1(new_n933), .A2(new_n936), .A3(new_n1118), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1113), .A2(new_n1116), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT125), .B1(new_n1108), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n939), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1068), .A2(new_n1103), .A3(new_n1106), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1037), .A2(new_n1049), .A3(new_n1041), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1126), .A2(new_n1127), .A3(new_n1120), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1122), .A2(new_n1128), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g704(.A(G227), .ZN(new_n1131));
  NAND3_X1  g705(.A1(new_n625), .A2(G319), .A3(new_n1131), .ZN(new_n1132));
  AOI22_X1  g706(.A1(new_n857), .A2(new_n861), .B1(KEYINPUT126), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g707(.A1(new_n911), .A2(new_n914), .A3(new_n916), .ZN(new_n1134));
  NOR2_X1   g708(.A1(new_n1132), .A2(KEYINPUT126), .ZN(new_n1135));
  NOR2_X1   g709(.A1(new_n1135), .A2(G229), .ZN(new_n1136));
  AND3_X1   g710(.A1(new_n1133), .A2(new_n1134), .A3(new_n1136), .ZN(G308));
  NAND3_X1  g711(.A1(new_n1133), .A2(new_n1134), .A3(new_n1136), .ZN(G225));
endmodule


