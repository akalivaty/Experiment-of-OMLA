

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773;

  XNOR2_X1 U371 ( .A(n622), .B(n451), .ZN(n725) );
  BUF_X1 U372 ( .A(n700), .Z(n349) );
  NOR2_X1 U373 ( .A1(n436), .A2(n428), .ZN(n683) );
  NOR2_X1 U374 ( .A1(n592), .A2(n591), .ZN(n688) );
  XNOR2_X1 U375 ( .A(n557), .B(n556), .ZN(n348) );
  OR2_X1 U376 ( .A1(n737), .A2(G902), .ZN(n534) );
  OR2_X1 U377 ( .A1(G902), .A2(G237), .ZN(n514) );
  XOR2_X1 U378 ( .A(KEYINPUT8), .B(n528), .Z(n564) );
  XOR2_X2 U379 ( .A(G140), .B(G131), .Z(n554) );
  XNOR2_X2 U380 ( .A(n593), .B(KEYINPUT102), .ZN(n642) );
  XNOR2_X1 U381 ( .A(n348), .B(n431), .ZN(n657) );
  NOR2_X1 U382 ( .A1(G953), .A2(G237), .ZN(n543) );
  AND2_X1 U383 ( .A1(G898), .A2(G953), .ZN(n497) );
  XNOR2_X1 U384 ( .A(G110), .B(G140), .ZN(n527) );
  INV_X1 U385 ( .A(G953), .ZN(n739) );
  XNOR2_X1 U386 ( .A(n574), .B(n573), .ZN(n585) );
  AND2_X2 U387 ( .A1(n383), .A2(n392), .ZN(n390) );
  OR2_X2 U388 ( .A1(n526), .A2(G902), .ZN(n468) );
  NOR2_X1 U389 ( .A1(n621), .A2(n370), .ZN(n628) );
  AND2_X2 U390 ( .A1(n418), .A2(n747), .ZN(n419) );
  XNOR2_X2 U391 ( .A(n510), .B(n500), .ZN(n568) );
  OR2_X1 U392 ( .A1(n404), .A2(n651), .ZN(n353) );
  AND2_X1 U393 ( .A1(n403), .A2(n488), .ZN(n401) );
  NAND2_X1 U394 ( .A1(n485), .A2(n487), .ZN(n484) );
  AND2_X1 U395 ( .A1(n411), .A2(n409), .ZN(n408) );
  INV_X1 U396 ( .A(KEYINPUT16), .ZN(n442) );
  NAND2_X1 U397 ( .A1(n401), .A2(n400), .ZN(n395) );
  INV_X1 U398 ( .A(n484), .ZN(n386) );
  NAND2_X1 U399 ( .A1(n572), .A2(n633), .ZN(n574) );
  XNOR2_X1 U400 ( .A(n364), .B(n358), .ZN(n572) );
  NAND2_X1 U401 ( .A1(n425), .A2(n456), .ZN(n724) );
  NAND2_X2 U402 ( .A1(n408), .A2(n405), .ZN(n595) );
  NAND2_X1 U403 ( .A1(n407), .A2(n406), .ZN(n405) );
  XNOR2_X1 U404 ( .A(KEYINPUT69), .B(n608), .ZN(n619) );
  XNOR2_X1 U405 ( .A(n438), .B(n441), .ZN(n710) );
  NOR2_X1 U406 ( .A1(n698), .A2(n711), .ZN(n626) );
  XNOR2_X1 U407 ( .A(n618), .B(n440), .ZN(n609) );
  XNOR2_X1 U408 ( .A(n412), .B(n554), .ZN(n752) );
  XNOR2_X1 U409 ( .A(n483), .B(G137), .ZN(n412) );
  XNOR2_X1 U410 ( .A(n442), .B(G122), .ZN(n378) );
  XNOR2_X1 U411 ( .A(G146), .B(G125), .ZN(n509) );
  INV_X2 U412 ( .A(G128), .ZN(n427) );
  NOR2_X2 U413 ( .A1(n649), .A2(n691), .ZN(n758) );
  XNOR2_X2 U414 ( .A(n437), .B(n575), .ZN(n581) );
  XNOR2_X2 U415 ( .A(n630), .B(KEYINPUT40), .ZN(n773) );
  XNOR2_X1 U416 ( .A(n631), .B(KEYINPUT46), .ZN(n403) );
  XNOR2_X1 U417 ( .A(n446), .B(KEYINPUT73), .ZN(n402) );
  INV_X1 U418 ( .A(KEYINPUT86), .ZN(n489) );
  XOR2_X1 U419 ( .A(KEYINPUT4), .B(KEYINPUT64), .Z(n507) );
  INV_X1 U420 ( .A(KEYINPUT68), .ZN(n483) );
  XNOR2_X1 U421 ( .A(n515), .B(KEYINPUT79), .ZN(n516) );
  XNOR2_X1 U422 ( .A(n445), .B(n553), .ZN(n556) );
  OR2_X1 U423 ( .A1(n667), .A2(G902), .ZN(n479) );
  XNOR2_X1 U424 ( .A(G902), .B(KEYINPUT15), .ZN(n650) );
  XNOR2_X1 U425 ( .A(n374), .B(n373), .ZN(n613) );
  INV_X1 U426 ( .A(KEYINPUT108), .ZN(n373) );
  NAND2_X1 U427 ( .A1(n609), .A2(n375), .ZN(n374) );
  AND2_X1 U428 ( .A1(n685), .A2(n619), .ZN(n375) );
  NAND2_X1 U429 ( .A1(n724), .A2(n595), .ZN(n364) );
  XNOR2_X1 U430 ( .A(KEYINPUT22), .B(KEYINPUT65), .ZN(n575) );
  NAND2_X1 U431 ( .A1(n486), .A2(KEYINPUT48), .ZN(n394) );
  AND2_X1 U432 ( .A1(n402), .A2(n646), .ZN(n400) );
  XNOR2_X1 U433 ( .A(G113), .B(G116), .ZN(n362) );
  XNOR2_X1 U434 ( .A(n466), .B(n422), .ZN(n421) );
  INV_X1 U435 ( .A(KEYINPUT66), .ZN(n422) );
  INV_X1 U436 ( .A(G146), .ZN(n540) );
  INV_X1 U437 ( .A(n509), .ZN(n382) );
  XNOR2_X1 U438 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n473) );
  INV_X1 U439 ( .A(KEYINPUT70), .ZN(n430) );
  INV_X1 U440 ( .A(n627), .ZN(n371) );
  INV_X1 U441 ( .A(KEYINPUT13), .ZN(n559) );
  XNOR2_X1 U442 ( .A(G128), .B(KEYINPUT24), .ZN(n481) );
  XNOR2_X1 U443 ( .A(G119), .B(KEYINPUT23), .ZN(n482) );
  XNOR2_X1 U444 ( .A(n527), .B(n412), .ZN(n381) );
  NAND2_X1 U445 ( .A1(n761), .A2(G234), .ZN(n528) );
  AND2_X1 U446 ( .A1(n453), .A2(n454), .ZN(n425) );
  XNOR2_X1 U447 ( .A(n623), .B(KEYINPUT111), .ZN(n451) );
  NAND2_X1 U448 ( .A1(n714), .A2(n712), .ZN(n622) );
  XNOR2_X1 U449 ( .A(n696), .B(KEYINPUT91), .ZN(n615) );
  NAND2_X1 U450 ( .A1(n613), .A2(n476), .ZN(n475) );
  INV_X1 U451 ( .A(KEYINPUT104), .ZN(n398) );
  XNOR2_X1 U452 ( .A(n571), .B(KEYINPUT107), .ZN(n633) );
  NAND2_X1 U453 ( .A1(n424), .A2(n423), .ZN(n436) );
  AND2_X1 U454 ( .A1(n524), .A2(n410), .ZN(n406) );
  XOR2_X1 U455 ( .A(KEYINPUT25), .B(KEYINPUT77), .Z(n532) );
  INV_X1 U456 ( .A(KEYINPUT6), .ZN(n440) );
  AND2_X2 U457 ( .A1(n420), .A2(n353), .ZN(n369) );
  NAND2_X1 U458 ( .A1(n658), .A2(n660), .ZN(n496) );
  OR2_X1 U459 ( .A1(n658), .A2(n660), .ZN(n495) );
  AND2_X1 U460 ( .A1(n492), .A2(n738), .ZN(n416) );
  NAND2_X1 U461 ( .A1(n494), .A2(n493), .ZN(n492) );
  OR2_X1 U462 ( .A1(n658), .A2(KEYINPUT59), .ZN(n493) );
  INV_X1 U463 ( .A(n692), .ZN(n487) );
  NAND2_X1 U464 ( .A1(n484), .A2(n393), .ZN(n392) );
  NOR2_X1 U465 ( .A1(n389), .A2(n388), .ZN(n387) );
  XNOR2_X1 U466 ( .A(KEYINPUT80), .B(n606), .ZN(n627) );
  XNOR2_X1 U467 ( .A(n552), .B(n351), .ZN(n445) );
  XOR2_X1 U468 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n552) );
  XNOR2_X1 U469 ( .A(KEYINPUT0), .B(KEYINPUT89), .ZN(n525) );
  XOR2_X1 U470 ( .A(KEYINPUT95), .B(KEYINPUT21), .Z(n537) );
  INV_X1 U471 ( .A(KEYINPUT71), .ZN(n470) );
  XNOR2_X1 U472 ( .A(KEYINPUT74), .B(KEYINPUT38), .ZN(n441) );
  INV_X1 U473 ( .A(n525), .ZN(n410) );
  OR2_X1 U474 ( .A1(n524), .A2(n410), .ZN(n409) );
  INV_X1 U475 ( .A(G469), .ZN(n490) );
  XNOR2_X1 U476 ( .A(n480), .B(n546), .ZN(n667) );
  XNOR2_X1 U477 ( .A(n396), .B(n542), .ZN(n480) );
  INV_X1 U478 ( .A(KEYINPUT84), .ZN(n434) );
  XNOR2_X1 U479 ( .A(G107), .B(G116), .ZN(n562) );
  XNOR2_X1 U480 ( .A(n432), .B(G122), .ZN(n563) );
  INV_X1 U481 ( .A(KEYINPUT9), .ZN(n432) );
  XOR2_X1 U482 ( .A(KEYINPUT101), .B(KEYINPUT7), .Z(n566) );
  XNOR2_X1 U483 ( .A(n511), .B(n512), .ZN(n376) );
  XNOR2_X1 U484 ( .A(n513), .B(n741), .ZN(n377) );
  NAND2_X1 U485 ( .A1(n747), .A2(n758), .ZN(n404) );
  XNOR2_X1 U486 ( .A(n570), .B(G478), .ZN(n592) );
  NOR2_X1 U487 ( .A1(G902), .A2(n657), .ZN(n561) );
  BUF_X1 U488 ( .A(n698), .Z(n367) );
  NAND2_X1 U489 ( .A1(n369), .A2(G472), .ZN(n671) );
  XNOR2_X1 U490 ( .A(n529), .B(n381), .ZN(n380) );
  NAND2_X1 U491 ( .A1(n369), .A2(G217), .ZN(n465) );
  NAND2_X1 U492 ( .A1(n369), .A2(G469), .ZN(n478) );
  XNOR2_X1 U493 ( .A(n652), .B(KEYINPUT57), .ZN(n477) );
  NAND2_X1 U494 ( .A1(n369), .A2(G210), .ZN(n664) );
  INV_X1 U495 ( .A(n736), .ZN(n738) );
  INV_X1 U496 ( .A(n436), .ZN(n638) );
  XNOR2_X1 U497 ( .A(n617), .B(KEYINPUT113), .ZN(n766) );
  INV_X1 U498 ( .A(KEYINPUT36), .ZN(n474) );
  INV_X1 U499 ( .A(KEYINPUT35), .ZN(n573) );
  XNOR2_X1 U500 ( .A(n399), .B(n398), .ZN(n397) );
  BUF_X1 U501 ( .A(n639), .Z(n428) );
  AND2_X2 U502 ( .A1(n591), .A2(n592), .ZN(n685) );
  XNOR2_X1 U503 ( .A(n732), .B(n450), .ZN(n735) );
  XNOR2_X1 U504 ( .A(n734), .B(n733), .ZN(n450) );
  NAND2_X1 U505 ( .A1(n415), .A2(n414), .ZN(n413) );
  XOR2_X1 U506 ( .A(KEYINPUT96), .B(n701), .Z(n350) );
  XOR2_X1 U507 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n351) );
  XOR2_X2 U508 ( .A(G104), .B(G107), .Z(n352) );
  OR2_X1 U509 ( .A1(n691), .A2(n650), .ZN(n354) );
  AND2_X1 U510 ( .A1(n452), .A2(n548), .ZN(n355) );
  XOR2_X1 U511 ( .A(n482), .B(n481), .Z(n356) );
  NOR2_X1 U512 ( .A1(n696), .A2(n695), .ZN(n357) );
  INV_X1 U513 ( .A(n548), .ZN(n455) );
  XOR2_X1 U514 ( .A(KEYINPUT34), .B(KEYINPUT78), .Z(n358) );
  XOR2_X1 U515 ( .A(KEYINPUT28), .B(KEYINPUT109), .Z(n359) );
  NAND2_X1 U516 ( .A1(n496), .A2(n495), .ZN(n360) );
  XNOR2_X1 U517 ( .A(n377), .B(n376), .ZN(n661) );
  OR2_X1 U518 ( .A1(n650), .A2(n651), .ZN(n361) );
  NAND2_X1 U519 ( .A1(n579), .A2(n578), .ZN(n363) );
  INV_X1 U520 ( .A(n362), .ZN(n505) );
  NAND2_X1 U521 ( .A1(n363), .A2(n580), .ZN(n769) );
  AND2_X2 U522 ( .A1(n429), .A2(n350), .ZN(n452) );
  XNOR2_X1 U523 ( .A(n555), .B(n365), .ZN(n431) );
  NAND2_X1 U524 ( .A1(n549), .A2(G214), .ZN(n365) );
  NAND2_X1 U525 ( .A1(n448), .A2(n366), .ZN(n637) );
  XNOR2_X1 U526 ( .A(n682), .B(KEYINPUT83), .ZN(n366) );
  INV_X1 U527 ( .A(n452), .ZN(n695) );
  NAND2_X1 U528 ( .A1(n452), .A2(n371), .ZN(n370) );
  AND2_X1 U529 ( .A1(n355), .A2(n609), .ZN(n457) );
  XNOR2_X1 U530 ( .A(n583), .B(KEYINPUT32), .ZN(n772) );
  NAND2_X1 U531 ( .A1(n439), .A2(n368), .ZN(n636) );
  XNOR2_X1 U532 ( .A(n626), .B(KEYINPUT30), .ZN(n368) );
  NAND2_X1 U533 ( .A1(n369), .A2(G475), .ZN(n659) );
  NAND2_X1 U534 ( .A1(n369), .A2(G478), .ZN(n732) );
  NAND2_X1 U535 ( .A1(n423), .A2(n452), .ZN(n372) );
  NOR2_X1 U536 ( .A1(n596), .A2(n372), .ZN(n676) );
  INV_X1 U537 ( .A(n685), .ZN(n629) );
  NAND2_X1 U538 ( .A1(n661), .A2(n650), .ZN(n517) );
  XNOR2_X2 U539 ( .A(n545), .B(n378), .ZN(n741) );
  XNOR2_X2 U540 ( .A(n740), .B(n430), .ZN(n513) );
  XNOR2_X1 U541 ( .A(n380), .B(n379), .ZN(n737) );
  XNOR2_X1 U542 ( .A(n356), .B(n755), .ZN(n379) );
  XNOR2_X1 U543 ( .A(n509), .B(KEYINPUT10), .ZN(n755) );
  INV_X1 U544 ( .A(n700), .ZN(n429) );
  XNOR2_X2 U545 ( .A(n534), .B(n533), .ZN(n700) );
  XNOR2_X1 U546 ( .A(n478), .B(n477), .ZN(n654) );
  XNOR2_X1 U547 ( .A(n465), .B(n464), .ZN(n463) );
  XNOR2_X1 U548 ( .A(n510), .B(n382), .ZN(n511) );
  XNOR2_X2 U549 ( .A(n427), .B(G143), .ZN(n510) );
  NOR2_X1 U550 ( .A1(n649), .A2(n354), .ZN(n418) );
  NAND2_X1 U551 ( .A1(n654), .A2(n738), .ZN(n656) );
  NAND2_X1 U552 ( .A1(n394), .A2(KEYINPUT85), .ZN(n388) );
  NAND2_X1 U553 ( .A1(n387), .A2(n386), .ZN(n385) );
  INV_X1 U554 ( .A(KEYINPUT85), .ZN(n393) );
  NAND2_X1 U555 ( .A1(n390), .A2(n385), .ZN(n649) );
  XNOR2_X1 U556 ( .A(n419), .B(n434), .ZN(n433) );
  NAND2_X1 U557 ( .A1(n391), .A2(n393), .ZN(n383) );
  NAND2_X1 U558 ( .A1(n384), .A2(n455), .ZN(n453) );
  NAND2_X1 U559 ( .A1(n609), .A2(n452), .ZN(n384) );
  INV_X1 U560 ( .A(n395), .ZN(n389) );
  NAND2_X1 U561 ( .A1(n395), .A2(n394), .ZN(n391) );
  XNOR2_X1 U562 ( .A(n396), .B(n540), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n396), .B(n753), .ZN(n754) );
  XNOR2_X2 U564 ( .A(n568), .B(n507), .ZN(n396) );
  NAND2_X1 U565 ( .A1(n581), .A2(n397), .ZN(n582) );
  NAND2_X1 U566 ( .A1(n615), .A2(n349), .ZN(n399) );
  XNOR2_X1 U567 ( .A(n766), .B(n489), .ZN(n488) );
  NAND2_X1 U568 ( .A1(n403), .A2(n402), .ZN(n486) );
  XNOR2_X1 U569 ( .A(n404), .B(n651), .ZN(n693) );
  INV_X1 U570 ( .A(n639), .ZN(n407) );
  NAND2_X1 U571 ( .A1(n639), .A2(n525), .ZN(n411) );
  NAND2_X1 U572 ( .A1(n472), .A2(n595), .ZN(n437) );
  XNOR2_X1 U573 ( .A(n413), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U574 ( .A1(n659), .A2(n416), .ZN(n414) );
  NAND2_X1 U575 ( .A1(n491), .A2(n417), .ZN(n415) );
  AND2_X1 U576 ( .A1(n360), .A2(n738), .ZN(n417) );
  XNOR2_X2 U577 ( .A(n459), .B(KEYINPUT45), .ZN(n747) );
  NAND2_X1 U578 ( .A1(n433), .A2(n361), .ZN(n420) );
  NAND2_X1 U579 ( .A1(n471), .A2(n421), .ZN(n461) );
  INV_X1 U580 ( .A(n621), .ZN(n423) );
  XNOR2_X1 U581 ( .A(n620), .B(n359), .ZN(n424) );
  XNOR2_X2 U582 ( .A(n621), .B(KEYINPUT1), .ZN(n696) );
  NAND2_X1 U583 ( .A1(n463), .A2(n738), .ZN(n462) );
  XNOR2_X1 U584 ( .A(n426), .B(n666), .ZN(G51) );
  NAND2_X1 U585 ( .A1(n665), .A2(n738), .ZN(n426) );
  XNOR2_X1 U586 ( .A(n473), .B(n506), .ZN(n508) );
  XNOR2_X1 U587 ( .A(n443), .B(KEYINPUT39), .ZN(n647) );
  NOR2_X1 U588 ( .A1(n647), .A2(n629), .ZN(n630) );
  XNOR2_X2 U589 ( .A(n352), .B(n499), .ZN(n740) );
  NAND2_X1 U590 ( .A1(n460), .A2(n602), .ZN(n459) );
  AND2_X1 U591 ( .A1(n712), .A2(n350), .ZN(n472) );
  INV_X1 U592 ( .A(n592), .ZN(n590) );
  XNOR2_X1 U593 ( .A(n567), .B(n566), .ZN(n449) );
  XNOR2_X1 U594 ( .A(n449), .B(n565), .ZN(n569) );
  NOR2_X2 U595 ( .A1(n636), .A2(n635), .ZN(n682) );
  BUF_X1 U596 ( .A(n634), .Z(n438) );
  XNOR2_X1 U597 ( .A(n502), .B(n469), .ZN(n526) );
  XNOR2_X1 U598 ( .A(n628), .B(KEYINPUT76), .ZN(n439) );
  XNOR2_X1 U599 ( .A(n475), .B(n474), .ZN(n616) );
  XNOR2_X2 U600 ( .A(n505), .B(n504), .ZN(n545) );
  NOR2_X2 U601 ( .A1(n636), .A2(n710), .ZN(n443) );
  NOR2_X2 U602 ( .A1(n773), .A2(n765), .ZN(n631) );
  NAND2_X1 U603 ( .A1(n444), .A2(n645), .ZN(n446) );
  XNOR2_X1 U604 ( .A(n637), .B(KEYINPUT81), .ZN(n444) );
  INV_X1 U605 ( .A(n642), .ZN(n715) );
  NAND2_X1 U606 ( .A1(n642), .A2(KEYINPUT47), .ZN(n632) );
  XNOR2_X2 U607 ( .A(n614), .B(n518), .ZN(n639) );
  NAND2_X2 U608 ( .A1(n634), .A2(n603), .ZN(n614) );
  XNOR2_X1 U609 ( .A(n584), .B(KEYINPUT88), .ZN(n471) );
  XNOR2_X1 U610 ( .A(n447), .B(n673), .ZN(G57) );
  NAND2_X1 U611 ( .A1(n672), .A2(n738), .ZN(n447) );
  XNOR2_X1 U612 ( .A(n632), .B(KEYINPUT82), .ZN(n448) );
  NAND2_X1 U613 ( .A1(n696), .A2(n455), .ZN(n454) );
  NAND2_X1 U614 ( .A1(n458), .A2(n457), .ZN(n456) );
  INV_X1 U615 ( .A(n696), .ZN(n458) );
  XNOR2_X1 U616 ( .A(n461), .B(n470), .ZN(n460) );
  XNOR2_X1 U617 ( .A(n462), .B(KEYINPUT123), .ZN(G66) );
  INV_X1 U618 ( .A(n737), .ZN(n464) );
  INV_X1 U619 ( .A(n585), .ZN(n768) );
  NAND2_X1 U620 ( .A1(n585), .A2(n467), .ZN(n466) );
  INV_X1 U621 ( .A(KEYINPUT44), .ZN(n467) );
  XNOR2_X2 U622 ( .A(n468), .B(n490), .ZN(n621) );
  XNOR2_X1 U623 ( .A(n501), .B(n513), .ZN(n469) );
  NOR2_X2 U624 ( .A1(n769), .A2(n772), .ZN(n584) );
  INV_X1 U625 ( .A(n614), .ZN(n476) );
  XNOR2_X2 U626 ( .A(n479), .B(n547), .ZN(n618) );
  NAND2_X2 U627 ( .A1(n588), .A2(n576), .ZN(n577) );
  OR2_X1 U628 ( .A1(n488), .A2(n646), .ZN(n485) );
  INV_X1 U629 ( .A(n659), .ZN(n491) );
  NAND2_X1 U630 ( .A1(n658), .A2(KEYINPUT59), .ZN(n494) );
  AND2_X1 U631 ( .A1(n739), .A2(G227), .ZN(n498) );
  INV_X1 U632 ( .A(KEYINPUT48), .ZN(n646) );
  XNOR2_X1 U633 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U634 ( .A(n752), .B(n498), .ZN(n501) );
  XNOR2_X1 U635 ( .A(n545), .B(n544), .ZN(n546) );
  NOR2_X1 U636 ( .A1(n523), .A2(n497), .ZN(n524) );
  INV_X1 U637 ( .A(G475), .ZN(n558) );
  INV_X1 U638 ( .A(G134), .ZN(n500) );
  XNOR2_X1 U639 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U640 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U641 ( .A(n661), .B(n662), .ZN(n663) );
  XNOR2_X1 U642 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U643 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U644 ( .A(G110), .B(G101), .ZN(n499) );
  XNOR2_X1 U645 ( .A(n526), .B(KEYINPUT58), .ZN(n652) );
  INV_X1 U646 ( .A(KEYINPUT19), .ZN(n518) );
  NAND2_X1 U647 ( .A1(G214), .A2(n514), .ZN(n503) );
  XNOR2_X1 U648 ( .A(KEYINPUT94), .B(n503), .ZN(n603) );
  XNOR2_X1 U649 ( .A(G119), .B(KEYINPUT3), .ZN(n504) );
  NAND2_X1 U650 ( .A1(G224), .A2(n739), .ZN(n506) );
  XNOR2_X1 U651 ( .A(n508), .B(n507), .ZN(n512) );
  NAND2_X1 U652 ( .A1(G210), .A2(n514), .ZN(n515) );
  XNOR2_X2 U653 ( .A(n517), .B(n516), .ZN(n634) );
  NAND2_X1 U654 ( .A1(G237), .A2(G234), .ZN(n519) );
  XNOR2_X1 U655 ( .A(n519), .B(KEYINPUT14), .ZN(n694) );
  INV_X2 U656 ( .A(G953), .ZN(n761) );
  OR2_X1 U657 ( .A1(n739), .A2(G902), .ZN(n520) );
  NAND2_X1 U658 ( .A1(n694), .A2(n520), .ZN(n522) );
  NOR2_X1 U659 ( .A1(G953), .A2(G952), .ZN(n521) );
  NOR2_X1 U660 ( .A1(n522), .A2(n521), .ZN(n605) );
  INV_X1 U661 ( .A(n605), .ZN(n523) );
  XOR2_X1 U662 ( .A(KEYINPUT106), .B(KEYINPUT33), .Z(n548) );
  NAND2_X1 U663 ( .A1(G221), .A2(n564), .ZN(n529) );
  NAND2_X1 U664 ( .A1(n650), .A2(G234), .ZN(n530) );
  XNOR2_X1 U665 ( .A(n530), .B(KEYINPUT20), .ZN(n535) );
  NAND2_X1 U666 ( .A1(n535), .A2(G217), .ZN(n531) );
  XNOR2_X1 U667 ( .A(n532), .B(n531), .ZN(n533) );
  NAND2_X1 U668 ( .A1(n535), .A2(G221), .ZN(n536) );
  XNOR2_X1 U669 ( .A(n537), .B(n536), .ZN(n701) );
  XNOR2_X1 U670 ( .A(KEYINPUT72), .B(G472), .ZN(n547) );
  XOR2_X1 U671 ( .A(KEYINPUT5), .B(G131), .Z(n539) );
  XNOR2_X1 U672 ( .A(G137), .B(G101), .ZN(n538) );
  XNOR2_X1 U673 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U674 ( .A(KEYINPUT75), .B(n543), .Z(n549) );
  NAND2_X1 U675 ( .A1(G210), .A2(n549), .ZN(n544) );
  XNOR2_X1 U676 ( .A(n755), .B(G104), .ZN(n557) );
  XOR2_X1 U677 ( .A(KEYINPUT100), .B(KEYINPUT12), .Z(n551) );
  XNOR2_X1 U678 ( .A(G113), .B(G122), .ZN(n550) );
  XNOR2_X1 U679 ( .A(n551), .B(n550), .ZN(n553) );
  XOR2_X1 U680 ( .A(n554), .B(G143), .Z(n555) );
  XNOR2_X2 U681 ( .A(n561), .B(n560), .ZN(n591) );
  XNOR2_X1 U682 ( .A(n563), .B(n562), .ZN(n567) );
  NAND2_X1 U683 ( .A1(G217), .A2(n564), .ZN(n565) );
  XOR2_X1 U684 ( .A(n568), .B(n569), .Z(n734) );
  NOR2_X1 U685 ( .A1(G902), .A2(n734), .ZN(n570) );
  NAND2_X1 U686 ( .A1(n591), .A2(n590), .ZN(n571) );
  NOR2_X1 U687 ( .A1(n590), .A2(n591), .ZN(n712) );
  AND2_X2 U688 ( .A1(n581), .A2(n696), .ZN(n588) );
  INV_X1 U689 ( .A(n618), .ZN(n698) );
  AND2_X1 U690 ( .A1(n367), .A2(n349), .ZN(n576) );
  NAND2_X1 U691 ( .A1(KEYINPUT105), .A2(n577), .ZN(n580) );
  INV_X1 U692 ( .A(n577), .ZN(n579) );
  INV_X1 U693 ( .A(KEYINPUT105), .ZN(n578) );
  NOR2_X1 U694 ( .A1(n582), .A2(n609), .ZN(n583) );
  NAND2_X1 U695 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U696 ( .A1(n586), .A2(KEYINPUT44), .ZN(n600) );
  NOR2_X1 U697 ( .A1(n609), .A2(n349), .ZN(n587) );
  NAND2_X1 U698 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U699 ( .A(KEYINPUT103), .B(n589), .ZN(n771) );
  NOR2_X1 U700 ( .A1(n685), .A2(n688), .ZN(n593) );
  AND2_X1 U701 ( .A1(n618), .A2(n357), .ZN(n706) );
  NAND2_X1 U702 ( .A1(n706), .A2(n595), .ZN(n594) );
  XNOR2_X1 U703 ( .A(KEYINPUT31), .B(n594), .ZN(n689) );
  NAND2_X1 U704 ( .A1(n367), .A2(n595), .ZN(n596) );
  NOR2_X1 U705 ( .A1(n689), .A2(n676), .ZN(n597) );
  NOR2_X1 U706 ( .A1(n642), .A2(n597), .ZN(n598) );
  NOR2_X1 U707 ( .A1(n771), .A2(n598), .ZN(n599) );
  NAND2_X1 U708 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U709 ( .A(KEYINPUT87), .B(n601), .ZN(n602) );
  INV_X1 U710 ( .A(n603), .ZN(n711) );
  NAND2_X1 U711 ( .A1(G953), .A2(G900), .ZN(n604) );
  NAND2_X1 U712 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U713 ( .A1(n627), .A2(n701), .ZN(n607) );
  NAND2_X1 U714 ( .A1(n700), .A2(n607), .ZN(n608) );
  NAND2_X1 U715 ( .A1(n696), .A2(n613), .ZN(n610) );
  NOR2_X1 U716 ( .A1(n711), .A2(n610), .ZN(n611) );
  XNOR2_X1 U717 ( .A(n611), .B(KEYINPUT43), .ZN(n612) );
  NOR2_X1 U718 ( .A1(n438), .A2(n612), .ZN(n692) );
  NAND2_X1 U719 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U720 ( .A(KEYINPUT112), .B(KEYINPUT42), .Z(n625) );
  AND2_X1 U721 ( .A1(n618), .A2(n619), .ZN(n620) );
  XOR2_X1 U722 ( .A(KEYINPUT41), .B(KEYINPUT110), .Z(n623) );
  NOR2_X1 U723 ( .A1(n710), .A2(n711), .ZN(n714) );
  NAND2_X1 U724 ( .A1(n638), .A2(n725), .ZN(n624) );
  XNOR2_X1 U725 ( .A(n625), .B(n624), .ZN(n765) );
  NAND2_X1 U726 ( .A1(n438), .A2(n633), .ZN(n635) );
  INV_X1 U727 ( .A(KEYINPUT67), .ZN(n640) );
  NAND2_X1 U728 ( .A1(n640), .A2(n683), .ZN(n641) );
  XNOR2_X1 U729 ( .A(n641), .B(KEYINPUT47), .ZN(n644) );
  NAND2_X1 U730 ( .A1(n642), .A2(n683), .ZN(n643) );
  NAND2_X1 U731 ( .A1(n644), .A2(n643), .ZN(n645) );
  INV_X1 U732 ( .A(n688), .ZN(n648) );
  NOR2_X1 U733 ( .A1(n648), .A2(n647), .ZN(n691) );
  INV_X1 U734 ( .A(KEYINPUT2), .ZN(n651) );
  NOR2_X1 U735 ( .A1(n761), .A2(G952), .ZN(n653) );
  XOR2_X1 U736 ( .A(n653), .B(KEYINPUT93), .Z(n736) );
  INV_X1 U737 ( .A(KEYINPUT120), .ZN(n655) );
  XNOR2_X1 U738 ( .A(n656), .B(n655), .ZN(G54) );
  XNOR2_X1 U739 ( .A(n657), .B(KEYINPUT92), .ZN(n658) );
  INV_X1 U740 ( .A(KEYINPUT59), .ZN(n660) );
  INV_X1 U741 ( .A(KEYINPUT56), .ZN(n666) );
  XOR2_X1 U742 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n662) );
  XOR2_X1 U743 ( .A(KEYINPUT63), .B(KEYINPUT115), .Z(n673) );
  XNOR2_X1 U744 ( .A(n667), .B(KEYINPUT114), .ZN(n669) );
  XOR2_X1 U745 ( .A(KEYINPUT62), .B(KEYINPUT90), .Z(n668) );
  NAND2_X1 U746 ( .A1(n676), .A2(n685), .ZN(n674) );
  XNOR2_X1 U747 ( .A(n674), .B(KEYINPUT116), .ZN(n675) );
  XNOR2_X1 U748 ( .A(G104), .B(n675), .ZN(G6) );
  XOR2_X1 U749 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n678) );
  NAND2_X1 U750 ( .A1(n676), .A2(n688), .ZN(n677) );
  XNOR2_X1 U751 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U752 ( .A(G107), .B(n679), .ZN(G9) );
  XOR2_X1 U753 ( .A(G128), .B(KEYINPUT29), .Z(n681) );
  NAND2_X1 U754 ( .A1(n683), .A2(n688), .ZN(n680) );
  XNOR2_X1 U755 ( .A(n681), .B(n680), .ZN(G30) );
  XOR2_X1 U756 ( .A(G143), .B(n682), .Z(G45) );
  NAND2_X1 U757 ( .A1(n683), .A2(n685), .ZN(n684) );
  XNOR2_X1 U758 ( .A(n684), .B(G146), .ZN(G48) );
  XOR2_X1 U759 ( .A(G113), .B(KEYINPUT117), .Z(n687) );
  NAND2_X1 U760 ( .A1(n689), .A2(n685), .ZN(n686) );
  XNOR2_X1 U761 ( .A(n687), .B(n686), .ZN(G15) );
  NAND2_X1 U762 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U763 ( .A(n690), .B(G116), .ZN(G18) );
  XOR2_X1 U764 ( .A(G134), .B(n691), .Z(G36) );
  XOR2_X1 U765 ( .A(G140), .B(n692), .Z(G42) );
  NAND2_X1 U766 ( .A1(n693), .A2(n739), .ZN(n730) );
  NAND2_X1 U767 ( .A1(G952), .A2(n694), .ZN(n723) );
  NAND2_X1 U768 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U769 ( .A(KEYINPUT50), .B(n697), .ZN(n699) );
  NAND2_X1 U770 ( .A1(n699), .A2(n367), .ZN(n704) );
  NAND2_X1 U771 ( .A1(n701), .A2(n349), .ZN(n702) );
  XNOR2_X1 U772 ( .A(KEYINPUT49), .B(n702), .ZN(n703) );
  NOR2_X1 U773 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U774 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U775 ( .A(n707), .B(KEYINPUT51), .ZN(n708) );
  NAND2_X1 U776 ( .A1(n708), .A2(n725), .ZN(n709) );
  XNOR2_X1 U777 ( .A(n709), .B(KEYINPUT118), .ZN(n720) );
  NAND2_X1 U778 ( .A1(n711), .A2(n710), .ZN(n713) );
  NAND2_X1 U779 ( .A1(n713), .A2(n712), .ZN(n717) );
  NAND2_X1 U780 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U781 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U782 ( .A1(n718), .A2(n724), .ZN(n719) );
  NAND2_X1 U783 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U784 ( .A(KEYINPUT52), .B(n721), .Z(n722) );
  NOR2_X1 U785 ( .A1(n723), .A2(n722), .ZN(n727) );
  AND2_X1 U786 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U787 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U788 ( .A(n728), .B(KEYINPUT119), .ZN(n729) );
  NOR2_X1 U789 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U790 ( .A(KEYINPUT53), .B(n731), .ZN(G75) );
  XOR2_X1 U791 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n733) );
  NOR2_X1 U792 ( .A1(n736), .A2(n735), .ZN(G63) );
  NOR2_X1 U793 ( .A1(G898), .A2(n739), .ZN(n743) );
  XOR2_X1 U794 ( .A(n741), .B(n740), .Z(n742) );
  NOR2_X1 U795 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U796 ( .A(KEYINPUT124), .B(n744), .Z(n751) );
  NAND2_X1 U797 ( .A1(G953), .A2(G224), .ZN(n745) );
  XNOR2_X1 U798 ( .A(KEYINPUT61), .B(n745), .ZN(n746) );
  NAND2_X1 U799 ( .A1(n746), .A2(G898), .ZN(n749) );
  NAND2_X1 U800 ( .A1(n747), .A2(n761), .ZN(n748) );
  NAND2_X1 U801 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U802 ( .A(n751), .B(n750), .Z(G69) );
  XOR2_X1 U803 ( .A(KEYINPUT125), .B(n752), .Z(n753) );
  XOR2_X1 U804 ( .A(n755), .B(n754), .Z(n759) );
  XOR2_X1 U805 ( .A(G227), .B(n759), .Z(n756) );
  NAND2_X1 U806 ( .A1(n756), .A2(G900), .ZN(n757) );
  NAND2_X1 U807 ( .A1(n757), .A2(G953), .ZN(n764) );
  XNOR2_X1 U808 ( .A(n759), .B(n758), .ZN(n760) );
  XNOR2_X1 U809 ( .A(n760), .B(KEYINPUT126), .ZN(n762) );
  NAND2_X1 U810 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U811 ( .A1(n764), .A2(n763), .ZN(G72) );
  XOR2_X1 U812 ( .A(n765), .B(G137), .Z(G39) );
  XNOR2_X1 U813 ( .A(n766), .B(G125), .ZN(n767) );
  XNOR2_X1 U814 ( .A(n767), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U815 ( .A(G122), .B(n768), .Z(G24) );
  BUF_X1 U816 ( .A(n769), .Z(n770) );
  XOR2_X1 U817 ( .A(G110), .B(n770), .Z(G12) );
  XOR2_X1 U818 ( .A(G101), .B(n771), .Z(G3) );
  XOR2_X1 U819 ( .A(n772), .B(G119), .Z(G21) );
  XOR2_X1 U820 ( .A(n773), .B(G131), .Z(G33) );
endmodule

