//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n527, new_n528, new_n529, new_n531, new_n532, new_n533, new_n534,
    new_n536, new_n538, new_n539, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n584, new_n585, new_n588, new_n590, new_n591,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT66), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT67), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT68), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT69), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n453), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n463), .B(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  OR2_X1    g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n470), .A2(G137), .B1(G101), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n467), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n470), .A2(G136), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n461), .A2(G2105), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT71), .ZN(new_n482));
  AOI211_X1 g057(.A(new_n477), .B(new_n480), .C1(new_n482), .C2(G124), .ZN(G162));
  AND2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  OAI211_X1 g060(.A(G138), .B(new_n471), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT72), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n461), .A2(G138), .A3(new_n471), .A4(new_n488), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n471), .B1(new_n468), .B2(new_n469), .ZN(new_n493));
  OR2_X1    g068(.A1(new_n471), .A2(G114), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n493), .A2(G126), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(KEYINPUT73), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .A3(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n508), .A2(new_n514), .ZN(G166));
  NAND3_X1  g090(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  INV_X1    g093(.A(G89), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n516), .B(new_n518), .C1(new_n510), .C2(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n509), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT74), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT74), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n512), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n520), .B1(new_n525), .B2(G51), .ZN(G168));
  AOI22_X1  g101(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n527), .A2(new_n507), .B1(new_n528), .B2(new_n510), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n529), .B1(G52), .B2(new_n525), .ZN(G171));
  AOI22_X1  g105(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT75), .B(G81), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n531), .A2(new_n507), .B1(new_n510), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n533), .B1(G43), .B2(new_n525), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G860), .ZN(G153));
  AND3_X1   g110(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G36), .ZN(G176));
  NAND2_X1  g112(.A1(G1), .A2(G3), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT8), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n536), .A2(new_n539), .ZN(G188));
  NAND2_X1  g115(.A1(G78), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(new_n505), .ZN(new_n542));
  INV_X1    g117(.A(G65), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n505), .A2(new_n509), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n544), .A2(G651), .B1(new_n545), .B2(G91), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT9), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n521), .A2(new_n547), .A3(G53), .ZN(new_n548));
  INV_X1    g123(.A(G53), .ZN(new_n549));
  OAI21_X1  g124(.A(KEYINPUT9), .B1(new_n512), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n546), .A2(new_n551), .ZN(G299));
  INV_X1    g127(.A(G171), .ZN(G301));
  INV_X1    g128(.A(G168), .ZN(G286));
  INV_X1    g129(.A(G166), .ZN(G303));
  OAI21_X1  g130(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n505), .A2(G87), .A3(new_n509), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n509), .A2(G49), .A3(G543), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(G288));
  AOI22_X1  g134(.A1(new_n545), .A2(G86), .B1(new_n521), .B2(G48), .ZN(new_n560));
  AND2_X1   g135(.A1(new_n505), .A2(G61), .ZN(new_n561));
  NAND2_X1  g136(.A1(G73), .A2(G543), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT76), .Z(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n560), .A2(new_n564), .ZN(G305));
  XOR2_X1   g140(.A(KEYINPUT77), .B(G47), .Z(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(new_n522), .B2(new_n524), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n568));
  XOR2_X1   g143(.A(KEYINPUT78), .B(G85), .Z(new_n569));
  OAI22_X1  g144(.A1(new_n568), .A2(new_n507), .B1(new_n510), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G290));
  NAND2_X1  g147(.A1(G301), .A2(G868), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n545), .A2(G92), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT10), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n574), .B(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n505), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(new_n507), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n525), .B2(G54), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n573), .B1(new_n581), .B2(G868), .ZN(G284));
  OAI21_X1  g157(.A(new_n573), .B1(new_n581), .B2(G868), .ZN(G321));
  INV_X1    g158(.A(G868), .ZN(new_n584));
  NAND2_X1  g159(.A1(G299), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n585), .B1(new_n584), .B2(G168), .ZN(G297));
  XNOR2_X1  g161(.A(G297), .B(KEYINPUT79), .ZN(G280));
  INV_X1    g162(.A(G559), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n581), .B1(new_n588), .B2(G860), .ZN(G148));
  NAND2_X1  g164(.A1(new_n581), .A2(new_n588), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G868), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n591), .B1(G868), .B2(new_n534), .ZN(G323));
  XNOR2_X1  g167(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g168(.A1(new_n470), .A2(G2104), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT12), .ZN(new_n595));
  XOR2_X1   g170(.A(new_n595), .B(KEYINPUT13), .Z(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(G2100), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(G2100), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n470), .A2(G135), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n471), .A2(G111), .ZN(new_n600));
  OAI21_X1  g175(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n493), .B(KEYINPUT71), .ZN(new_n602));
  INV_X1    g177(.A(G123), .ZN(new_n603));
  OAI221_X1 g178(.A(new_n599), .B1(new_n600), .B2(new_n601), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(G2096), .Z(new_n605));
  NAND3_X1  g180(.A1(new_n597), .A2(new_n598), .A3(new_n605), .ZN(G156));
  INV_X1    g181(.A(KEYINPUT14), .ZN(new_n607));
  XNOR2_X1  g182(.A(G2427), .B(G2438), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(G2430), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT15), .B(G2435), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(new_n610), .B2(new_n609), .ZN(new_n612));
  XNOR2_X1  g187(.A(G2451), .B(G2454), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT16), .ZN(new_n614));
  XNOR2_X1  g189(.A(G1341), .B(G1348), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n612), .B(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(G2443), .B(G2446), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(G14), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(new_n620), .B2(new_n618), .ZN(G401));
  XOR2_X1   g197(.A(G2067), .B(G2678), .Z(new_n623));
  XNOR2_X1  g198(.A(G2084), .B(G2090), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT80), .B(KEYINPUT17), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT18), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2072), .B(G2078), .Z(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(new_n625), .B2(KEYINPUT18), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n630), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT81), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2096), .B(G2100), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(G227));
  XNOR2_X1  g211(.A(G1971), .B(G1976), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT19), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G1956), .B(G2474), .Z(new_n640));
  XOR2_X1   g215(.A(G1961), .B(G1966), .Z(new_n641));
  NOR2_X1   g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g217(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n640), .A2(new_n641), .ZN(new_n644));
  NOR3_X1   g219(.A1(new_n639), .A2(new_n644), .A3(new_n642), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n639), .A2(new_n644), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n647));
  AOI211_X1 g222(.A(new_n643), .B(new_n645), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n646), .B2(new_n647), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT83), .ZN(new_n650));
  XOR2_X1   g225(.A(G1981), .B(G1986), .Z(new_n651));
  XNOR2_X1  g226(.A(G1991), .B(G1996), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n650), .B(new_n655), .ZN(G229));
  INV_X1    g231(.A(G29), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(G25), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n470), .A2(G131), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n471), .A2(G107), .ZN(new_n660));
  OAI21_X1  g235(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n661));
  INV_X1    g236(.A(G119), .ZN(new_n662));
  OAI221_X1 g237(.A(new_n659), .B1(new_n660), .B2(new_n661), .C1(new_n602), .C2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT84), .Z(new_n664));
  OAI21_X1  g239(.A(new_n658), .B1(new_n664), .B2(new_n657), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT35), .B(G1991), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT85), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n665), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(G16), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(G24), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(new_n571), .B2(new_n670), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT86), .B(G1986), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(G16), .A2(G23), .ZN(new_n675));
  NAND2_X1  g250(.A1(G288), .A2(KEYINPUT87), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT87), .ZN(new_n677));
  NAND4_X1  g252(.A1(new_n556), .A2(new_n557), .A3(new_n677), .A4(new_n558), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n675), .B1(new_n679), .B2(G16), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT33), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n670), .A2(G22), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(G166), .B2(new_n670), .ZN(new_n684));
  INV_X1    g259(.A(G1971), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  MUX2_X1   g261(.A(G6), .B(G305), .S(G16), .Z(new_n687));
  XOR2_X1   g262(.A(KEYINPUT32), .B(G1981), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n682), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n669), .B(new_n674), .C1(new_n690), .C2(KEYINPUT34), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT88), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(KEYINPUT36), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n690), .A2(KEYINPUT34), .ZN(new_n695));
  OR3_X1    g270(.A1(new_n691), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n694), .B1(new_n691), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n657), .A2(G33), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT25), .Z(new_n701));
  NAND2_X1  g276(.A1(new_n470), .A2(G139), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT93), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n703), .B2(new_n702), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT94), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n461), .A2(G127), .ZN(new_n708));
  AND2_X1   g283(.A1(G115), .A2(G2104), .ZN(new_n709));
  OAI21_X1  g284(.A(G2105), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n699), .B1(new_n711), .B2(new_n657), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G2072), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT95), .ZN(new_n714));
  NOR2_X1   g289(.A1(G29), .A2(G35), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G162), .B2(G29), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n718), .A2(G2090), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT99), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n670), .A2(G5), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G171), .B2(new_n670), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(G1961), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT31), .B(G11), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT30), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n726), .A2(G28), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n657), .B1(new_n726), .B2(G28), .ZN(new_n728));
  OAI221_X1 g303(.A(new_n725), .B1(new_n727), .B2(new_n728), .C1(new_n604), .C2(new_n657), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT24), .ZN(new_n730));
  INV_X1    g305(.A(G34), .ZN(new_n731));
  AOI21_X1  g306(.A(G29), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n730), .B2(new_n731), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G160), .B2(new_n657), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n729), .B1(G2084), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n723), .A2(G1961), .ZN(new_n736));
  NOR2_X1   g311(.A1(G168), .A2(new_n670), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n670), .B2(G21), .ZN(new_n738));
  INV_X1    g313(.A(G1966), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n735), .A2(new_n736), .A3(new_n740), .ZN(new_n741));
  NOR3_X1   g316(.A1(new_n721), .A2(new_n724), .A3(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n712), .A2(G2072), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n719), .A2(new_n720), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n734), .A2(G2084), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT96), .Z(new_n747));
  AND2_X1   g322(.A1(new_n657), .A2(G32), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n482), .A2(G129), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n472), .A2(G105), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT26), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n750), .B(new_n752), .C1(G141), .C2(new_n470), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n748), .B1(new_n754), .B2(G29), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT27), .B(G1996), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G164), .A2(new_n657), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G27), .B2(new_n657), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT97), .B(G2078), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n747), .A2(new_n757), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n670), .A2(G20), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT23), .Z(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G299), .B2(G16), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1956), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n718), .B2(G2090), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n759), .A2(new_n760), .ZN(new_n768));
  OAI22_X1  g343(.A1(new_n738), .A2(new_n739), .B1(new_n755), .B2(new_n756), .ZN(new_n769));
  NOR4_X1   g344(.A1(new_n762), .A2(new_n767), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n714), .A2(new_n742), .A3(new_n745), .A4(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G4), .A2(G16), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n581), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT89), .B(G1348), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n657), .A2(G26), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT28), .ZN(new_n777));
  OAI21_X1  g352(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n778));
  INV_X1    g353(.A(G116), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(G2105), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G140), .B2(new_n470), .ZN(new_n781));
  INV_X1    g356(.A(G128), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n602), .B2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n777), .B1(new_n785), .B2(new_n657), .ZN(new_n786));
  INV_X1    g361(.A(G2067), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n670), .A2(G19), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n534), .B2(new_n670), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT90), .B(G1341), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n775), .A2(new_n788), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT92), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n771), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n698), .A2(new_n795), .ZN(G150));
  INV_X1    g371(.A(G150), .ZN(G311));
  XNOR2_X1  g372(.A(KEYINPUT100), .B(G55), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n525), .A2(new_n798), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(new_n507), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n545), .A2(G93), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n799), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(G860), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT37), .Z(new_n805));
  NAND2_X1  g380(.A1(new_n581), .A2(G559), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT101), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT38), .ZN(new_n808));
  AND3_X1   g383(.A1(new_n799), .A2(new_n801), .A3(new_n802), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(new_n534), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n808), .B(new_n810), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n811), .A2(KEYINPUT39), .ZN(new_n812));
  INV_X1    g387(.A(G860), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n811), .B2(KEYINPUT39), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n805), .B1(new_n812), .B2(new_n814), .ZN(G145));
  XNOR2_X1  g390(.A(new_n604), .B(new_n474), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G162), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n783), .B(KEYINPUT91), .ZN(new_n818));
  AND3_X1   g393(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT102), .ZN(new_n819));
  AOI21_X1  g394(.A(KEYINPUT102), .B1(new_n490), .B2(new_n491), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n497), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n818), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(new_n711), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n785), .B(new_n821), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n707), .A2(new_n710), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(new_n754), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n823), .A2(new_n826), .A3(new_n749), .A4(new_n753), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n470), .A2(G142), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n471), .A2(G118), .ZN(new_n832));
  OAI21_X1  g407(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n482), .B2(G130), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(new_n595), .Z(new_n836));
  XOR2_X1   g411(.A(new_n664), .B(new_n836), .Z(new_n837));
  AOI21_X1  g412(.A(new_n817), .B1(new_n830), .B2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n837), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n828), .A2(new_n829), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(G37), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT103), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n830), .B1(new_n842), .B2(new_n839), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n828), .A2(KEYINPUT103), .A3(new_n829), .A4(new_n837), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n843), .A2(new_n844), .A3(new_n817), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n841), .A2(KEYINPUT40), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(KEYINPUT40), .B1(new_n841), .B2(new_n845), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(G395));
  INV_X1    g423(.A(KEYINPUT106), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n580), .A2(G299), .ZN(new_n850));
  INV_X1    g425(.A(G299), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n851), .A2(new_n576), .A3(new_n579), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT41), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n850), .A2(KEYINPUT41), .A3(new_n852), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n580), .A2(G559), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n810), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n803), .B(new_n534), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n859), .A2(new_n590), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n855), .B(new_n856), .C1(new_n858), .C2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT105), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n855), .A2(new_n856), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT105), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n863), .B(new_n864), .C1(new_n860), .C2(new_n858), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n810), .A2(new_n857), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n859), .A2(new_n590), .ZN(new_n867));
  INV_X1    g442(.A(new_n853), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT104), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n862), .B(new_n865), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n679), .B(G305), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(G303), .A2(new_n571), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(G303), .A2(new_n571), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT42), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT42), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n880), .A2(new_n884), .A3(new_n881), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n873), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n869), .B(new_n870), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n889), .A2(new_n865), .A3(new_n862), .A4(new_n886), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(G868), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n809), .A2(G868), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n849), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n584), .B1(new_n888), .B2(new_n890), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n896), .A2(KEYINPUT106), .A3(new_n893), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n895), .A2(new_n897), .ZN(G295));
  NAND2_X1  g473(.A1(new_n892), .A2(new_n894), .ZN(G331));
  XNOR2_X1  g474(.A(G171), .B(G168), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n810), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n900), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n859), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT108), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n901), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n902), .A2(new_n859), .A3(KEYINPUT108), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(new_n863), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT109), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n901), .A2(new_n903), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n810), .A2(KEYINPUT109), .A3(new_n900), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n882), .B(new_n907), .C1(new_n911), .C2(new_n853), .ZN(new_n912));
  INV_X1    g487(.A(G37), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n915));
  INV_X1    g490(.A(new_n882), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n909), .A2(new_n863), .A3(new_n910), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n853), .B1(new_n905), .B2(new_n906), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n914), .A2(KEYINPUT110), .A3(new_n915), .A4(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n905), .A2(new_n863), .A3(new_n906), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n853), .B1(new_n909), .B2(new_n910), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n916), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(new_n912), .A3(new_n913), .ZN(new_n925));
  INV_X1    g500(.A(new_n915), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n919), .A2(new_n912), .A3(new_n913), .A4(new_n915), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n920), .B(new_n921), .C1(new_n927), .C2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n919), .A2(new_n912), .A3(new_n913), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT111), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n924), .A2(new_n912), .A3(new_n913), .A4(new_n915), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n936), .A2(KEYINPUT44), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n932), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n931), .A2(new_n939), .ZN(G397));
  XNOR2_X1  g515(.A(new_n664), .B(new_n668), .ZN(new_n941));
  XOR2_X1   g516(.A(new_n754), .B(G1996), .Z(new_n942));
  NAND2_X1  g517(.A1(new_n818), .A2(G2067), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n785), .A2(new_n787), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n571), .B(G1986), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n497), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT102), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n488), .B1(new_n470), .B2(G138), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n486), .A2(new_n489), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT102), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n949), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT112), .B1(new_n955), .B2(G1384), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT112), .ZN(new_n958));
  INV_X1    g533(.A(G1384), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n821), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n956), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n467), .A2(G40), .A3(new_n473), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n948), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT62), .ZN(new_n965));
  INV_X1    g540(.A(G2084), .ZN(new_n966));
  INV_X1    g541(.A(new_n962), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n968));
  AOI21_X1  g543(.A(G1384), .B1(new_n492), .B2(new_n497), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT114), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n953), .A2(new_n954), .ZN(new_n973));
  AOI21_X1  g548(.A(G1384), .B1(new_n973), .B2(new_n497), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n972), .B1(new_n974), .B2(new_n968), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n821), .A2(new_n972), .A3(new_n968), .A4(new_n959), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n966), .B(new_n971), .C1(new_n975), .C2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n821), .A2(new_n959), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n957), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n962), .B1(KEYINPUT45), .B2(new_n969), .ZN(new_n981));
  AOI21_X1  g556(.A(G1966), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n978), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(KEYINPUT115), .B(G8), .ZN(new_n985));
  NOR2_X1   g560(.A1(G168), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n821), .A2(new_n968), .A3(new_n959), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT114), .ZN(new_n990));
  AOI211_X1 g565(.A(G2084), .B(new_n970), .C1(new_n990), .C2(new_n976), .ZN(new_n991));
  OAI21_X1  g566(.A(G8), .B1(new_n991), .B2(new_n982), .ZN(new_n992));
  INV_X1    g567(.A(new_n986), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n988), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n988), .ZN(new_n995));
  INV_X1    g570(.A(new_n985), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n995), .B1(new_n984), .B2(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n965), .B(new_n987), .C1(new_n994), .C2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(G2078), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n980), .A2(new_n981), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n971), .B1(new_n975), .B2(new_n977), .ZN(new_n1002));
  INV_X1    g577(.A(G1961), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT45), .B1(new_n498), .B2(new_n959), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n962), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G2078), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n821), .A2(KEYINPUT45), .A3(new_n959), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT113), .B1(new_n969), .B2(KEYINPUT45), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1011), .A2(new_n999), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(G301), .B1(new_n1004), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(G303), .A2(G8), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT55), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n968), .B1(new_n821), .B2(new_n959), .ZN(new_n1017));
  INV_X1    g592(.A(new_n969), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n967), .B1(new_n1018), .B2(KEYINPUT50), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1017), .A2(new_n1019), .A3(G2090), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1020), .B1(new_n685), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1016), .B1(new_n1022), .B2(new_n985), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1016), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(new_n685), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  AOI211_X1 g601(.A(G2090), .B(new_n970), .C1(new_n990), .C2(new_n976), .ZN(new_n1027));
  OAI211_X1 g602(.A(G8), .B(new_n1024), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(G305), .A2(KEYINPUT49), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n564), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G1981), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT49), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1033), .B1(new_n560), .B2(new_n564), .ZN(new_n1034));
  OR3_X1    g609(.A1(new_n1029), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n985), .B1(new_n974), .B2(new_n967), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1032), .B1(new_n1029), .B2(new_n1034), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n676), .A2(KEYINPUT116), .A3(G1976), .A4(new_n678), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n676), .A2(G1976), .A3(new_n678), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT117), .B(G1976), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT52), .B1(G288), .B2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1036), .A2(new_n1039), .A3(new_n1042), .A4(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n967), .A2(new_n821), .A3(new_n959), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1042), .A2(new_n1046), .A3(new_n996), .A4(new_n1039), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT52), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1038), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  AND4_X1   g625(.A1(new_n1014), .A2(new_n1023), .A3(new_n1028), .A4(new_n1050), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n998), .A2(new_n1051), .A3(KEYINPUT126), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT126), .B1(new_n998), .B2(new_n1051), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n986), .B1(new_n984), .B2(G8), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n970), .B1(new_n990), .B2(new_n976), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n982), .B1(new_n1055), .B2(new_n966), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1056), .A2(new_n985), .ZN(new_n1057));
  OAI22_X1  g632(.A1(new_n1054), .A2(new_n988), .B1(new_n1057), .B2(new_n995), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n965), .B1(new_n1058), .B2(new_n987), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1052), .A2(new_n1053), .A3(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(G288), .A2(G1976), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1038), .A2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(G305), .A2(G1981), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1036), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1064), .B1(new_n1028), .B2(new_n1049), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT63), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1023), .A2(new_n1028), .A3(new_n1050), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1057), .A2(G168), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G8), .ZN(new_n1070));
  INV_X1    g645(.A(G2090), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1055), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1070), .B1(new_n1072), .B2(new_n1025), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1049), .B1(new_n1073), .B2(new_n1024), .ZN(new_n1074));
  NOR4_X1   g649(.A1(new_n1056), .A2(new_n1066), .A3(G286), .A4(new_n985), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1074), .B(new_n1075), .C1(new_n1024), .C2(new_n1073), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1065), .B1(new_n1069), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT57), .B1(new_n551), .B2(KEYINPUT119), .ZN(new_n1078));
  XNOR2_X1  g653(.A(G299), .B(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1956), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT56), .B(G2072), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1079), .B1(new_n1084), .B2(KEYINPUT120), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(KEYINPUT120), .B2(new_n1084), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1046), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n787), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n1055), .B2(G1348), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1079), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(new_n581), .A3(new_n1090), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1086), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT60), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1093), .B1(new_n581), .B2(KEYINPUT122), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1094), .B(new_n1088), .C1(new_n1055), .C2(G1348), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(new_n1096), .A3(new_n580), .ZN(new_n1097));
  INV_X1    g672(.A(G1348), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1002), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n580), .A2(new_n1096), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1099), .A2(new_n1088), .A3(new_n1094), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1097), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1079), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT61), .B1(new_n1084), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT61), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT121), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1090), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1079), .B1(new_n1083), .B2(new_n1081), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1090), .B(new_n1107), .C1(new_n1110), .C2(KEYINPUT61), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT58), .B(G1341), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n1021), .A2(G1996), .B1(new_n1087), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n534), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(KEYINPUT59), .A3(new_n534), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1109), .A2(new_n1111), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1092), .B1(new_n1103), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1067), .B1(new_n1058), .B2(new_n987), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1000), .A2(G40), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n466), .A2(KEYINPUT123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(G2105), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n466), .A2(KEYINPUT123), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n473), .B(new_n1123), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1127), .B1(new_n974), .B2(KEYINPUT45), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n961), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(new_n1055), .B2(G1961), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1130), .A2(G171), .A3(new_n1012), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1122), .B1(new_n1014), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g709(.A(KEYINPUT124), .B(new_n1122), .C1(new_n1014), .C2(new_n1131), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n980), .A2(new_n981), .A3(new_n1000), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1055), .B2(G1961), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1137), .A2(new_n1012), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1122), .B1(new_n1138), .B2(G301), .ZN(new_n1139));
  OAI21_X1  g714(.A(G171), .B1(new_n1130), .B2(new_n1012), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT125), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT125), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1142), .B(G171), .C1(new_n1130), .C2(new_n1012), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1139), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1134), .A2(new_n1135), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1077), .B1(new_n1121), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n964), .B1(new_n1060), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n943), .A2(new_n944), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n963), .B1(new_n1148), .B2(new_n754), .ZN(new_n1149));
  INV_X1    g724(.A(new_n963), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1150), .A2(G1996), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1149), .B1(new_n1151), .B2(KEYINPUT46), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1152), .B1(KEYINPUT46), .B2(new_n1151), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT47), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n664), .A2(new_n668), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n944), .B1(new_n945), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n963), .ZN(new_n1157));
  OR3_X1    g732(.A1(new_n1150), .A2(G1986), .A3(G290), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT48), .ZN(new_n1159));
  OAI22_X1  g734(.A1(new_n946), .A2(new_n1150), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1157), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1154), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1147), .A2(new_n1163), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g739(.A1(G227), .A2(new_n459), .ZN(new_n1166));
  OR2_X1    g740(.A1(new_n1166), .A2(KEYINPUT127), .ZN(new_n1167));
  NAND2_X1  g741(.A1(new_n1166), .A2(KEYINPUT127), .ZN(new_n1168));
  NOR2_X1   g742(.A1(G229), .A2(G401), .ZN(new_n1169));
  NAND3_X1  g743(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g744(.A(new_n1170), .B1(new_n841), .B2(new_n845), .ZN(new_n1171));
  NAND2_X1  g745(.A1(new_n925), .A2(new_n926), .ZN(new_n1172));
  NAND3_X1  g746(.A1(new_n1172), .A2(new_n929), .A3(new_n928), .ZN(new_n1173));
  AND3_X1   g747(.A1(new_n1171), .A2(new_n1173), .A3(new_n920), .ZN(G308));
  NAND3_X1  g748(.A1(new_n1171), .A2(new_n1173), .A3(new_n920), .ZN(G225));
endmodule


