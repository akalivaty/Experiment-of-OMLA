//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  AND3_X1   g001(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n188));
  AOI21_X1  g002(.A(G143), .B1(new_n187), .B2(G214), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT18), .ZN(new_n191));
  INV_X1    g005(.A(G131), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n190), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  OAI211_X1 g007(.A(KEYINPUT18), .B(G131), .C1(new_n188), .C2(new_n189), .ZN(new_n194));
  XNOR2_X1  g008(.A(G125), .B(G140), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n195), .B(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n193), .A2(new_n194), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G125), .ZN(new_n200));
  NOR3_X1   g014(.A1(new_n200), .A2(KEYINPUT16), .A3(G140), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n201), .B1(new_n195), .B2(KEYINPUT16), .ZN(new_n202));
  XNOR2_X1  g016(.A(new_n202), .B(G146), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT85), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G131), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n190), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n205), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n207), .B(KEYINPUT85), .C1(new_n188), .C2(new_n189), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n203), .B1(new_n209), .B2(KEYINPUT17), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT17), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n190), .A2(new_n205), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n206), .A2(new_n211), .A3(new_n208), .A4(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n199), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G113), .B(G122), .ZN(new_n215));
  INV_X1    g029(.A(G104), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n215), .B(new_n216), .ZN(new_n217));
  XOR2_X1   g031(.A(new_n217), .B(KEYINPUT86), .Z(new_n218));
  INV_X1    g032(.A(new_n217), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n206), .A2(new_n208), .A3(new_n212), .ZN(new_n220));
  INV_X1    g034(.A(new_n201), .ZN(new_n221));
  INV_X1    g035(.A(G140), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G125), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n200), .A2(G140), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT16), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n221), .A2(new_n225), .A3(G146), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n195), .B(KEYINPUT19), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n226), .B1(new_n227), .B2(new_n196), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n220), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n198), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n214), .A2(new_n218), .B1(new_n219), .B2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(G475), .A2(G902), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT20), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n209), .A2(KEYINPUT17), .ZN(new_n235));
  INV_X1    g049(.A(new_n203), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n213), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n198), .A3(new_n218), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n230), .A2(new_n219), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT20), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(new_n241), .A3(new_n232), .ZN(new_n242));
  INV_X1    g056(.A(G902), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n237), .A2(new_n198), .A3(new_n218), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n217), .B1(new_n237), .B2(new_n198), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n234), .A2(new_n242), .B1(new_n246), .B2(G475), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT13), .ZN(new_n248));
  INV_X1    g062(.A(G128), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(G143), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(G143), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G128), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(new_n248), .ZN(new_n255));
  OAI21_X1  g069(.A(G134), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G134), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n254), .A2(new_n251), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G122), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G116), .ZN(new_n260));
  INV_X1    g074(.A(G116), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G122), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G107), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n263), .A2(G107), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n256), .B(new_n258), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT9), .B(G234), .ZN(new_n269));
  INV_X1    g083(.A(G217), .ZN(new_n270));
  NOR3_X1   g084(.A1(new_n269), .A2(new_n270), .A3(G953), .ZN(new_n271));
  INV_X1    g085(.A(new_n258), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n257), .B1(new_n254), .B2(new_n251), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT87), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n254), .A2(new_n251), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G134), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT87), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n277), .A3(new_n258), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT14), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n260), .A2(new_n262), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n261), .A2(KEYINPUT14), .A3(G122), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n280), .A2(KEYINPUT88), .A3(G107), .A4(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n274), .A2(new_n278), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(G107), .A3(new_n281), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT88), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n267), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n268), .B(new_n271), .C1(new_n283), .C2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n267), .B1(new_n284), .B2(new_n285), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n291), .A2(new_n278), .A3(new_n282), .A4(new_n274), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n271), .B1(new_n292), .B2(new_n268), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n243), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G478), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(KEYINPUT15), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n294), .B(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G952), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n298), .A2(G953), .ZN(new_n299));
  NAND2_X1  g113(.A1(G234), .A2(G237), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT21), .B(G898), .Z(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(G902), .A3(G953), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  XOR2_X1   g118(.A(new_n304), .B(KEYINPUT89), .Z(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n297), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n247), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT90), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n247), .A2(KEYINPUT90), .A3(new_n307), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(G221), .B1(new_n269), .B2(G902), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G469), .ZN(new_n315));
  XNOR2_X1  g129(.A(G110), .B(G140), .ZN(new_n316));
  INV_X1    g130(.A(G953), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G227), .ZN(new_n318));
  XOR2_X1   g132(.A(new_n316), .B(new_n318), .Z(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(KEYINPUT3), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n216), .A2(G107), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(KEYINPUT3), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n326), .A2(new_n265), .A3(KEYINPUT74), .A4(G104), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n216), .A2(G107), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(G101), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n265), .A2(G104), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(new_n322), .B2(new_n323), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT75), .B(G101), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n326), .A2(KEYINPUT74), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n326), .A2(KEYINPUT74), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n265), .A2(G104), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n332), .A2(new_n333), .A3(new_n337), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n330), .A2(KEYINPUT4), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n196), .A2(G143), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n253), .A2(G146), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT0), .A4(G128), .ZN(new_n342));
  XNOR2_X1  g156(.A(G143), .B(G146), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT0), .B(G128), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n347), .B(G101), .C1(new_n325), .C2(new_n329), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT10), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n340), .B(new_n341), .C1(KEYINPUT1), .C2(new_n249), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT1), .B1(new_n253), .B2(G146), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n253), .A2(G146), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n196), .A2(G143), .ZN(new_n354));
  OAI211_X1 g168(.A(G128), .B(new_n352), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G101), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n336), .B2(new_n328), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n338), .A2(new_n351), .A3(new_n355), .A4(new_n358), .ZN(new_n359));
  OAI22_X1  g173(.A1(new_n339), .A2(new_n349), .B1(new_n350), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n350), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT76), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT76), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n359), .A2(new_n363), .A3(new_n350), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n360), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G137), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT64), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT64), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G137), .ZN(new_n369));
  AND2_X1   g183(.A1(KEYINPUT11), .A2(G134), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(KEYINPUT11), .A2(G134), .ZN(new_n372));
  NOR2_X1   g186(.A1(KEYINPUT11), .A2(G134), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n372), .B1(new_n373), .B2(G137), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G131), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT66), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n371), .A2(new_n374), .A3(new_n205), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT66), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n375), .A2(new_n379), .A3(G131), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT78), .B1(new_n365), .B2(new_n382), .ZN(new_n383));
  XOR2_X1   g197(.A(KEYINPUT75), .B(G101), .Z(new_n384));
  NOR3_X1   g198(.A1(new_n325), .A2(new_n329), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n355), .A2(new_n351), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n385), .A2(new_n386), .A3(new_n357), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n356), .B1(new_n332), .B2(new_n337), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n345), .B1(new_n388), .B2(new_n347), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n330), .A2(KEYINPUT4), .A3(new_n338), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n387), .A2(KEYINPUT10), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n363), .B1(new_n359), .B2(new_n350), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n359), .A2(new_n363), .A3(new_n350), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT78), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(new_n381), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n383), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n391), .B(new_n382), .C1(new_n392), .C2(new_n393), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n320), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT12), .B1(new_n381), .B2(KEYINPUT77), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n338), .A2(new_n358), .B1(new_n351), .B2(new_n355), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n381), .B1(new_n387), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT79), .ZN(new_n404));
  OAI221_X1 g218(.A(new_n381), .B1(KEYINPUT77), .B2(KEYINPUT12), .C1(new_n387), .C2(new_n401), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n398), .A2(new_n320), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n404), .B1(new_n403), .B2(new_n405), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n315), .B(new_n243), .C1(new_n399), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n403), .A2(new_n405), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n320), .B1(new_n411), .B2(new_n398), .ZN(new_n412));
  INV_X1    g226(.A(new_n407), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n412), .B1(new_n397), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(G469), .B1(new_n414), .B2(G902), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n314), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n312), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(G210), .B1(G237), .B2(G902), .ZN(new_n418));
  INV_X1    g232(.A(G119), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G116), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n261), .A2(G119), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT2), .B(G113), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n423), .ZN(new_n425));
  XNOR2_X1  g239(.A(G116), .B(G119), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n388), .A2(new_n347), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n325), .A2(new_n329), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n357), .B1(new_n429), .B2(new_n333), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n422), .A2(new_n423), .ZN(new_n431));
  INV_X1    g245(.A(G113), .ZN(new_n432));
  XOR2_X1   g246(.A(KEYINPUT80), .B(KEYINPUT5), .Z(new_n433));
  INV_X1    g247(.A(new_n420), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n426), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n431), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n428), .A2(new_n390), .B1(new_n430), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G122), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT81), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n442), .B1(new_n439), .B2(new_n440), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n427), .A2(new_n424), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n348), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n338), .A2(new_n358), .ZN(new_n446));
  INV_X1    g260(.A(new_n437), .ZN(new_n447));
  OAI21_X1  g261(.A(G113), .B1(new_n436), .B2(new_n420), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n427), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI22_X1  g263(.A1(new_n339), .A2(new_n445), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT81), .ZN(new_n451));
  INV_X1    g265(.A(new_n440), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n441), .A2(new_n443), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n345), .A2(G125), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n355), .A2(new_n351), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n455), .B1(new_n456), .B2(G125), .ZN(new_n457));
  INV_X1    g271(.A(G224), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(G953), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n457), .B(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n439), .A2(new_n440), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT82), .B1(new_n461), .B2(new_n442), .ZN(new_n462));
  AND4_X1   g276(.A1(KEYINPUT82), .A2(new_n450), .A3(new_n442), .A4(new_n452), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n454), .B(new_n460), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT7), .B1(new_n458), .B2(G953), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n457), .B(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n448), .B1(KEYINPUT5), .B2(new_n426), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n430), .B1(new_n431), .B2(new_n467), .ZN(new_n468));
  XOR2_X1   g282(.A(new_n440), .B(KEYINPUT8), .Z(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(new_n438), .B2(new_n446), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n466), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n439), .A2(new_n440), .ZN(new_n472));
  AOI21_X1  g286(.A(G902), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n418), .B1(new_n464), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(KEYINPUT83), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT83), .ZN(new_n476));
  AOI211_X1 g290(.A(new_n476), .B(new_n418), .C1(new_n464), .C2(new_n473), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n464), .A2(new_n473), .A3(new_n418), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT84), .ZN(new_n481));
  OAI21_X1  g295(.A(G214), .B1(G237), .B2(G902), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n464), .A2(new_n473), .ZN(new_n485));
  INV_X1    g299(.A(new_n418), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n476), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n474), .A2(KEYINPUT83), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(new_n478), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT84), .B1(new_n490), .B2(new_n482), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n417), .B1(new_n484), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n380), .A2(new_n378), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n192), .B1(new_n371), .B2(new_n374), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n494), .A2(new_n379), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n346), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n444), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n367), .A2(new_n369), .A3(new_n257), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n498), .B(G131), .C1(new_n257), .C2(new_n366), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n456), .A2(new_n378), .A3(new_n499), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n496), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n497), .B1(new_n496), .B2(new_n500), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT28), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n496), .A2(new_n497), .A3(new_n500), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT28), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT68), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n504), .A2(KEYINPUT68), .A3(new_n505), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n503), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n187), .A2(G210), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(KEYINPUT27), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT26), .B(G101), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n510), .A2(KEYINPUT69), .A3(KEYINPUT29), .A4(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT69), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n503), .A2(new_n508), .A3(new_n509), .A4(new_n514), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT29), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n514), .ZN(new_n520));
  INV_X1    g334(.A(new_n375), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n521), .A2(new_n205), .B1(new_n494), .B2(new_n379), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n345), .B1(new_n522), .B2(new_n377), .ZN(new_n523));
  INV_X1    g337(.A(new_n500), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT30), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT30), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n496), .A2(new_n526), .A3(new_n500), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n497), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n520), .B1(new_n528), .B2(new_n501), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n517), .A2(new_n529), .A3(new_n518), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n515), .A2(new_n519), .A3(new_n243), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G472), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT32), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n496), .A2(new_n526), .A3(new_n500), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n526), .B1(new_n496), .B2(new_n500), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n444), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT31), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n504), .A2(new_n514), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT67), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n536), .A2(new_n539), .A3(KEYINPUT67), .A4(new_n537), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n503), .A2(new_n508), .A3(new_n509), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n536), .A2(new_n539), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n545), .A2(new_n520), .B1(new_n546), .B2(KEYINPUT31), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(G472), .A2(G902), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n533), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n549), .ZN(new_n551));
  AOI211_X1 g365(.A(KEYINPUT32), .B(new_n551), .C1(new_n544), .C2(new_n547), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n532), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n317), .A2(G221), .A3(G234), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT71), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT22), .B(G137), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n555), .B(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT70), .B1(new_n419), .B2(G128), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT23), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n249), .A2(G119), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT23), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(KEYINPUT70), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n419), .A2(G128), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n559), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(G110), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n560), .A2(new_n563), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT24), .B(G110), .ZN(new_n567));
  OR2_X1    g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n202), .A2(G146), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n565), .B(new_n568), .C1(new_n569), .C2(new_n226), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT72), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n566), .A2(new_n567), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n572), .B1(new_n564), .B2(G110), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n223), .A2(new_n224), .A3(new_n196), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n202), .B2(G146), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n570), .A2(new_n571), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n571), .B1(new_n570), .B2(new_n576), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n557), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n570), .A2(new_n576), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT72), .ZN(new_n581));
  INV_X1    g395(.A(new_n557), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n579), .A2(new_n243), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT73), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT25), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n270), .B1(G234), .B2(new_n243), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n584), .A2(new_n586), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n579), .A2(KEYINPUT25), .A3(new_n583), .A4(new_n243), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(KEYINPUT73), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n588), .A2(G902), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n579), .A2(new_n583), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n553), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n492), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(new_n333), .ZN(G3));
  AOI21_X1  g414(.A(G902), .B1(new_n544), .B2(new_n547), .ZN(new_n601));
  NAND2_X1  g415(.A1(KEYINPUT91), .A2(G472), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n410), .A2(new_n415), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n313), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n603), .A2(new_n605), .A3(new_n596), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n483), .B1(new_n487), .B2(new_n478), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT93), .B(G478), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n294), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT92), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT33), .B1(new_n290), .B2(new_n293), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n268), .B1(new_n283), .B2(new_n288), .ZN(new_n612));
  INV_X1    g426(.A(new_n271), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n614), .A2(new_n615), .A3(new_n289), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n295), .A2(G902), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n610), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n618), .ZN(new_n620));
  AOI211_X1 g434(.A(KEYINPUT92), .B(new_n620), .C1(new_n611), .C2(new_n616), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n609), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(KEYINPUT94), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n290), .A2(new_n293), .A3(KEYINPUT33), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n615), .B1(new_n614), .B2(new_n289), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n618), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT92), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n617), .A2(new_n610), .A3(new_n618), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT94), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n629), .A2(new_n630), .A3(new_n609), .ZN(new_n631));
  AOI211_X1 g445(.A(new_n247), .B(new_n306), .C1(new_n623), .C2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n606), .A2(new_n607), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G104), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT95), .B(KEYINPUT34), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  INV_X1    g450(.A(KEYINPUT96), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n246), .A2(G475), .ZN(new_n638));
  INV_X1    g452(.A(new_n242), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n241), .B1(new_n240), .B2(new_n232), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n638), .B(new_n297), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n637), .B1(new_n641), .B2(new_n306), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n247), .A2(KEYINPUT96), .A3(new_n297), .A4(new_n305), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n606), .A2(new_n607), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT35), .B(G107), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G9));
  INV_X1    g461(.A(new_n594), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n557), .A2(KEYINPUT36), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n649), .A2(KEYINPUT97), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(KEYINPUT97), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n580), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n650), .A2(new_n570), .A3(new_n576), .A4(new_n651), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n648), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n589), .B2(new_n592), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n603), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n657), .B(new_n417), .C1(new_n491), .C2(new_n484), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT98), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT37), .B(G110), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  NAND2_X1  g475(.A1(new_n525), .A2(new_n527), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n538), .B1(new_n662), .B2(new_n444), .ZN(new_n663));
  AOI21_X1  g477(.A(KEYINPUT67), .B1(new_n663), .B2(new_n537), .ZN(new_n664));
  NOR4_X1   g478(.A1(new_n528), .A2(new_n541), .A3(KEYINPUT31), .A4(new_n538), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n546), .A2(KEYINPUT31), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n667), .B1(new_n510), .B2(new_n514), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n549), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT32), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n551), .B1(new_n544), .B2(new_n547), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n533), .ZN(new_n672));
  AOI22_X1  g486(.A1(new_n670), .A2(new_n672), .B1(G472), .B2(new_n531), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n605), .ZN(new_n674));
  OR2_X1    g488(.A1(new_n303), .A2(G900), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n301), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n641), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n653), .A2(new_n654), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n594), .ZN(new_n680));
  INV_X1    g494(.A(new_n592), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n587), .A2(new_n588), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n607), .A2(new_n678), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n674), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  INV_X1    g500(.A(KEYINPUT102), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n490), .B(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n297), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n234), .A2(new_n242), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n690), .B1(new_n691), .B2(new_n638), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n656), .A2(new_n482), .A3(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n520), .B1(new_n536), .B2(new_n504), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n501), .A2(new_n502), .A3(new_n514), .ZN(new_n697));
  OAI21_X1  g511(.A(KEYINPUT100), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT100), .ZN(new_n699));
  INV_X1    g513(.A(new_n697), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n528), .A2(new_n501), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n699), .B(new_n700), .C1(new_n701), .C2(new_n520), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n698), .A2(new_n702), .A3(new_n243), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(G472), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(KEYINPUT101), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT101), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n703), .A2(new_n706), .A3(G472), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n705), .B(new_n707), .C1(new_n550), .C2(new_n552), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n695), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n676), .B(KEYINPUT39), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n605), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT40), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n687), .B1(new_n709), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n712), .B(KEYINPUT40), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n716), .A2(KEYINPUT102), .A3(new_n708), .A4(new_n695), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n253), .ZN(G45));
  INV_X1    g533(.A(new_n247), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n630), .B1(new_n629), .B2(new_n609), .ZN(new_n721));
  INV_X1    g535(.A(new_n609), .ZN(new_n722));
  AOI211_X1 g536(.A(KEYINPUT94), .B(new_n722), .C1(new_n627), .C2(new_n628), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n720), .B(new_n676), .C1(new_n721), .C2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n607), .A2(new_n683), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n674), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G146), .ZN(G48));
  NAND2_X1  g542(.A1(new_n362), .A2(new_n364), .ZN(new_n729));
  AOI211_X1 g543(.A(KEYINPUT78), .B(new_n382), .C1(new_n729), .C2(new_n391), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n395), .B1(new_n394), .B2(new_n381), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n398), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n406), .A2(new_n407), .ZN(new_n733));
  INV_X1    g547(.A(new_n408), .ZN(new_n734));
  AOI22_X1  g548(.A1(new_n732), .A2(new_n319), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(G469), .B1(new_n735), .B2(G902), .ZN(new_n736));
  AND4_X1   g550(.A1(new_n313), .A2(new_n607), .A3(new_n736), .A4(new_n410), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n737), .A2(new_n553), .A3(new_n597), .A4(new_n632), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT41), .B(G113), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT103), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n738), .B(new_n740), .ZN(G15));
  NAND4_X1  g555(.A1(new_n737), .A2(new_n553), .A3(new_n597), .A4(new_n644), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G116), .ZN(G18));
  AOI21_X1  g557(.A(new_n656), .B1(new_n310), .B2(new_n311), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n737), .A2(new_n553), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G119), .ZN(G21));
  INV_X1    g560(.A(KEYINPUT104), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n671), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(G472), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n601), .A2(new_n749), .ZN(new_n750));
  AOI211_X1 g564(.A(KEYINPUT104), .B(new_n551), .C1(new_n544), .C2(new_n547), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n748), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n736), .A2(new_n313), .A3(new_n410), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n487), .A2(new_n478), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(new_n692), .A3(new_n482), .A4(new_n305), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n752), .A2(new_n597), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G122), .ZN(G24));
  INV_X1    g572(.A(new_n724), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n752), .A2(new_n683), .A3(new_n759), .A4(new_n737), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G125), .ZN(G27));
  INV_X1    g575(.A(KEYINPUT106), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n762), .B1(new_n673), .B2(new_n596), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n478), .A2(new_n482), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n488), .A2(new_n764), .A3(new_n489), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT105), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n488), .A2(new_n764), .A3(KEYINPUT105), .A4(new_n489), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n767), .A2(new_n416), .A3(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n553), .A2(KEYINPUT106), .A3(new_n597), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT42), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n724), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n763), .A2(new_n769), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n767), .A2(new_n416), .A3(new_n768), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n774), .A2(new_n598), .A3(new_n724), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n773), .B1(new_n775), .B2(KEYINPUT42), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G131), .ZN(G33));
  NAND2_X1  g591(.A1(new_n670), .A2(new_n672), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n596), .B1(new_n778), .B2(new_n532), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n769), .A2(new_n779), .A3(new_n678), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT107), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT107), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n769), .A2(new_n779), .A3(new_n782), .A4(new_n678), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G134), .ZN(G36));
  NAND2_X1  g599(.A1(new_n623), .A2(new_n631), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n247), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT43), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n601), .A2(new_n602), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n601), .A2(new_n602), .ZN(new_n791));
  OAI211_X1 g605(.A(KEYINPUT108), .B(new_n683), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT108), .B1(new_n603), .B2(new_n683), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n789), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT44), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n410), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n397), .A2(new_n413), .ZN(new_n799));
  INV_X1    g613(.A(new_n412), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(KEYINPUT45), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT45), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n407), .B1(new_n383), .B2(new_n396), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n802), .B1(new_n803), .B2(new_n412), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n801), .A2(new_n804), .A3(G469), .ZN(new_n805));
  NAND2_X1  g619(.A1(G469), .A2(G902), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT46), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n798), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n805), .A2(KEYINPUT46), .A3(new_n806), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n313), .A3(new_n710), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n767), .A2(new_n768), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n789), .B(KEYINPUT44), .C1(new_n793), .C2(new_n794), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n797), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G137), .ZN(G39));
  NOR4_X1   g631(.A1(new_n813), .A2(new_n553), .A3(new_n597), .A4(new_n724), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT47), .B1(new_n811), .B2(new_n313), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT47), .ZN(new_n820));
  AOI211_X1 g634(.A(new_n820), .B(new_n314), .C1(new_n809), .C2(new_n810), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n818), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G140), .ZN(G42));
  INV_X1    g637(.A(new_n301), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n789), .A2(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n825), .A2(new_n753), .A3(new_n813), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n763), .A2(new_n770), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n826), .A2(KEYINPUT48), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n752), .A2(new_n597), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n737), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n708), .A2(new_n596), .A3(new_n301), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n247), .B1(new_n623), .B2(new_n631), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n813), .A2(new_n753), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n831), .A2(new_n299), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT48), .B1(new_n826), .B2(new_n827), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n753), .A2(new_n482), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n689), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n830), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(KEYINPUT113), .A2(KEYINPUT50), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n832), .A2(new_n834), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n845), .A2(new_n720), .A3(new_n786), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n752), .A2(new_n683), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n846), .B1(new_n847), .B2(new_n826), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n839), .B1(new_n844), .B2(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n825), .A2(new_n829), .A3(new_n813), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n819), .A2(new_n821), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n736), .A2(new_n410), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n313), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n850), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n854), .B1(new_n855), .B2(KEYINPUT51), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n828), .B(new_n838), .C1(new_n849), .C2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n844), .A2(new_n848), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n844), .A2(new_n848), .A3(KEYINPUT114), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n854), .A2(new_n855), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n857), .B1(new_n839), .B2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n757), .A2(new_n738), .A3(new_n742), .A4(new_n745), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n750), .A2(new_n751), .ZN(new_n866));
  INV_X1    g680(.A(new_n748), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n759), .A2(new_n866), .A3(new_n683), .A4(new_n867), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n720), .A2(new_n297), .A3(new_n677), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n553), .A2(new_n683), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n774), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n865), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n784), .A2(new_n776), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n632), .B1(new_n484), .B2(new_n491), .ZN(new_n874));
  INV_X1    g688(.A(new_n641), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n305), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n481), .B1(new_n480), .B2(new_n483), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n490), .A2(KEYINPUT84), .A3(new_n482), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT109), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n874), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI211_X1 g695(.A(KEYINPUT109), .B(new_n876), .C1(new_n877), .C2(new_n878), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n606), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n658), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n599), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  AOI211_X1 g700(.A(new_n677), .B(new_n655), .C1(new_n589), .C2(new_n592), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n604), .A2(new_n887), .A3(new_n313), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT111), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT111), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n416), .A2(new_n890), .A3(new_n887), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n607), .A2(new_n692), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n889), .A2(new_n708), .A3(new_n891), .A4(new_n893), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n553), .B(new_n416), .C1(new_n726), .C2(new_n684), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n895), .A3(new_n760), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT52), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT52), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n894), .A2(new_n895), .A3(new_n760), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n873), .A2(new_n886), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT53), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n784), .A2(new_n776), .A3(new_n872), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n904), .A2(new_n900), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT53), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n906), .A3(new_n886), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n901), .A2(KEYINPUT110), .A3(new_n906), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n902), .A2(KEYINPUT110), .A3(new_n906), .A4(new_n901), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT54), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT54), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n906), .B1(new_n905), .B2(new_n886), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n883), .A2(new_n885), .ZN(new_n915));
  NOR4_X1   g729(.A1(new_n904), .A2(new_n915), .A3(new_n900), .A4(KEYINPUT53), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n913), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n864), .A2(new_n912), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(G952), .A2(G953), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT115), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n597), .A2(new_n482), .A3(new_n313), .ZN(new_n922));
  AOI211_X1 g736(.A(new_n787), .B(new_n922), .C1(KEYINPUT49), .C2(new_n852), .ZN(new_n923));
  INV_X1    g737(.A(new_n708), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n852), .A2(KEYINPUT49), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n923), .A2(new_n924), .A3(new_n689), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n921), .A2(new_n926), .ZN(G75));
  NAND2_X1  g741(.A1(new_n298), .A2(G953), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT118), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n914), .A2(new_n916), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n931), .A2(G210), .A3(G902), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT56), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n454), .B1(new_n462), .B2(new_n463), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT116), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n460), .B(KEYINPUT55), .Z(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n930), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n908), .A2(new_n243), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT117), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n940), .A2(new_n941), .A3(G210), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n932), .A2(KEYINPUT117), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n938), .A2(KEYINPUT56), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n939), .A2(new_n945), .ZN(G51));
  NAND2_X1  g760(.A1(new_n931), .A2(G902), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(new_n805), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n735), .B(KEYINPUT119), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n903), .A2(KEYINPUT54), .A3(new_n907), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n917), .A2(new_n950), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n806), .B(KEYINPUT57), .Z(new_n952));
  AOI21_X1  g766(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n948), .B1(new_n953), .B2(KEYINPUT120), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT120), .ZN(new_n955));
  INV_X1    g769(.A(new_n952), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n917), .B2(new_n950), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n955), .B1(new_n957), .B2(new_n949), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n930), .B1(new_n954), .B2(new_n958), .ZN(G54));
  NAND4_X1  g773(.A1(new_n940), .A2(KEYINPUT58), .A3(G475), .A4(new_n231), .ZN(new_n960));
  NAND2_X1  g774(.A1(KEYINPUT58), .A2(G475), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n240), .B1(new_n947), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n930), .B1(new_n960), .B2(new_n962), .ZN(G60));
  XNOR2_X1  g777(.A(new_n617), .B(KEYINPUT121), .ZN(new_n964));
  NAND2_X1  g778(.A1(G478), .A2(G902), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT59), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n951), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n929), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n912), .A2(new_n917), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n966), .ZN(new_n970));
  INV_X1    g784(.A(new_n964), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(G63));
  NAND2_X1  g786(.A1(new_n579), .A2(new_n583), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT122), .Z(new_n974));
  NAND2_X1  g788(.A1(G217), .A2(G902), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT60), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n974), .B1(new_n908), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n976), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n903), .A2(new_n907), .A3(new_n679), .A4(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n977), .A2(new_n929), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n979), .A2(KEYINPUT123), .A3(new_n929), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(KEYINPUT61), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n980), .B(new_n982), .ZN(G66));
  AOI21_X1  g797(.A(new_n317), .B1(new_n302), .B2(G224), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n915), .A2(new_n865), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(new_n317), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n936), .B1(G898), .B2(new_n317), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT124), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n986), .B(new_n988), .ZN(G69));
  NAND2_X1  g803(.A1(new_n895), .A2(new_n760), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n769), .A2(new_n779), .A3(new_n759), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n771), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n990), .B1(new_n992), .B2(new_n773), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n816), .A2(new_n993), .ZN(new_n994));
  AOI211_X1 g808(.A(new_n314), .B(new_n711), .C1(new_n809), .C2(new_n810), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n995), .A2(new_n893), .A3(new_n763), .A4(new_n770), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n784), .A2(new_n822), .A3(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT126), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n994), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n816), .A2(new_n993), .ZN(new_n1001));
  OAI21_X1  g815(.A(KEYINPUT126), .B1(new_n1001), .B2(new_n997), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n317), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT127), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n317), .A2(G900), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(G953), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1009));
  OAI21_X1  g823(.A(KEYINPUT127), .B1(new_n1009), .B2(new_n1006), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n662), .B(new_n227), .Z(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1008), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n990), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n715), .A2(new_n717), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(KEYINPUT62), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT62), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n715), .A2(new_n717), .A3(new_n1014), .A4(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n710), .B1(new_n833), .B2(new_n875), .ZN(new_n1020));
  NOR3_X1   g834(.A1(new_n774), .A2(new_n598), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1021), .B1(new_n851), .B2(new_n818), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1019), .A2(new_n816), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n317), .B1(new_n1017), .B2(new_n1023), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n1024), .A2(KEYINPUT125), .A3(new_n1011), .ZN(new_n1025));
  AOI21_X1  g839(.A(KEYINPUT125), .B1(new_n1024), .B2(new_n1011), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n317), .B1(G227), .B2(G900), .ZN(new_n1028));
  AND3_X1   g842(.A1(new_n1013), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1028), .B1(new_n1013), .B2(new_n1027), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1029), .A2(new_n1030), .ZN(G72));
  NAND2_X1  g845(.A1(G472), .A2(G902), .ZN(new_n1032));
  XOR2_X1   g846(.A(new_n1032), .B(KEYINPUT63), .Z(new_n1033));
  OR2_X1    g847(.A1(new_n1017), .A2(new_n1023), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1033), .B1(new_n1034), .B2(new_n985), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1035), .A2(new_n696), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1033), .B1(new_n1003), .B2(new_n985), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1037), .A2(new_n520), .A3(new_n701), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1036), .A2(new_n929), .A3(new_n1038), .ZN(new_n1039));
  AND2_X1   g853(.A1(new_n910), .A2(new_n911), .ZN(new_n1040));
  INV_X1    g854(.A(new_n1033), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1041), .B1(new_n529), .B2(new_n546), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1039), .B1(new_n1040), .B2(new_n1042), .ZN(G57));
endmodule


