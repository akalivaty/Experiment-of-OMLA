

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U556 ( .A1(n538), .A2(n537), .ZN(G160) );
  NOR2_X2 U557 ( .A1(n546), .A2(n545), .ZN(G164) );
  XOR2_X1 U558 ( .A(KEYINPUT95), .B(n600), .Z(n710) );
  NOR2_X1 U559 ( .A1(n659), .A2(n934), .ZN(n604) );
  BUF_X1 U560 ( .A(n908), .Z(n525) );
  AND2_X2 U561 ( .A1(G2105), .A2(G2104), .ZN(n904) );
  XNOR2_X1 U562 ( .A(n529), .B(n528), .ZN(n908) );
  AND2_X1 U563 ( .A1(n618), .A2(n617), .ZN(n629) );
  AND2_X1 U564 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U565 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  NOR2_X1 U566 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U567 ( .A1(n904), .A2(G114), .ZN(n539) );
  XOR2_X1 U568 ( .A(n712), .B(KEYINPUT103), .Z(n526) );
  OR2_X1 U569 ( .A1(n704), .A2(n962), .ZN(n527) );
  NOR2_X2 U570 ( .A1(n735), .A2(n599), .ZN(n653) );
  XNOR2_X1 U571 ( .A(n663), .B(KEYINPUT30), .ZN(n664) );
  INV_X1 U572 ( .A(KEYINPUT31), .ZN(n668) );
  NAND2_X1 U573 ( .A1(n809), .A2(G54), .ZN(n619) );
  NOR2_X1 U574 ( .A1(G164), .A2(G1384), .ZN(n598) );
  XNOR2_X1 U575 ( .A(n622), .B(KEYINPUT76), .ZN(n626) );
  XOR2_X1 U576 ( .A(KEYINPUT0), .B(G543), .Z(n583) );
  INV_X1 U577 ( .A(KEYINPUT17), .ZN(n528) );
  NOR2_X2 U578 ( .A1(G651), .A2(n583), .ZN(n809) );
  NOR2_X1 U579 ( .A1(G651), .A2(G543), .ZN(n813) );
  NAND2_X1 U580 ( .A1(n908), .A2(G138), .ZN(n541) );
  NAND2_X1 U581 ( .A1(n525), .A2(G137), .ZN(n532) );
  INV_X1 U582 ( .A(G2105), .ZN(n533) );
  AND2_X1 U583 ( .A1(n533), .A2(G2104), .ZN(n910) );
  NAND2_X1 U584 ( .A1(G101), .A2(n910), .ZN(n530) );
  XOR2_X1 U585 ( .A(KEYINPUT23), .B(n530), .Z(n531) );
  NAND2_X1 U586 ( .A1(n532), .A2(n531), .ZN(n538) );
  NAND2_X1 U587 ( .A1(G113), .A2(n904), .ZN(n536) );
  NOR2_X1 U588 ( .A1(n533), .A2(G2104), .ZN(n534) );
  XNOR2_X1 U589 ( .A(n534), .B(KEYINPUT66), .ZN(n542) );
  BUF_X1 U590 ( .A(n542), .Z(n905) );
  NAND2_X1 U591 ( .A1(G125), .A2(n905), .ZN(n535) );
  NAND2_X1 U592 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U593 ( .A(n539), .B(KEYINPUT88), .ZN(n540) );
  NAND2_X1 U594 ( .A1(n541), .A2(n540), .ZN(n546) );
  NAND2_X1 U595 ( .A1(G126), .A2(n542), .ZN(n544) );
  NAND2_X1 U596 ( .A1(G102), .A2(n910), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U598 ( .A1(n813), .A2(G86), .ZN(n555) );
  INV_X1 U599 ( .A(G651), .ZN(n550) );
  NOR2_X1 U600 ( .A1(G543), .A2(n550), .ZN(n547) );
  XOR2_X1 U601 ( .A(KEYINPUT1), .B(n547), .Z(n808) );
  NAND2_X1 U602 ( .A1(G61), .A2(n808), .ZN(n549) );
  NAND2_X1 U603 ( .A1(G48), .A2(n809), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n549), .A2(n548), .ZN(n553) );
  NOR2_X1 U605 ( .A1(n583), .A2(n550), .ZN(n812) );
  NAND2_X1 U606 ( .A1(G73), .A2(n812), .ZN(n551) );
  XOR2_X1 U607 ( .A(KEYINPUT2), .B(n551), .Z(n552) );
  NOR2_X1 U608 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U609 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U610 ( .A(n556), .B(KEYINPUT84), .ZN(G305) );
  NAND2_X1 U611 ( .A1(n813), .A2(G90), .ZN(n557) );
  XNOR2_X1 U612 ( .A(n557), .B(KEYINPUT70), .ZN(n559) );
  NAND2_X1 U613 ( .A1(G77), .A2(n812), .ZN(n558) );
  NAND2_X1 U614 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U615 ( .A(n560), .B(KEYINPUT9), .ZN(n562) );
  NAND2_X1 U616 ( .A1(G52), .A2(n809), .ZN(n561) );
  NAND2_X1 U617 ( .A1(n562), .A2(n561), .ZN(n565) );
  NAND2_X1 U618 ( .A1(G64), .A2(n808), .ZN(n563) );
  XNOR2_X1 U619 ( .A(KEYINPUT69), .B(n563), .ZN(n564) );
  NOR2_X1 U620 ( .A1(n565), .A2(n564), .ZN(G171) );
  NAND2_X1 U621 ( .A1(n813), .A2(G89), .ZN(n566) );
  XNOR2_X1 U622 ( .A(n566), .B(KEYINPUT4), .ZN(n568) );
  NAND2_X1 U623 ( .A1(G76), .A2(n812), .ZN(n567) );
  NAND2_X1 U624 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U625 ( .A(n569), .B(KEYINPUT5), .ZN(n575) );
  XNOR2_X1 U626 ( .A(KEYINPUT6), .B(KEYINPUT77), .ZN(n573) );
  NAND2_X1 U627 ( .A1(G63), .A2(n808), .ZN(n571) );
  NAND2_X1 U628 ( .A1(G51), .A2(n809), .ZN(n570) );
  NAND2_X1 U629 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U630 ( .A(n573), .B(n572), .ZN(n574) );
  NAND2_X1 U631 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U632 ( .A(KEYINPUT7), .B(n576), .ZN(G168) );
  XOR2_X1 U633 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U634 ( .A1(G75), .A2(n812), .ZN(n578) );
  NAND2_X1 U635 ( .A1(G88), .A2(n813), .ZN(n577) );
  NAND2_X1 U636 ( .A1(n578), .A2(n577), .ZN(n582) );
  NAND2_X1 U637 ( .A1(G62), .A2(n808), .ZN(n580) );
  NAND2_X1 U638 ( .A1(G50), .A2(n809), .ZN(n579) );
  NAND2_X1 U639 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U640 ( .A1(n582), .A2(n581), .ZN(G166) );
  INV_X1 U641 ( .A(G166), .ZN(G303) );
  NAND2_X1 U642 ( .A1(G651), .A2(G74), .ZN(n588) );
  NAND2_X1 U643 ( .A1(G49), .A2(n809), .ZN(n585) );
  NAND2_X1 U644 ( .A1(G87), .A2(n583), .ZN(n584) );
  NAND2_X1 U645 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U646 ( .A1(n808), .A2(n586), .ZN(n587) );
  NAND2_X1 U647 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U648 ( .A(KEYINPUT83), .B(n589), .Z(G288) );
  NAND2_X1 U649 ( .A1(n809), .A2(G47), .ZN(n590) );
  XOR2_X1 U650 ( .A(KEYINPUT67), .B(n590), .Z(n592) );
  NAND2_X1 U651 ( .A1(n808), .A2(G60), .ZN(n591) );
  NAND2_X1 U652 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U653 ( .A(KEYINPUT68), .B(n593), .Z(n597) );
  NAND2_X1 U654 ( .A1(n812), .A2(G72), .ZN(n595) );
  NAND2_X1 U655 ( .A1(G85), .A2(n813), .ZN(n594) );
  AND2_X1 U656 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U657 ( .A1(n597), .A2(n596), .ZN(G290) );
  NAND2_X1 U658 ( .A1(G160), .A2(G40), .ZN(n735) );
  XNOR2_X1 U659 ( .A(n598), .B(KEYINPUT64), .ZN(n736) );
  INV_X1 U660 ( .A(n736), .ZN(n599) );
  INV_X1 U661 ( .A(n653), .ZN(n659) );
  NAND2_X1 U662 ( .A1(n659), .A2(G8), .ZN(n600) );
  NOR2_X1 U663 ( .A1(G1981), .A2(G305), .ZN(n601) );
  XOR2_X1 U664 ( .A(n601), .B(KEYINPUT24), .Z(n602) );
  NOR2_X1 U665 ( .A1(n710), .A2(n602), .ZN(n715) );
  XNOR2_X1 U666 ( .A(KEYINPUT29), .B(KEYINPUT98), .ZN(n652) );
  XOR2_X1 U667 ( .A(KEYINPUT96), .B(G1996), .Z(n934) );
  XNOR2_X1 U668 ( .A(KEYINPUT65), .B(KEYINPUT26), .ZN(n603) );
  XNOR2_X1 U669 ( .A(n604), .B(n603), .ZN(n618) );
  AND2_X1 U670 ( .A1(n659), .A2(G1341), .ZN(n616) );
  NAND2_X1 U671 ( .A1(n809), .A2(G43), .ZN(n605) );
  XNOR2_X1 U672 ( .A(KEYINPUT74), .B(n605), .ZN(n615) );
  XNOR2_X1 U673 ( .A(KEYINPUT13), .B(KEYINPUT73), .ZN(n610) );
  NAND2_X1 U674 ( .A1(n813), .A2(G81), .ZN(n606) );
  XNOR2_X1 U675 ( .A(n606), .B(KEYINPUT12), .ZN(n608) );
  NAND2_X1 U676 ( .A1(G68), .A2(n812), .ZN(n607) );
  NAND2_X1 U677 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U678 ( .A(n610), .B(n609), .ZN(n613) );
  NAND2_X1 U679 ( .A1(n808), .A2(G56), .ZN(n611) );
  XOR2_X1 U680 ( .A(KEYINPUT14), .B(n611), .Z(n612) );
  NOR2_X1 U681 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U682 ( .A1(n615), .A2(n614), .ZN(n954) );
  NOR2_X1 U683 ( .A1(n616), .A2(n954), .ZN(n617) );
  XOR2_X1 U684 ( .A(KEYINPUT75), .B(n619), .Z(n621) );
  NAND2_X1 U685 ( .A1(n812), .A2(G79), .ZN(n620) );
  NAND2_X1 U686 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U687 ( .A1(G66), .A2(n808), .ZN(n624) );
  NAND2_X1 U688 ( .A1(G92), .A2(n813), .ZN(n623) );
  NAND2_X1 U689 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X2 U690 ( .A(KEYINPUT15), .B(n627), .Z(n968) );
  NOR2_X1 U691 ( .A1(n629), .A2(n968), .ZN(n628) );
  XNOR2_X1 U692 ( .A(n628), .B(KEYINPUT97), .ZN(n635) );
  NAND2_X1 U693 ( .A1(n629), .A2(n968), .ZN(n633) );
  NOR2_X1 U694 ( .A1(n653), .A2(G1348), .ZN(n631) );
  NOR2_X1 U695 ( .A1(G2067), .A2(n659), .ZN(n630) );
  NOR2_X1 U696 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U697 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U698 ( .A1(n635), .A2(n634), .ZN(n646) );
  NAND2_X1 U699 ( .A1(G65), .A2(n808), .ZN(n637) );
  NAND2_X1 U700 ( .A1(G53), .A2(n809), .ZN(n636) );
  NAND2_X1 U701 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U702 ( .A1(G78), .A2(n812), .ZN(n639) );
  NAND2_X1 U703 ( .A1(G91), .A2(n813), .ZN(n638) );
  NAND2_X1 U704 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U705 ( .A1(n641), .A2(n640), .ZN(n951) );
  NAND2_X1 U706 ( .A1(n653), .A2(G2072), .ZN(n642) );
  XNOR2_X1 U707 ( .A(n642), .B(KEYINPUT27), .ZN(n644) );
  INV_X1 U708 ( .A(G1956), .ZN(n986) );
  NOR2_X1 U709 ( .A1(n986), .A2(n653), .ZN(n643) );
  NOR2_X1 U710 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U711 ( .A1(n951), .A2(n647), .ZN(n645) );
  NAND2_X1 U712 ( .A1(n646), .A2(n645), .ZN(n650) );
  NOR2_X1 U713 ( .A1(n951), .A2(n647), .ZN(n648) );
  XOR2_X1 U714 ( .A(n648), .B(KEYINPUT28), .Z(n649) );
  NAND2_X1 U715 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U716 ( .A(n652), .B(n651), .ZN(n657) );
  XNOR2_X1 U717 ( .A(KEYINPUT25), .B(G2078), .ZN(n935) );
  NOR2_X1 U718 ( .A1(n659), .A2(n935), .ZN(n655) );
  AND2_X1 U719 ( .A1(n659), .A2(G1961), .ZN(n654) );
  NOR2_X1 U720 ( .A1(n655), .A2(n654), .ZN(n665) );
  AND2_X1 U721 ( .A1(G171), .A2(n665), .ZN(n656) );
  NOR2_X2 U722 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U723 ( .A(n658), .B(KEYINPUT99), .ZN(n681) );
  OR2_X1 U724 ( .A1(G1966), .A2(n710), .ZN(n662) );
  NOR2_X1 U725 ( .A1(G2084), .A2(n659), .ZN(n682) );
  INV_X1 U726 ( .A(G8), .ZN(n660) );
  NOR2_X1 U727 ( .A1(n682), .A2(n660), .ZN(n661) );
  NAND2_X1 U728 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U729 ( .A1(n664), .A2(G168), .ZN(n667) );
  NOR2_X1 U730 ( .A1(G171), .A2(n665), .ZN(n666) );
  NOR2_X1 U731 ( .A1(n667), .A2(n666), .ZN(n669) );
  XNOR2_X1 U732 ( .A(n669), .B(n668), .ZN(n680) );
  NAND2_X1 U733 ( .A1(n681), .A2(n680), .ZN(n671) );
  AND2_X1 U734 ( .A1(G286), .A2(G8), .ZN(n670) );
  NAND2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n678) );
  NOR2_X1 U736 ( .A1(G1971), .A2(n710), .ZN(n673) );
  NOR2_X1 U737 ( .A1(G2090), .A2(n659), .ZN(n672) );
  NOR2_X1 U738 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U739 ( .A(n674), .B(KEYINPUT100), .ZN(n675) );
  NAND2_X1 U740 ( .A1(n675), .A2(G303), .ZN(n676) );
  OR2_X1 U741 ( .A1(n660), .A2(n676), .ZN(n677) );
  XNOR2_X1 U742 ( .A(n679), .B(KEYINPUT32), .ZN(n705) );
  AND2_X1 U743 ( .A1(n681), .A2(n680), .ZN(n686) );
  AND2_X1 U744 ( .A1(G8), .A2(n682), .ZN(n684) );
  NOR2_X1 U745 ( .A1(G1966), .A2(n710), .ZN(n683) );
  OR2_X1 U746 ( .A1(n684), .A2(n683), .ZN(n685) );
  OR2_X1 U747 ( .A1(n686), .A2(n685), .ZN(n706) );
  NOR2_X1 U748 ( .A1(G1976), .A2(G288), .ZN(n696) );
  INV_X1 U749 ( .A(n710), .ZN(n689) );
  NAND2_X1 U750 ( .A1(n696), .A2(n689), .ZN(n687) );
  NAND2_X1 U751 ( .A1(n687), .A2(KEYINPUT33), .ZN(n697) );
  INV_X1 U752 ( .A(n697), .ZN(n692) );
  INV_X1 U753 ( .A(KEYINPUT33), .ZN(n688) );
  NAND2_X1 U754 ( .A1(G1976), .A2(G288), .ZN(n959) );
  AND2_X1 U755 ( .A1(n688), .A2(n959), .ZN(n690) );
  AND2_X1 U756 ( .A1(n690), .A2(n689), .ZN(n691) );
  OR2_X1 U757 ( .A1(n692), .A2(n691), .ZN(n694) );
  AND2_X1 U758 ( .A1(n706), .A2(n694), .ZN(n693) );
  NAND2_X1 U759 ( .A1(n705), .A2(n693), .ZN(n701) );
  INV_X1 U760 ( .A(n694), .ZN(n699) );
  NOR2_X1 U761 ( .A1(G1971), .A2(G303), .ZN(n695) );
  NOR2_X1 U762 ( .A1(n696), .A2(n695), .ZN(n956) );
  AND2_X1 U763 ( .A1(n956), .A2(n697), .ZN(n698) );
  OR2_X1 U764 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U765 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U766 ( .A(n702), .B(KEYINPUT101), .ZN(n704) );
  XNOR2_X1 U767 ( .A(G1981), .B(G305), .ZN(n703) );
  XNOR2_X1 U768 ( .A(n703), .B(KEYINPUT102), .ZN(n962) );
  NAND2_X1 U769 ( .A1(n706), .A2(n705), .ZN(n709) );
  NOR2_X1 U770 ( .A1(G2090), .A2(G303), .ZN(n707) );
  NAND2_X1 U771 ( .A1(G8), .A2(n707), .ZN(n708) );
  NAND2_X1 U772 ( .A1(n709), .A2(n708), .ZN(n711) );
  NAND2_X1 U773 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U774 ( .A1(n527), .A2(n526), .ZN(n713) );
  XNOR2_X1 U775 ( .A(n713), .B(KEYINPUT104), .ZN(n714) );
  NOR2_X1 U776 ( .A1(n715), .A2(n714), .ZN(n749) );
  NAND2_X1 U777 ( .A1(G131), .A2(n525), .ZN(n717) );
  NAND2_X1 U778 ( .A1(G95), .A2(n910), .ZN(n716) );
  NAND2_X1 U779 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U780 ( .A(KEYINPUT92), .B(n718), .ZN(n723) );
  NAND2_X1 U781 ( .A1(G107), .A2(n904), .ZN(n720) );
  NAND2_X1 U782 ( .A1(G119), .A2(n905), .ZN(n719) );
  NAND2_X1 U783 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U784 ( .A(KEYINPUT91), .B(n721), .Z(n722) );
  NOR2_X1 U785 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U786 ( .A(KEYINPUT93), .B(n724), .ZN(n896) );
  NAND2_X1 U787 ( .A1(n896), .A2(G1991), .ZN(n734) );
  NAND2_X1 U788 ( .A1(n905), .A2(G129), .ZN(n731) );
  NAND2_X1 U789 ( .A1(G117), .A2(n904), .ZN(n726) );
  NAND2_X1 U790 ( .A1(G141), .A2(n525), .ZN(n725) );
  NAND2_X1 U791 ( .A1(n726), .A2(n725), .ZN(n729) );
  NAND2_X1 U792 ( .A1(n910), .A2(G105), .ZN(n727) );
  XOR2_X1 U793 ( .A(KEYINPUT38), .B(n727), .Z(n728) );
  NOR2_X1 U794 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U795 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U796 ( .A(n732), .B(KEYINPUT94), .ZN(n901) );
  NAND2_X1 U797 ( .A1(n901), .A2(G1996), .ZN(n733) );
  NAND2_X1 U798 ( .A1(n734), .A2(n733), .ZN(n1016) );
  NOR2_X1 U799 ( .A1(n736), .A2(n735), .ZN(n764) );
  NAND2_X1 U800 ( .A1(n1016), .A2(n764), .ZN(n752) );
  XNOR2_X1 U801 ( .A(G2067), .B(KEYINPUT37), .ZN(n761) );
  NAND2_X1 U802 ( .A1(n910), .A2(G104), .ZN(n737) );
  XOR2_X1 U803 ( .A(KEYINPUT89), .B(n737), .Z(n739) );
  NAND2_X1 U804 ( .A1(n525), .A2(G140), .ZN(n738) );
  NAND2_X1 U805 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U806 ( .A(KEYINPUT34), .B(n740), .ZN(n746) );
  NAND2_X1 U807 ( .A1(G116), .A2(n904), .ZN(n742) );
  NAND2_X1 U808 ( .A1(G128), .A2(n905), .ZN(n741) );
  NAND2_X1 U809 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U810 ( .A(KEYINPUT90), .B(n743), .Z(n744) );
  XNOR2_X1 U811 ( .A(KEYINPUT35), .B(n744), .ZN(n745) );
  NOR2_X1 U812 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U813 ( .A(KEYINPUT36), .B(n747), .ZN(n918) );
  NOR2_X1 U814 ( .A1(n761), .A2(n918), .ZN(n1023) );
  NAND2_X1 U815 ( .A1(n764), .A2(n1023), .ZN(n759) );
  NAND2_X1 U816 ( .A1(n752), .A2(n759), .ZN(n748) );
  NOR2_X1 U817 ( .A1(n749), .A2(n748), .ZN(n751) );
  XNOR2_X1 U818 ( .A(G1986), .B(G290), .ZN(n973) );
  NAND2_X1 U819 ( .A1(n973), .A2(n764), .ZN(n750) );
  NAND2_X1 U820 ( .A1(n751), .A2(n750), .ZN(n767) );
  NOR2_X1 U821 ( .A1(G1996), .A2(n901), .ZN(n1011) );
  INV_X1 U822 ( .A(n752), .ZN(n755) );
  NOR2_X1 U823 ( .A1(G1986), .A2(G290), .ZN(n753) );
  NOR2_X1 U824 ( .A1(G1991), .A2(n896), .ZN(n1020) );
  NOR2_X1 U825 ( .A1(n753), .A2(n1020), .ZN(n754) );
  NOR2_X1 U826 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U827 ( .A(KEYINPUT105), .B(n756), .Z(n757) );
  NOR2_X1 U828 ( .A1(n1011), .A2(n757), .ZN(n758) );
  XNOR2_X1 U829 ( .A(n758), .B(KEYINPUT39), .ZN(n760) );
  NAND2_X1 U830 ( .A1(n760), .A2(n759), .ZN(n762) );
  NAND2_X1 U831 ( .A1(n761), .A2(n918), .ZN(n1027) );
  NAND2_X1 U832 ( .A1(n762), .A2(n1027), .ZN(n763) );
  NAND2_X1 U833 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U834 ( .A(KEYINPUT106), .B(n765), .ZN(n766) );
  NAND2_X1 U835 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U836 ( .A(n768), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U837 ( .A(G2435), .B(G2427), .ZN(n778) );
  XOR2_X1 U838 ( .A(G2454), .B(G2430), .Z(n770) );
  XNOR2_X1 U839 ( .A(G2443), .B(G2451), .ZN(n769) );
  XNOR2_X1 U840 ( .A(n770), .B(n769), .ZN(n774) );
  XOR2_X1 U841 ( .A(G2446), .B(KEYINPUT107), .Z(n772) );
  XNOR2_X1 U842 ( .A(G1348), .B(G1341), .ZN(n771) );
  XNOR2_X1 U843 ( .A(n772), .B(n771), .ZN(n773) );
  XOR2_X1 U844 ( .A(n774), .B(n773), .Z(n776) );
  XNOR2_X1 U845 ( .A(KEYINPUT108), .B(G2438), .ZN(n775) );
  XNOR2_X1 U846 ( .A(n776), .B(n775), .ZN(n777) );
  XNOR2_X1 U847 ( .A(n778), .B(n777), .ZN(n779) );
  AND2_X1 U848 ( .A1(n779), .A2(G14), .ZN(G401) );
  AND2_X1 U849 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U850 ( .A1(G123), .A2(n905), .ZN(n780) );
  XNOR2_X1 U851 ( .A(n780), .B(KEYINPUT18), .ZN(n782) );
  NAND2_X1 U852 ( .A1(G135), .A2(n525), .ZN(n781) );
  NAND2_X1 U853 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U854 ( .A(KEYINPUT80), .B(n783), .ZN(n786) );
  NAND2_X1 U855 ( .A1(G111), .A2(n904), .ZN(n784) );
  XNOR2_X1 U856 ( .A(KEYINPUT81), .B(n784), .ZN(n785) );
  NOR2_X1 U857 ( .A1(n786), .A2(n785), .ZN(n788) );
  NAND2_X1 U858 ( .A1(n910), .A2(G99), .ZN(n787) );
  NAND2_X1 U859 ( .A1(n788), .A2(n787), .ZN(n1017) );
  XNOR2_X1 U860 ( .A(G2096), .B(n1017), .ZN(n789) );
  OR2_X1 U861 ( .A1(G2100), .A2(n789), .ZN(G156) );
  INV_X1 U862 ( .A(G108), .ZN(G238) );
  INV_X1 U863 ( .A(G120), .ZN(G236) );
  INV_X1 U864 ( .A(G57), .ZN(G237) );
  INV_X1 U865 ( .A(G132), .ZN(G219) );
  NAND2_X1 U866 ( .A1(G7), .A2(G661), .ZN(n790) );
  XNOR2_X1 U867 ( .A(n790), .B(KEYINPUT72), .ZN(n791) );
  XNOR2_X1 U868 ( .A(KEYINPUT10), .B(n791), .ZN(G223) );
  INV_X1 U869 ( .A(G567), .ZN(n841) );
  NOR2_X1 U870 ( .A1(G223), .A2(n841), .ZN(n792) );
  XNOR2_X1 U871 ( .A(n792), .B(KEYINPUT11), .ZN(G234) );
  INV_X1 U872 ( .A(G860), .ZN(n807) );
  OR2_X1 U873 ( .A1(n954), .A2(n807), .ZN(G153) );
  INV_X1 U874 ( .A(G171), .ZN(G301) );
  NAND2_X1 U875 ( .A1(G868), .A2(G301), .ZN(n794) );
  OR2_X1 U876 ( .A1(n968), .A2(G868), .ZN(n793) );
  NAND2_X1 U877 ( .A1(n794), .A2(n793), .ZN(G284) );
  INV_X1 U878 ( .A(n951), .ZN(G299) );
  NOR2_X1 U879 ( .A1(G868), .A2(G299), .ZN(n795) );
  XNOR2_X1 U880 ( .A(n795), .B(KEYINPUT78), .ZN(n798) );
  INV_X1 U881 ( .A(G868), .ZN(n796) );
  NOR2_X1 U882 ( .A1(n796), .A2(G286), .ZN(n797) );
  NOR2_X1 U883 ( .A1(n798), .A2(n797), .ZN(G297) );
  NAND2_X1 U884 ( .A1(n807), .A2(G559), .ZN(n799) );
  NAND2_X1 U885 ( .A1(n799), .A2(n968), .ZN(n800) );
  XNOR2_X1 U886 ( .A(n800), .B(KEYINPUT79), .ZN(n801) );
  XOR2_X1 U887 ( .A(KEYINPUT16), .B(n801), .Z(G148) );
  NOR2_X1 U888 ( .A1(G868), .A2(n954), .ZN(n804) );
  NAND2_X1 U889 ( .A1(G868), .A2(n968), .ZN(n802) );
  NOR2_X1 U890 ( .A1(G559), .A2(n802), .ZN(n803) );
  NOR2_X1 U891 ( .A1(n804), .A2(n803), .ZN(G282) );
  NAND2_X1 U892 ( .A1(G559), .A2(n968), .ZN(n805) );
  XOR2_X1 U893 ( .A(KEYINPUT82), .B(n805), .Z(n806) );
  XNOR2_X1 U894 ( .A(n954), .B(n806), .ZN(n825) );
  NAND2_X1 U895 ( .A1(n807), .A2(n825), .ZN(n818) );
  NAND2_X1 U896 ( .A1(G67), .A2(n808), .ZN(n811) );
  NAND2_X1 U897 ( .A1(G55), .A2(n809), .ZN(n810) );
  NAND2_X1 U898 ( .A1(n811), .A2(n810), .ZN(n817) );
  NAND2_X1 U899 ( .A1(G80), .A2(n812), .ZN(n815) );
  NAND2_X1 U900 ( .A1(G93), .A2(n813), .ZN(n814) );
  NAND2_X1 U901 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U902 ( .A1(n817), .A2(n816), .ZN(n827) );
  XOR2_X1 U903 ( .A(n818), .B(n827), .Z(G145) );
  XNOR2_X1 U904 ( .A(KEYINPUT85), .B(KEYINPUT19), .ZN(n820) );
  XNOR2_X1 U905 ( .A(G288), .B(G166), .ZN(n819) );
  XNOR2_X1 U906 ( .A(n820), .B(n819), .ZN(n821) );
  XOR2_X1 U907 ( .A(n821), .B(n827), .Z(n823) );
  XNOR2_X1 U908 ( .A(G305), .B(n951), .ZN(n822) );
  XNOR2_X1 U909 ( .A(n823), .B(n822), .ZN(n824) );
  XOR2_X1 U910 ( .A(n824), .B(G290), .Z(n856) );
  XNOR2_X1 U911 ( .A(n825), .B(n856), .ZN(n826) );
  NAND2_X1 U912 ( .A1(n826), .A2(G868), .ZN(n829) );
  OR2_X1 U913 ( .A1(n827), .A2(G868), .ZN(n828) );
  NAND2_X1 U914 ( .A1(n829), .A2(n828), .ZN(G295) );
  XOR2_X1 U915 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n831) );
  NAND2_X1 U916 ( .A1(G2084), .A2(G2078), .ZN(n830) );
  XNOR2_X1 U917 ( .A(n831), .B(n830), .ZN(n832) );
  NAND2_X1 U918 ( .A1(G2090), .A2(n832), .ZN(n833) );
  XNOR2_X1 U919 ( .A(KEYINPUT21), .B(n833), .ZN(n834) );
  NAND2_X1 U920 ( .A1(n834), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U921 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U922 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NOR2_X1 U923 ( .A1(G219), .A2(G220), .ZN(n835) );
  XOR2_X1 U924 ( .A(KEYINPUT22), .B(n835), .Z(n836) );
  NOR2_X1 U925 ( .A1(G218), .A2(n836), .ZN(n837) );
  NAND2_X1 U926 ( .A1(G96), .A2(n837), .ZN(n851) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n851), .ZN(n838) );
  XNOR2_X1 U928 ( .A(n838), .B(KEYINPUT87), .ZN(n843) );
  NOR2_X1 U929 ( .A1(G236), .A2(G238), .ZN(n839) );
  NAND2_X1 U930 ( .A1(G69), .A2(n839), .ZN(n840) );
  NOR2_X1 U931 ( .A1(G237), .A2(n840), .ZN(n850) );
  NOR2_X1 U932 ( .A1(n841), .A2(n850), .ZN(n842) );
  NOR2_X1 U933 ( .A1(n843), .A2(n842), .ZN(G319) );
  INV_X1 U934 ( .A(G319), .ZN(n924) );
  NAND2_X1 U935 ( .A1(G483), .A2(G661), .ZN(n844) );
  NOR2_X1 U936 ( .A1(n924), .A2(n844), .ZN(n849) );
  NAND2_X1 U937 ( .A1(n849), .A2(G36), .ZN(G176) );
  INV_X1 U938 ( .A(G223), .ZN(n845) );
  NAND2_X1 U939 ( .A1(G2106), .A2(n845), .ZN(G217) );
  AND2_X1 U940 ( .A1(G15), .A2(G2), .ZN(n846) );
  NAND2_X1 U941 ( .A1(G661), .A2(n846), .ZN(G259) );
  NAND2_X1 U942 ( .A1(G3), .A2(G1), .ZN(n847) );
  XOR2_X1 U943 ( .A(KEYINPUT109), .B(n847), .Z(n848) );
  NAND2_X1 U944 ( .A1(n849), .A2(n848), .ZN(G188) );
  INV_X1 U946 ( .A(G96), .ZN(G221) );
  INV_X1 U947 ( .A(n850), .ZN(n852) );
  NOR2_X1 U948 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U949 ( .A(KEYINPUT110), .B(n853), .ZN(G325) );
  INV_X1 U950 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U951 ( .A(n954), .B(G286), .ZN(n855) );
  XNOR2_X1 U952 ( .A(G171), .B(n968), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n857) );
  XNOR2_X1 U954 ( .A(n857), .B(n856), .ZN(n858) );
  NOR2_X1 U955 ( .A1(G37), .A2(n858), .ZN(G397) );
  XOR2_X1 U956 ( .A(KEYINPUT42), .B(G2090), .Z(n860) );
  XNOR2_X1 U957 ( .A(G2067), .B(G2084), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U959 ( .A(n861), .B(G2100), .Z(n863) );
  XNOR2_X1 U960 ( .A(G2078), .B(G2072), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U962 ( .A(G2096), .B(KEYINPUT43), .Z(n865) );
  XNOR2_X1 U963 ( .A(KEYINPUT111), .B(G2678), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U965 ( .A(n867), .B(n866), .Z(G227) );
  XNOR2_X1 U966 ( .A(G1966), .B(KEYINPUT41), .ZN(n877) );
  XOR2_X1 U967 ( .A(G1956), .B(G1961), .Z(n869) );
  XNOR2_X1 U968 ( .A(G1981), .B(G1971), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n873) );
  XOR2_X1 U970 ( .A(G1991), .B(G1986), .Z(n871) );
  XNOR2_X1 U971 ( .A(G1976), .B(G1996), .ZN(n870) );
  XNOR2_X1 U972 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U973 ( .A(n873), .B(n872), .Z(n875) );
  XNOR2_X1 U974 ( .A(KEYINPUT112), .B(G2474), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U976 ( .A(n877), .B(n876), .ZN(G229) );
  NAND2_X1 U977 ( .A1(G100), .A2(n910), .ZN(n884) );
  NAND2_X1 U978 ( .A1(G112), .A2(n904), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G136), .A2(n525), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n882) );
  NAND2_X1 U981 ( .A1(n905), .A2(G124), .ZN(n880) );
  XOR2_X1 U982 ( .A(KEYINPUT44), .B(n880), .Z(n881) );
  NOR2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U985 ( .A(n885), .B(KEYINPUT113), .ZN(G162) );
  NAND2_X1 U986 ( .A1(G103), .A2(n910), .ZN(n886) );
  XNOR2_X1 U987 ( .A(n886), .B(KEYINPUT116), .ZN(n889) );
  NAND2_X1 U988 ( .A1(G139), .A2(n525), .ZN(n887) );
  XOR2_X1 U989 ( .A(KEYINPUT117), .B(n887), .Z(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n894) );
  NAND2_X1 U991 ( .A1(G115), .A2(n904), .ZN(n891) );
  NAND2_X1 U992 ( .A1(G127), .A2(n905), .ZN(n890) );
  NAND2_X1 U993 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n892), .Z(n893) );
  NOR2_X1 U995 ( .A1(n894), .A2(n893), .ZN(n1006) );
  XOR2_X1 U996 ( .A(G160), .B(n1006), .Z(n895) );
  XNOR2_X1 U997 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U998 ( .A(n897), .B(KEYINPUT115), .Z(n899) );
  XNOR2_X1 U999 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n898) );
  XNOR2_X1 U1000 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U1001 ( .A(n900), .B(G162), .Z(n903) );
  XNOR2_X1 U1002 ( .A(G164), .B(n901), .ZN(n902) );
  XNOR2_X1 U1003 ( .A(n903), .B(n902), .ZN(n917) );
  NAND2_X1 U1004 ( .A1(G118), .A2(n904), .ZN(n907) );
  NAND2_X1 U1005 ( .A1(G130), .A2(n905), .ZN(n906) );
  NAND2_X1 U1006 ( .A1(n907), .A2(n906), .ZN(n915) );
  NAND2_X1 U1007 ( .A1(n525), .A2(G142), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n909), .B(KEYINPUT114), .ZN(n912) );
  NAND2_X1 U1009 ( .A1(G106), .A2(n910), .ZN(n911) );
  NAND2_X1 U1010 ( .A1(n912), .A2(n911), .ZN(n913) );
  XOR2_X1 U1011 ( .A(n913), .B(KEYINPUT45), .Z(n914) );
  NOR2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1013 ( .A(n917), .B(n916), .Z(n919) );
  XNOR2_X1 U1014 ( .A(n919), .B(n918), .ZN(n920) );
  XNOR2_X1 U1015 ( .A(n920), .B(n1017), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n921), .ZN(G395) );
  NOR2_X1 U1017 ( .A1(G227), .A2(G229), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(KEYINPUT49), .B(n922), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(G397), .A2(n923), .ZN(n928) );
  NOR2_X1 U1020 ( .A1(n924), .A2(G401), .ZN(n925) );
  XOR2_X1 U1021 ( .A(KEYINPUT118), .B(n925), .Z(n926) );
  NOR2_X1 U1022 ( .A1(G395), .A2(n926), .ZN(n927) );
  NAND2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1026 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n1037) );
  INV_X1 U1027 ( .A(KEYINPUT55), .ZN(n1031) );
  XNOR2_X1 U1028 ( .A(KEYINPUT54), .B(G34), .ZN(n929) );
  XNOR2_X1 U1029 ( .A(n929), .B(KEYINPUT121), .ZN(n930) );
  XNOR2_X1 U1030 ( .A(G2084), .B(n930), .ZN(n946) );
  XNOR2_X1 U1031 ( .A(G2090), .B(G35), .ZN(n944) );
  XOR2_X1 U1032 ( .A(G1991), .B(G25), .Z(n931) );
  NAND2_X1 U1033 ( .A1(n931), .A2(G28), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(G2067), .B(G26), .ZN(n933) );
  XNOR2_X1 U1035 ( .A(G33), .B(G2072), .ZN(n932) );
  NOR2_X1 U1036 ( .A1(n933), .A2(n932), .ZN(n939) );
  XOR2_X1 U1037 ( .A(n934), .B(G32), .Z(n937) );
  XOR2_X1 U1038 ( .A(n935), .B(G27), .Z(n936) );
  NOR2_X1 U1039 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1041 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1042 ( .A(KEYINPUT53), .B(n942), .ZN(n943) );
  NOR2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1045 ( .A(n1031), .B(n947), .ZN(n949) );
  INV_X1 U1046 ( .A(G29), .ZN(n948) );
  NAND2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(G11), .A2(n950), .ZN(n1005) );
  XNOR2_X1 U1049 ( .A(G16), .B(KEYINPUT56), .ZN(n977) );
  XNOR2_X1 U1050 ( .A(G1956), .B(n951), .ZN(n953) );
  NAND2_X1 U1051 ( .A1(G1971), .A2(G303), .ZN(n952) );
  NAND2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n958) );
  XOR2_X1 U1053 ( .A(G1341), .B(n954), .Z(n955) );
  NAND2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n967) );
  XOR2_X1 U1057 ( .A(G1966), .B(G168), .Z(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1059 ( .A(KEYINPUT123), .B(n963), .Z(n965) );
  XNOR2_X1 U1060 ( .A(KEYINPUT122), .B(KEYINPUT57), .ZN(n964) );
  XNOR2_X1 U1061 ( .A(n965), .B(n964), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n975) );
  XOR2_X1 U1063 ( .A(G1348), .B(n968), .Z(n970) );
  XOR2_X1 U1064 ( .A(G171), .B(G1961), .Z(n969) );
  NOR2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1066 ( .A(KEYINPUT124), .B(n971), .Z(n972) );
  NOR2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n1003) );
  INV_X1 U1070 ( .A(G16), .ZN(n1001) );
  XNOR2_X1 U1071 ( .A(G1986), .B(G24), .ZN(n982) );
  XNOR2_X1 U1072 ( .A(G1976), .B(G23), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(G22), .B(G1971), .ZN(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(KEYINPUT125), .B(n980), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(KEYINPUT58), .B(n983), .ZN(n985) );
  XOR2_X1 U1078 ( .A(G1961), .B(G5), .Z(n984) );
  NAND2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n998) );
  XOR2_X1 U1080 ( .A(G1966), .B(G21), .Z(n996) );
  XNOR2_X1 U1081 ( .A(G20), .B(n986), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(G1981), .B(G6), .ZN(n988) );
  XNOR2_X1 U1083 ( .A(G19), .B(G1341), .ZN(n987) );
  NOR2_X1 U1084 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1085 ( .A1(n990), .A2(n989), .ZN(n993) );
  XOR2_X1 U1086 ( .A(KEYINPUT59), .B(G1348), .Z(n991) );
  XNOR2_X1 U1087 ( .A(G4), .B(n991), .ZN(n992) );
  NOR2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1089 ( .A(n994), .B(KEYINPUT60), .ZN(n995) );
  NAND2_X1 U1090 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1092 ( .A(KEYINPUT61), .B(n999), .ZN(n1000) );
  NAND2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1035) );
  XOR2_X1 U1096 ( .A(G2072), .B(n1006), .Z(n1008) );
  XOR2_X1 U1097 ( .A(G164), .B(G2078), .Z(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(KEYINPUT50), .B(n1009), .ZN(n1015) );
  XOR2_X1 U1100 ( .A(G2090), .B(G162), .Z(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1102 ( .A(KEYINPUT51), .B(n1012), .Z(n1013) );
  XNOR2_X1 U1103 ( .A(KEYINPUT120), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1029) );
  INV_X1 U1105 ( .A(n1016), .ZN(n1022) );
  XNOR2_X1 U1106 ( .A(G160), .B(G2084), .ZN(n1018) );
  NAND2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  NOR2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1111 ( .A(KEYINPUT119), .B(n1025), .Z(n1026) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1114 ( .A(KEYINPUT52), .B(n1030), .ZN(n1032) );
  NAND2_X1 U1115 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1116 ( .A1(n1033), .A2(G29), .ZN(n1034) );
  NAND2_X1 U1117 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1118 ( .A(n1037), .B(n1036), .ZN(G311) );
  XNOR2_X1 U1119 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

