//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(KEYINPUT28), .A3(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G183gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT27), .B1(KEYINPUT66), .B2(G183gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND4_X1  g007(.A1(new_n205), .A2(KEYINPUT66), .A3(KEYINPUT27), .A4(G183gat), .ZN(new_n209));
  AOI21_X1  g008(.A(G190gat), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n211));
  OAI21_X1  g010(.A(new_n204), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT69), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT69), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n215), .B(new_n204), .C1(new_n210), .C2(new_n211), .ZN(new_n216));
  OR3_X1    g015(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n213), .A2(new_n214), .A3(new_n216), .A4(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(KEYINPUT64), .B(G176gat), .Z(new_n222));
  INV_X1    g021(.A(G169gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(KEYINPUT23), .A3(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n214), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n226), .B(new_n227), .C1(G183gat), .C2(G190gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT23), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(G169gat), .B2(G176gat), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n224), .A2(new_n218), .A3(new_n228), .A4(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT25), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G176gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n223), .A2(new_n234), .A3(KEYINPUT23), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n235), .A2(new_n236), .A3(new_n218), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n236), .B1(new_n235), .B2(new_n218), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT66), .B(G183gat), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n226), .B(new_n227), .C1(new_n240), .C2(G190gat), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n239), .A2(new_n241), .A3(KEYINPUT25), .A4(new_n230), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n233), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n221), .A2(new_n243), .ZN(new_n244));
  OR2_X1    g043(.A1(G127gat), .A2(G134gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n246));
  NAND2_X1  g045(.A1(G127gat), .A2(G134gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  AND2_X1   g047(.A1(G127gat), .A2(G134gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(G127gat), .A2(G134gat), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT70), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G120gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(KEYINPUT1), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT71), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n256));
  INV_X1    g055(.A(G113gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n257), .A2(G120gat), .ZN(new_n258));
  INV_X1    g057(.A(G120gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n259), .A2(G113gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n256), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n261), .A2(new_n262), .A3(new_n251), .A4(new_n248), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n255), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT72), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n253), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT72), .B1(new_n258), .B2(new_n260), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n245), .A2(new_n247), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n266), .A2(new_n267), .A3(new_n256), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n244), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n221), .A2(new_n243), .A3(new_n264), .A4(new_n269), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G227gat), .A2(G233gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n276), .A2(KEYINPUT73), .A3(KEYINPUT32), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT33), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n274), .B1(new_n271), .B2(new_n272), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT32), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(G15gat), .B(G43gat), .Z(new_n284));
  XNOR2_X1  g083(.A(G71gat), .B(G99gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n277), .A2(new_n279), .A3(new_n283), .A4(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT74), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n278), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(new_n288), .B2(new_n286), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n276), .A2(KEYINPUT32), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT34), .B1(new_n275), .B2(KEYINPUT75), .ZN(new_n293));
  INV_X1    g092(.A(new_n273), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n293), .B1(new_n294), .B2(new_n274), .ZN(new_n295));
  INV_X1    g094(.A(new_n293), .ZN(new_n296));
  NOR3_X1   g095(.A1(new_n273), .A2(new_n275), .A3(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n292), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n287), .A2(new_n291), .A3(new_n298), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT31), .B(G50gat), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G228gat), .ZN(new_n305));
  INV_X1    g104(.A(G233gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT76), .B(G211gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT77), .B(G218gat), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT22), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(G197gat), .B(G204gat), .Z(new_n311));
  XOR2_X1   g110(.A(G211gat), .B(G218gat), .Z(new_n312));
  OR3_X1    g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n312), .B1(new_n310), .B2(new_n311), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G148gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G141gat), .ZN(new_n318));
  INV_X1    g117(.A(G141gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G148gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT80), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT2), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n318), .A2(new_n320), .A3(KEYINPUT80), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n324), .ZN(new_n328));
  NOR2_X1   g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT81), .B(G141gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n318), .B1(new_n333), .B2(new_n317), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT82), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(new_n328), .B2(new_n329), .ZN(new_n336));
  INV_X1    g135(.A(new_n329), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(KEYINPUT82), .A3(new_n324), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n334), .A2(new_n325), .A3(new_n336), .A4(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n331), .A2(new_n332), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n316), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT87), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n316), .A2(new_n342), .A3(KEYINPUT87), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n330), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n318), .A2(new_n320), .A3(KEYINPUT80), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT80), .B1(new_n318), .B2(new_n320), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n348), .B1(new_n351), .B2(new_n325), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n319), .A2(KEYINPUT81), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT81), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G141gat), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n317), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n318), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n325), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n338), .A2(new_n336), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n352), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT29), .B1(new_n313), .B2(new_n314), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT86), .ZN(new_n363));
  OR2_X1    g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT3), .B1(new_n362), .B2(new_n363), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n361), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n307), .B1(new_n347), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G78gat), .B(G106gat), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n368), .B(G22gat), .Z(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n331), .A2(new_n339), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n371), .B1(new_n362), .B2(KEYINPUT3), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n372), .B(new_n343), .C1(new_n305), .C2(new_n306), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n367), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n370), .B1(new_n367), .B2(new_n373), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n304), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n367), .A2(new_n373), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n369), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n367), .A2(new_n370), .A3(new_n373), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(new_n303), .A3(new_n379), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n302), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n264), .A2(new_n269), .A3(new_n331), .A4(new_n339), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT3), .B1(new_n352), .B2(new_n360), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(new_n270), .A3(new_n340), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n361), .A2(KEYINPUT4), .A3(new_n264), .A4(new_n269), .ZN(new_n388));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n385), .A2(new_n387), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n270), .A2(new_n371), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n383), .ZN(new_n392));
  INV_X1    g191(.A(new_n389), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  XOR2_X1   g193(.A(KEYINPUT83), .B(KEYINPUT5), .Z(new_n395));
  NAND3_X1  g194(.A1(new_n390), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  AND4_X1   g195(.A1(new_n389), .A2(new_n385), .A3(new_n387), .A4(new_n388), .ZN(new_n397));
  INV_X1    g196(.A(new_n395), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT84), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT84), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n390), .A2(new_n400), .A3(new_n395), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n396), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G1gat), .B(G29gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(G85gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT0), .B(G57gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT6), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n406), .B(new_n396), .C1(new_n399), .C2(new_n401), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT85), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n402), .A2(KEYINPUT6), .A3(new_n407), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT85), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n408), .A2(new_n414), .A3(new_n409), .A4(new_n410), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n412), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n244), .A2(new_n341), .ZN(new_n417));
  NAND2_X1  g216(.A1(G226gat), .A2(G233gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(KEYINPUT78), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n244), .A2(new_n419), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n316), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n419), .B1(new_n244), .B2(new_n341), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT79), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n420), .B1(new_n221), .B2(new_n243), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT79), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n424), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n423), .B1(new_n429), .B2(new_n316), .ZN(new_n430));
  XNOR2_X1  g229(.A(G8gat), .B(G36gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(G64gat), .B(G92gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n424), .A2(new_n315), .A3(new_n427), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n427), .A2(KEYINPUT79), .ZN(new_n437));
  AOI211_X1 g236(.A(new_n425), .B(new_n420), .C1(new_n221), .C2(new_n243), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n421), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n436), .B1(new_n439), .B2(new_n315), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n433), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n435), .A2(new_n441), .A3(KEYINPUT30), .ZN(new_n442));
  OR3_X1    g241(.A1(new_n440), .A2(KEYINPUT30), .A3(new_n433), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n382), .A2(new_n416), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT35), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT90), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n411), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n408), .A2(KEYINPUT90), .A3(new_n409), .A4(new_n410), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n413), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n444), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT92), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n302), .A2(new_n381), .A3(KEYINPUT35), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n450), .A2(KEYINPUT92), .A3(new_n444), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n448), .A2(new_n449), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT91), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT38), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n459), .B(new_n433), .C1(new_n440), .C2(KEYINPUT37), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n429), .A2(new_n316), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n315), .B1(new_n424), .B2(new_n427), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(KEYINPUT37), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n458), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT37), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n434), .B1(new_n430), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n467), .A2(KEYINPUT91), .A3(new_n459), .A4(new_n463), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n435), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n430), .A2(new_n466), .ZN(new_n471));
  OAI211_X1 g270(.A(KEYINPUT37), .B(new_n423), .C1(new_n429), .C2(new_n316), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n433), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n470), .B1(new_n473), .B2(KEYINPUT38), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n457), .A2(new_n413), .A3(new_n469), .A4(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT39), .B1(new_n392), .B2(new_n393), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT88), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n385), .A2(new_n387), .A3(new_n388), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n393), .ZN(new_n480));
  OAI211_X1 g279(.A(KEYINPUT88), .B(KEYINPUT39), .C1(new_n392), .C2(new_n393), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT39), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n479), .A2(new_n483), .A3(new_n393), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(new_n484), .A3(new_n406), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT40), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n482), .A2(new_n484), .A3(KEYINPUT40), .A4(new_n406), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n408), .A3(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT89), .B1(new_n444), .B2(new_n489), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n487), .A2(new_n408), .A3(new_n488), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT89), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n443), .A4(new_n442), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n381), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n475), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT36), .ZN(new_n497));
  INV_X1    g296(.A(new_n301), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n298), .B1(new_n287), .B2(new_n291), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n300), .A2(KEYINPUT36), .A3(new_n301), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n416), .A2(new_n444), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n502), .B1(new_n503), .B2(new_n381), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n446), .A2(new_n456), .B1(new_n496), .B2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G43gat), .B(G50gat), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n506), .A2(KEYINPUT15), .ZN(new_n507));
  NOR3_X1   g306(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT94), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT95), .ZN(new_n513));
  INV_X1    g312(.A(G29gat), .ZN(new_n514));
  INV_X1    g313(.A(G36gat), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n507), .B(new_n509), .C1(new_n513), .C2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n516), .B1(new_n512), .B2(new_n509), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n506), .A2(KEYINPUT15), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n507), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT17), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT96), .ZN(new_n525));
  XOR2_X1   g324(.A(G15gat), .B(G22gat), .Z(new_n526));
  INV_X1    g325(.A(G1gat), .ZN(new_n527));
  OR3_X1    g326(.A1(new_n526), .A2(KEYINPUT97), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n527), .B1(new_n526), .B2(KEYINPUT97), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n528), .B(new_n529), .C1(KEYINPUT16), .C2(new_n526), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n530), .A2(G8gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(G8gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT98), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n517), .A2(KEYINPUT17), .A3(new_n521), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n533), .A2(KEYINPUT98), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n525), .A2(new_n534), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n533), .A2(new_n522), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(KEYINPUT18), .A3(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n533), .B(new_n522), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n540), .B(KEYINPUT13), .Z(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT18), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n541), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549));
  INV_X1    g348(.A(G197gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT11), .B(G169gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(KEYINPUT93), .Z(new_n554));
  XOR2_X1   g353(.A(new_n554), .B(KEYINPUT12), .Z(new_n555));
  NAND2_X1  g354(.A1(new_n548), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n555), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n541), .A2(new_n557), .A3(new_n544), .A4(new_n547), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G85gat), .A2(G92gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT7), .ZN(new_n562));
  INV_X1    g361(.A(G99gat), .ZN(new_n563));
  INV_X1    g362(.A(G106gat), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT8), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n562), .B(new_n565), .C1(G85gat), .C2(G92gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(G99gat), .B(G106gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G57gat), .B(G64gat), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G71gat), .B(G78gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n568), .B(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n568), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(new_n573), .ZN(new_n576));
  MUX2_X1   g375(.A(new_n574), .B(new_n576), .S(KEYINPUT10), .Z(new_n577));
  NAND2_X1  g376(.A1(G230gat), .A2(G233gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n579), .B1(new_n574), .B2(new_n578), .ZN(new_n580));
  XNOR2_X1  g379(.A(G176gat), .B(G204gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(new_n317), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT102), .B(G120gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n582), .B(new_n583), .Z(new_n584));
  XNOR2_X1  g383(.A(new_n580), .B(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n525), .A2(new_n535), .A3(new_n575), .ZN(new_n586));
  AND3_X1   g385(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n587), .B1(new_n522), .B2(new_n568), .ZN(new_n588));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n589), .B1(new_n586), .B2(new_n588), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G134gat), .B(G162gat), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n592), .A2(KEYINPUT100), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n586), .A2(new_n588), .ZN(new_n598));
  INV_X1    g397(.A(new_n589), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(KEYINPUT100), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(new_n595), .ZN(new_n603));
  AND3_X1   g402(.A1(new_n597), .A2(new_n603), .A3(KEYINPUT101), .ZN(new_n604));
  AOI22_X1  g403(.A1(new_n597), .A2(new_n603), .B1(KEYINPUT101), .B2(new_n592), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT21), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n531), .B(new_n532), .C1(new_n607), .C2(new_n573), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(G183gat), .ZN(new_n609));
  INV_X1    g408(.A(G231gat), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n609), .A2(new_n610), .A3(new_n306), .ZN(new_n611));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G127gat), .B(G155gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G211gat), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n616), .B1(new_n611), .B2(new_n613), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n573), .A2(new_n607), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT99), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n621), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n620), .B(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n606), .A2(new_n627), .ZN(new_n628));
  NOR4_X1   g427(.A1(new_n505), .A2(new_n560), .A3(new_n585), .A4(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n416), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(G1gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(G1324gat));
  INV_X1    g433(.A(new_n444), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n629), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n637));
  OR2_X1    g436(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n640), .A2(KEYINPUT42), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(KEYINPUT42), .ZN(new_n642));
  INV_X1    g441(.A(G8gat), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n641), .B(new_n642), .C1(new_n643), .C2(new_n636), .ZN(G1325gat));
  INV_X1    g443(.A(new_n302), .ZN(new_n645));
  AOI21_X1  g444(.A(G15gat), .B1(new_n629), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n502), .A2(G15gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT105), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n646), .B1(new_n629), .B2(new_n648), .ZN(G1326gat));
  NAND2_X1  g448(.A1(new_n629), .A2(new_n381), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT43), .B(G22gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1327gat));
  INV_X1    g451(.A(new_n502), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n503), .A2(new_n381), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n474), .A2(new_n413), .A3(new_n448), .A4(new_n449), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n465), .A2(new_n468), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n495), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n490), .A2(new_n493), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n653), .B(new_n654), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n450), .A2(KEYINPUT92), .A3(new_n444), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT92), .B1(new_n450), .B2(new_n444), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT35), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n382), .A2(new_n662), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n660), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n445), .A2(KEYINPUT35), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n659), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n606), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n585), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n559), .A2(new_n626), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n671), .A2(new_n514), .A3(new_n630), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT106), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT45), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT44), .B1(new_n505), .B2(new_n606), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT107), .B1(new_n604), .B2(new_n605), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n592), .A2(KEYINPUT101), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n596), .B1(new_n592), .B2(KEYINPUT100), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n602), .A2(new_n595), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT107), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n597), .A2(new_n603), .A3(KEYINPUT101), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n676), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n666), .ZN(new_n687));
  AOI211_X1 g486(.A(KEYINPUT108), .B(new_n670), .C1(new_n675), .C2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT108), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n456), .A2(new_n446), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n606), .B1(new_n690), .B2(new_n659), .ZN(new_n691));
  OAI22_X1  g490(.A1(new_n691), .A2(new_n684), .B1(new_n505), .B2(new_n685), .ZN(new_n692));
  INV_X1    g491(.A(new_n670), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n689), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n688), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(G29gat), .B1(new_n695), .B2(new_n416), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n674), .A2(new_n696), .ZN(G1328gat));
  OAI21_X1  g496(.A(G36gat), .B1(new_n695), .B2(new_n444), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n671), .A2(new_n515), .A3(new_n635), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(KEYINPUT46), .Z(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(G1329gat));
  INV_X1    g500(.A(G43gat), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n671), .A2(new_n702), .A3(new_n645), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n502), .B1(new_n688), .B2(new_n694), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n704), .B1(new_n705), .B2(G43gat), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n707));
  INV_X1    g506(.A(KEYINPUT47), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n692), .A2(new_n502), .A3(new_n693), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n708), .B1(new_n709), .B2(G43gat), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT110), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n710), .A2(new_n711), .A3(new_n703), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n711), .B1(new_n710), .B2(new_n703), .ZN(new_n713));
  OAI22_X1  g512(.A1(new_n706), .A2(new_n707), .B1(new_n712), .B2(new_n713), .ZN(G1330gat));
  INV_X1    g513(.A(KEYINPUT111), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n684), .B1(new_n666), .B2(new_n667), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n685), .B1(new_n690), .B2(new_n659), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n693), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT108), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n692), .A2(new_n689), .A3(new_n693), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n495), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(G50gat), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n715), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n671), .A2(new_n722), .A3(new_n381), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n381), .B1(new_n688), .B2(new_n694), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n725), .A2(KEYINPUT111), .A3(G50gat), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT48), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(G50gat), .B1(new_n718), .B2(new_n495), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n730), .A2(KEYINPUT48), .A3(new_n724), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(G1331gat));
  NOR4_X1   g531(.A1(new_n505), .A2(new_n559), .A3(new_n669), .A4(new_n628), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n630), .ZN(new_n734));
  XOR2_X1   g533(.A(KEYINPUT112), .B(G57gat), .Z(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1332gat));
  INV_X1    g535(.A(KEYINPUT49), .ZN(new_n737));
  INV_X1    g536(.A(G64gat), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n733), .B(new_n635), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT113), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n738), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1333gat));
  AOI21_X1  g541(.A(G71gat), .B1(new_n733), .B2(new_n645), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n502), .A2(G71gat), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n733), .B2(new_n744), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g545(.A1(new_n733), .A2(new_n381), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g547(.A1(new_n626), .A2(new_n556), .A3(new_n558), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT114), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n691), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT115), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n668), .A2(new_n751), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT115), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n756), .A2(new_n757), .A3(KEYINPUT51), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(KEYINPUT51), .B2(new_n756), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(new_n630), .A3(new_n585), .ZN(new_n761));
  INV_X1    g560(.A(G85gat), .ZN(new_n762));
  AOI22_X1  g561(.A1(new_n668), .A2(KEYINPUT44), .B1(new_n666), .B2(new_n686), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n763), .A2(new_n669), .A3(new_n751), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n416), .A2(new_n762), .ZN(new_n765));
  AOI22_X1  g564(.A1(new_n761), .A2(new_n762), .B1(new_n764), .B2(new_n765), .ZN(G1336gat));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n635), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT52), .B1(new_n767), .B2(G92gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n760), .A2(new_n585), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n444), .A2(G92gat), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n768), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n756), .A2(KEYINPUT116), .A3(KEYINPUT51), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n753), .B2(new_n754), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n669), .B1(new_n776), .B2(new_n759), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n777), .A2(new_n770), .B1(G92gat), .B2(new_n767), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n772), .B1(new_n778), .B2(new_n779), .ZN(G1337gat));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n502), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT117), .ZN(new_n782));
  XNOR2_X1  g581(.A(KEYINPUT118), .B(G99gat), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n645), .A2(new_n784), .ZN(new_n785));
  OAI22_X1  g584(.A1(new_n782), .A2(new_n784), .B1(new_n769), .B2(new_n785), .ZN(G1338gat));
  NOR2_X1   g585(.A1(new_n495), .A2(G106gat), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n760), .A2(new_n585), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n692), .A2(new_n585), .A3(new_n381), .A4(new_n752), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n564), .A2(KEYINPUT119), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n564), .A2(KEYINPUT119), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n788), .A2(new_n789), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n793), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n795), .B1(new_n777), .B2(new_n787), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n796), .B2(new_n789), .ZN(G1339gat));
  NOR3_X1   g596(.A1(new_n604), .A2(new_n605), .A3(KEYINPUT107), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n681), .B1(new_n680), .B2(new_n682), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n579), .A2(KEYINPUT54), .ZN(new_n800));
  INV_X1    g599(.A(new_n584), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n577), .A2(new_n578), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n803), .A2(KEYINPUT54), .A3(new_n579), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n802), .A2(new_n804), .A3(KEYINPUT55), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT55), .B1(new_n802), .B2(new_n804), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n580), .A2(new_n584), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n539), .A2(new_n540), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n542), .A2(new_n543), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n553), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n808), .A2(new_n558), .A3(new_n811), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n798), .A2(new_n799), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n559), .A2(new_n808), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n558), .A2(new_n811), .A3(new_n585), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n676), .A2(new_n683), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n626), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n628), .A2(new_n559), .A3(new_n585), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(new_n382), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n630), .A3(new_n444), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n822), .A2(KEYINPUT120), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(KEYINPUT120), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n823), .A2(new_n257), .A3(new_n559), .A4(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(G113gat), .B1(new_n822), .B2(new_n560), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(G1340gat));
  NAND4_X1  g626(.A1(new_n823), .A2(new_n259), .A3(new_n585), .A4(new_n824), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n821), .A2(new_n630), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n585), .A2(new_n444), .ZN(new_n830));
  OAI21_X1  g629(.A(G120gat), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n828), .A2(new_n831), .ZN(G1341gat));
  NOR2_X1   g631(.A1(new_n822), .A2(new_n626), .ZN(new_n833));
  XNOR2_X1  g632(.A(KEYINPUT121), .B(G127gat), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n833), .B(new_n834), .ZN(G1342gat));
  NAND4_X1  g634(.A1(new_n821), .A2(new_n630), .A3(new_n444), .A4(new_n667), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(G134gat), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(KEYINPUT56), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT56), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n836), .A2(new_n839), .A3(G134gat), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT122), .B1(new_n836), .B2(G134gat), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n836), .A2(KEYINPUT122), .A3(G134gat), .ZN(new_n842));
  OAI22_X1  g641(.A1(new_n838), .A2(new_n840), .B1(new_n841), .B2(new_n842), .ZN(G1343gat));
  INV_X1    g642(.A(KEYINPUT123), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n815), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n558), .A2(new_n811), .A3(KEYINPUT123), .A4(new_n585), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n814), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n606), .ZN(new_n848));
  INV_X1    g647(.A(new_n812), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n676), .A2(new_n683), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n818), .B1(new_n851), .B2(new_n626), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT57), .B1(new_n852), .B2(new_n495), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n820), .A2(new_n854), .A3(new_n381), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n502), .A2(new_n416), .A3(new_n635), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n853), .A2(new_n855), .A3(new_n559), .A4(new_n856), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n820), .A2(new_n381), .A3(new_n856), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n560), .A2(G141gat), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n857), .A2(new_n333), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT58), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(KEYINPUT58), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n862), .B1(new_n860), .B2(new_n863), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(G1344gat));
  NAND3_X1  g665(.A1(new_n858), .A2(new_n317), .A3(new_n585), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n798), .A2(new_n799), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n814), .A2(new_n815), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n850), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n818), .B1(new_n870), .B2(new_n626), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT57), .B1(new_n871), .B2(new_n495), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n667), .A2(new_n849), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n627), .B1(new_n848), .B2(new_n873), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n854), .B(new_n381), .C1(new_n874), .C2(new_n818), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n856), .A2(new_n585), .ZN(new_n877));
  OAI21_X1  g676(.A(G148gat), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n878), .A2(KEYINPUT59), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n669), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n881), .A2(KEYINPUT59), .A3(new_n317), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n867), .B1(new_n879), .B2(new_n882), .ZN(G1345gat));
  OAI21_X1  g682(.A(G155gat), .B1(new_n880), .B2(new_n626), .ZN(new_n884));
  INV_X1    g683(.A(G155gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n858), .A2(new_n885), .A3(new_n627), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(G1346gat));
  INV_X1    g686(.A(new_n868), .ZN(new_n888));
  OAI21_X1  g687(.A(G162gat), .B1(new_n880), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(G162gat), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n858), .A2(new_n890), .A3(new_n667), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(G1347gat));
  NAND2_X1  g691(.A1(new_n416), .A2(new_n635), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT126), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n821), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G169gat), .B1(new_n895), .B2(new_n560), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT125), .B1(new_n871), .B2(new_n630), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT125), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n820), .A2(new_n898), .A3(new_n416), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n444), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n382), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n559), .A2(new_n223), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n896), .B1(new_n901), .B2(new_n902), .ZN(G1348gat));
  NOR3_X1   g702(.A1(new_n895), .A2(new_n669), .A3(new_n222), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n900), .A2(new_n585), .A3(new_n382), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(new_n234), .ZN(G1349gat));
  OAI21_X1  g705(.A(new_n240), .B1(new_n895), .B2(new_n626), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n627), .A2(new_n202), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n901), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT60), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n911), .B(new_n907), .C1(new_n901), .C2(new_n908), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1350gat));
  NAND3_X1  g712(.A1(new_n821), .A2(new_n667), .A3(new_n894), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(new_n915), .A3(G190gat), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n915), .B1(new_n914), .B2(G190gat), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n868), .A2(new_n203), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n917), .A2(new_n918), .B1(new_n901), .B2(new_n919), .ZN(G1351gat));
  INV_X1    g719(.A(KEYINPUT127), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n876), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n872), .A2(KEYINPUT127), .A3(new_n875), .ZN(new_n923));
  AND4_X1   g722(.A1(G197gat), .A2(new_n922), .A3(new_n559), .A4(new_n923), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n894), .A2(new_n653), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n900), .A2(new_n559), .A3(new_n381), .A4(new_n653), .ZN(new_n926));
  AOI22_X1  g725(.A1(new_n924), .A2(new_n925), .B1(new_n550), .B2(new_n926), .ZN(G1352gat));
  AND3_X1   g726(.A1(new_n900), .A2(new_n381), .A3(new_n653), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT62), .ZN(new_n929));
  INV_X1    g728(.A(G204gat), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n928), .A2(new_n929), .A3(new_n930), .A4(new_n585), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n922), .A2(new_n585), .A3(new_n925), .A4(new_n923), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(G204gat), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n900), .A2(new_n930), .A3(new_n381), .A4(new_n653), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT62), .B1(new_n934), .B2(new_n669), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n931), .A2(new_n933), .A3(new_n935), .ZN(G1353gat));
  INV_X1    g735(.A(new_n308), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n928), .A2(new_n937), .A3(new_n627), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n872), .A2(new_n627), .A3(new_n875), .A4(new_n925), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT63), .B1(new_n939), .B2(G211gat), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n939), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G1354gat));
  AND4_X1   g741(.A1(new_n309), .A2(new_n922), .A3(new_n667), .A4(new_n923), .ZN(new_n943));
  INV_X1    g742(.A(G218gat), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n900), .A2(new_n381), .A3(new_n653), .A4(new_n868), .ZN(new_n945));
  AOI22_X1  g744(.A1(new_n943), .A2(new_n925), .B1(new_n944), .B2(new_n945), .ZN(G1355gat));
endmodule


