//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT74), .B(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT24), .B(G110), .ZN(new_n190));
  OR2_X1    g004(.A1(KEYINPUT68), .A2(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT68), .A2(G128), .ZN(new_n192));
  NAND4_X1  g006(.A1(new_n191), .A2(KEYINPUT75), .A3(G119), .A4(new_n192), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(G119), .A3(new_n192), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT75), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G119), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n190), .B(new_n193), .C1(new_n195), .C2(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT23), .B1(new_n197), .B2(G119), .ZN(new_n200));
  INV_X1    g014(.A(G119), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(G128), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(new_n194), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n199), .B1(new_n204), .B2(G110), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT16), .ZN(new_n206));
  INV_X1    g020(.A(G140), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(G125), .ZN(new_n209));
  INV_X1    g023(.A(G125), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G140), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  OAI211_X1 g026(.A(G146), .B(new_n208), .C1(new_n212), .C2(new_n206), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT76), .ZN(new_n214));
  XNOR2_X1  g028(.A(G125), .B(G140), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n215), .A2(new_n214), .A3(new_n216), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n205), .A2(new_n213), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n208), .B1(new_n212), .B2(new_n206), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n216), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n213), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n204), .A2(G110), .ZN(new_n225));
  MUX2_X1   g039(.A(new_n196), .B(new_n198), .S(new_n194), .Z(new_n226));
  OAI211_X1 g040(.A(new_n224), .B(new_n225), .C1(new_n226), .C2(new_n190), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT22), .B(G137), .ZN(new_n228));
  INV_X1    g042(.A(G953), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(G221), .A3(G234), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n228), .B(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n221), .A2(new_n227), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n231), .B1(new_n221), .B2(new_n227), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT25), .B1(new_n235), .B2(new_n188), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT25), .ZN(new_n237));
  INV_X1    g051(.A(new_n188), .ZN(new_n238));
  NOR4_X1   g052(.A1(new_n233), .A2(new_n234), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n189), .B1(new_n236), .B2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n189), .A2(G902), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n235), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT32), .ZN(new_n244));
  XOR2_X1   g058(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n245));
  INV_X1    g059(.A(G237), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(new_n229), .A3(G210), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n245), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G101), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT28), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT2), .B(G113), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n201), .A2(G116), .ZN(new_n255));
  INV_X1    g069(.A(G116), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G119), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n255), .A2(new_n257), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n253), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n259), .A2(KEYINPUT69), .A3(new_n261), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT65), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT11), .ZN(new_n268));
  INV_X1    g082(.A(G137), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n267), .A2(new_n268), .A3(new_n269), .A4(G134), .ZN(new_n270));
  INV_X1    g084(.A(G134), .ZN(new_n271));
  OAI22_X1  g085(.A1(new_n271), .A2(G137), .B1(KEYINPUT65), .B2(KEYINPUT11), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n274), .B1(new_n269), .B2(G134), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G131), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n273), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT66), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n275), .B1(new_n272), .B2(new_n270), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT66), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(new_n277), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n269), .A2(G134), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n271), .A2(G137), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT67), .ZN(new_n286));
  OAI21_X1  g100(.A(G131), .B1(new_n285), .B2(KEYINPUT67), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n216), .A2(G143), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT64), .ZN(new_n290));
  INV_X1    g104(.A(G143), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n290), .B1(new_n291), .B2(G146), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n216), .A2(KEYINPUT64), .A3(G143), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n289), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n191), .A2(new_n192), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n289), .A2(KEYINPUT1), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(G143), .B(G146), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT1), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n300), .A3(G128), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n288), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n283), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n280), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n279), .A2(new_n282), .B1(G131), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n306));
  XOR2_X1   g120(.A(KEYINPUT0), .B(G128), .Z(new_n307));
  NAND2_X1  g121(.A1(new_n291), .A2(G146), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n289), .A2(new_n308), .A3(G128), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n294), .A2(new_n307), .B1(new_n309), .B2(KEYINPUT0), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NOR3_X1   g125(.A1(new_n305), .A2(new_n306), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n304), .A2(G131), .ZN(new_n313));
  AND4_X1   g127(.A1(new_n281), .A2(new_n273), .A3(new_n277), .A4(new_n276), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n281), .B1(new_n280), .B2(new_n277), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT70), .B1(new_n316), .B2(new_n310), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n266), .B(new_n303), .C1(new_n312), .C2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n303), .B1(new_n305), .B2(new_n311), .ZN(new_n319));
  INV_X1    g133(.A(new_n266), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n252), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n252), .B1(new_n319), .B2(new_n320), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n251), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  OAI211_X1 g139(.A(KEYINPUT30), .B(new_n303), .C1(new_n312), .C2(new_n317), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT30), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n266), .B1(new_n319), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n283), .A2(new_n302), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n306), .B1(new_n305), .B2(new_n311), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n316), .A2(KEYINPUT70), .A3(new_n310), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n251), .B1(new_n333), .B2(new_n266), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT73), .B(KEYINPUT31), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n329), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n325), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n329), .A2(new_n334), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT72), .B1(new_n339), .B2(KEYINPUT31), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT72), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT31), .ZN(new_n342));
  AOI211_X1 g156(.A(new_n341), .B(new_n342), .C1(new_n329), .C2(new_n334), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n338), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(G472), .A2(G902), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n244), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n316), .A2(new_n310), .B1(new_n283), .B2(new_n302), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n320), .B1(new_n348), .B2(KEYINPUT30), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n349), .B1(KEYINPUT30), .B2(new_n333), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n318), .A2(new_n250), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT31), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n341), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n339), .A2(KEYINPUT72), .A3(KEYINPUT31), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n353), .A2(new_n325), .A3(new_n337), .A4(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n346), .A2(new_n244), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n333), .A2(new_n266), .ZN(new_n357));
  AOI211_X1 g171(.A(new_n320), .B(new_n330), .C1(new_n331), .C2(new_n332), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT28), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n323), .A2(new_n250), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT29), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n326), .A2(new_n328), .B1(new_n333), .B2(new_n266), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n361), .B1(new_n364), .B2(new_n250), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n322), .A2(new_n360), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n363), .B(new_n188), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  AOI22_X1  g181(.A1(new_n355), .A2(new_n356), .B1(new_n367), .B2(G472), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n243), .B1(new_n347), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT78), .ZN(new_n370));
  INV_X1    g184(.A(G104), .ZN(new_n371));
  AND2_X1   g185(.A1(KEYINPUT77), .A2(G107), .ZN(new_n372));
  NOR2_X1   g186(.A1(KEYINPUT77), .A2(G107), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n370), .B(new_n371), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G107), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G104), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT77), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n375), .ZN(new_n379));
  NAND2_X1  g193(.A1(KEYINPUT77), .A2(G107), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n370), .B1(new_n381), .B2(new_n371), .ZN(new_n382));
  OAI21_X1  g196(.A(G101), .B1(new_n377), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n197), .B1(new_n289), .B2(KEYINPUT1), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT79), .B1(new_n384), .B2(new_n299), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n289), .A2(new_n308), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT79), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n300), .B1(G143), .B2(new_n216), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n386), .B(new_n387), .C1(new_n197), .C2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n385), .A2(new_n389), .A3(new_n301), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT3), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n379), .A2(new_n391), .A3(G104), .A4(new_n380), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n391), .B1(new_n375), .B2(G104), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n376), .ZN(new_n394));
  INV_X1    g208(.A(G101), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n383), .A2(new_n390), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT10), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT64), .B1(new_n216), .B2(G143), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n290), .A2(new_n291), .A3(G146), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n400), .A2(new_n401), .B1(G143), .B2(new_n216), .ZN(new_n402));
  AOI22_X1  g216(.A1(new_n191), .A2(new_n192), .B1(new_n289), .B2(KEYINPUT1), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n301), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n383), .A2(KEYINPUT10), .A3(new_n404), .A4(new_n396), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n392), .A2(new_n394), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT4), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n407), .A3(G101), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n396), .A2(KEYINPUT4), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n395), .B1(new_n392), .B2(new_n394), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n310), .B(new_n408), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n399), .A2(new_n305), .A3(new_n405), .A4(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G110), .B(G140), .ZN(new_n413));
  INV_X1    g227(.A(G227), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(G953), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n413), .B(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT80), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n405), .A2(new_n411), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT78), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(new_n376), .A3(new_n374), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n421), .B1(new_n424), .B2(G101), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT10), .B1(new_n425), .B2(new_n390), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n316), .B1(new_n420), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT80), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n412), .A2(new_n428), .A3(new_n417), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n419), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n383), .A2(new_n390), .A3(new_n396), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n404), .B1(new_n383), .B2(new_n396), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n316), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT12), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(KEYINPUT12), .B(new_n316), .C1(new_n431), .C2(new_n432), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n437), .A2(new_n412), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n430), .B1(new_n438), .B2(new_n417), .ZN(new_n439));
  INV_X1    g253(.A(G902), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G469), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n418), .B1(new_n436), .B2(new_n435), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n417), .B1(new_n427), .B2(new_n412), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n442), .B(new_n188), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT81), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n420), .A2(new_n426), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n416), .B1(new_n447), .B2(new_n305), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n437), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n427), .A2(new_n412), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n416), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n238), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT81), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n453), .A3(new_n442), .ZN(new_n454));
  AOI22_X1  g268(.A1(G469), .A2(new_n441), .B1(new_n446), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(G214), .B1(G237), .B2(G902), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT82), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n298), .A2(new_n457), .A3(new_n210), .A4(new_n301), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n310), .A2(new_n210), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT82), .B1(new_n404), .B2(G125), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G224), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(G953), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n461), .B(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n258), .A2(KEYINPUT5), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n255), .A2(KEYINPUT5), .ZN(new_n467));
  INV_X1    g281(.A(G113), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n466), .A2(new_n469), .B1(new_n258), .B2(new_n254), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n383), .A2(new_n470), .A3(new_n396), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n471), .B1(new_n266), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(G110), .B(G122), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n471), .B(new_n474), .C1(new_n266), .C2(new_n472), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(KEYINPUT6), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT6), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n473), .A2(new_n479), .A3(new_n475), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n465), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n461), .A2(KEYINPUT7), .A3(new_n464), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n464), .A2(KEYINPUT7), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n458), .B(new_n483), .C1(new_n459), .C2(new_n460), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n477), .A2(new_n484), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n474), .B(KEYINPUT8), .Z(new_n486));
  NAND2_X1  g300(.A1(new_n383), .A2(new_n396), .ZN(new_n487));
  INV_X1    g301(.A(new_n470), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n486), .B1(new_n489), .B2(new_n471), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT83), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI211_X1 g306(.A(KEYINPUT83), .B(new_n486), .C1(new_n489), .C2(new_n471), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n482), .B(new_n485), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n481), .A2(new_n494), .A3(new_n440), .ZN(new_n495));
  OAI21_X1  g309(.A(G210), .B1(G237), .B2(G902), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n490), .B(new_n491), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n482), .A2(new_n477), .A3(new_n484), .ZN(new_n500));
  AOI21_X1  g314(.A(G902), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n496), .B1(new_n501), .B2(new_n481), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n456), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT84), .B(G143), .ZN(new_n504));
  INV_X1    g318(.A(G214), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n505), .A2(G237), .A3(G953), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n291), .A2(KEYINPUT84), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(G131), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT17), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT84), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n506), .B1(new_n512), .B2(G143), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n513), .B(new_n277), .C1(new_n506), .C2(new_n504), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n510), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(KEYINPUT17), .B(G131), .C1(new_n507), .C2(new_n509), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n515), .A2(new_n223), .A3(new_n213), .A4(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(KEYINPUT18), .B(G131), .C1(new_n507), .C2(new_n509), .ZN(new_n518));
  INV_X1    g332(.A(new_n507), .ZN(new_n519));
  NAND2_X1  g333(.A1(KEYINPUT18), .A2(G131), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n513), .A3(new_n520), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n218), .A2(new_n219), .ZN(new_n522));
  OR3_X1    g336(.A1(new_n215), .A2(KEYINPUT85), .A3(new_n216), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT85), .B1(new_n215), .B2(new_n216), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n518), .B(new_n521), .C1(new_n522), .C2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(G113), .B(G122), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(new_n371), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n517), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n510), .A2(new_n514), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n215), .B(KEYINPUT19), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n216), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(new_n213), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n528), .B1(new_n526), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(G475), .A2(G902), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT20), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT20), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n539), .B(new_n536), .C1(new_n529), .C2(new_n534), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n528), .B1(new_n517), .B2(new_n526), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n440), .B1(new_n529), .B2(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT86), .B(G475), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n538), .A2(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n191), .A2(G143), .A3(new_n192), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n197), .A2(G143), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT13), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n291), .A2(G128), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT13), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n545), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(G134), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n545), .A2(new_n271), .A3(new_n548), .ZN(new_n553));
  INV_X1    g367(.A(G122), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(G116), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n554), .A2(G116), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n381), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n256), .A2(G122), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n379), .A2(new_n555), .A3(new_n559), .A4(new_n380), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n552), .A2(new_n553), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT9), .B(G234), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n563), .A2(new_n187), .A3(G953), .ZN(new_n564));
  INV_X1    g378(.A(new_n553), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n271), .B1(new_n545), .B2(new_n548), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n560), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT14), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n568), .B1(new_n256), .B2(G122), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n559), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n570), .A2(KEYINPUT87), .B1(new_n568), .B2(new_n557), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT87), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n572), .A3(new_n559), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n375), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n562), .B(new_n564), .C1(new_n567), .C2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT88), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n562), .B1(new_n567), .B2(new_n574), .ZN(new_n578));
  INV_X1    g392(.A(new_n564), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT14), .B1(new_n554), .B2(G116), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT87), .B1(new_n581), .B2(new_n557), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n582), .B(new_n573), .C1(KEYINPUT14), .C2(new_n559), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G107), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n545), .A2(new_n548), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G134), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n553), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n584), .A2(new_n587), .A3(new_n560), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n588), .A2(KEYINPUT88), .A3(new_n562), .A4(new_n564), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n577), .A2(new_n580), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(G478), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(KEYINPUT15), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n590), .A2(new_n188), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n593), .B1(new_n590), .B2(new_n188), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(G952), .ZN(new_n598));
  AOI211_X1 g412(.A(G953), .B(new_n598), .C1(G234), .C2(G237), .ZN(new_n599));
  AOI211_X1 g413(.A(new_n229), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT21), .B(G898), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n544), .A2(new_n597), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(G221), .B1(new_n563), .B2(G902), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NOR4_X1   g420(.A1(new_n455), .A2(new_n503), .A3(new_n604), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n369), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G101), .ZN(G3));
  NAND2_X1  g423(.A1(new_n355), .A2(new_n345), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(G472), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n355), .B2(new_n188), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n455), .A2(new_n243), .A3(new_n606), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n590), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n564), .A2(KEYINPUT89), .ZN(new_n618));
  OR2_X1    g432(.A1(new_n578), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n578), .A2(new_n618), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(KEYINPUT33), .A3(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n617), .A2(G478), .A3(new_n188), .A4(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n590), .A2(new_n188), .ZN(new_n623));
  AOI21_X1  g437(.A(KEYINPUT90), .B1(new_n623), .B2(new_n591), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT90), .ZN(new_n625));
  AOI211_X1 g439(.A(new_n625), .B(G478), .C1(new_n590), .C2(new_n188), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n622), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT91), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g443(.A(KEYINPUT91), .B(new_n622), .C1(new_n624), .C2(new_n626), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n538), .A2(new_n540), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n542), .A2(new_n543), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n456), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n495), .A2(new_n497), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n501), .A2(new_n496), .A3(new_n481), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n603), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n614), .A2(new_n615), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  AOI21_X1  g458(.A(KEYINPUT92), .B1(new_n542), .B2(new_n543), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n542), .A2(KEYINPUT92), .A3(new_n543), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n632), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n596), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n594), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n640), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n614), .A2(new_n615), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NAND2_X1  g469(.A1(new_n221), .A2(new_n227), .ZN(new_n656));
  INV_X1    g470(.A(new_n231), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(KEYINPUT36), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n656), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n241), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n240), .A2(new_n660), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n661), .B(new_n456), .C1(new_n502), .C2(new_n498), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n455), .A2(new_n662), .A3(new_n606), .ZN(new_n663));
  INV_X1    g477(.A(new_n604), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n614), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT37), .B(G110), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  NAND2_X1  g481(.A1(new_n347), .A2(new_n368), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT93), .B(G900), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n600), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n599), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n651), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n663), .A2(new_n668), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G128), .ZN(G30));
  NAND2_X1  g490(.A1(new_n637), .A2(new_n638), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT38), .Z(new_n678));
  NAND3_X1  g492(.A1(new_n634), .A2(new_n650), .A3(new_n456), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n678), .A2(new_n661), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n446), .A2(new_n454), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n417), .B1(new_n437), .B2(new_n412), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n429), .A2(new_n427), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n682), .B1(new_n419), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(G469), .B1(new_n684), .B2(G902), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n606), .B1(new_n681), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n672), .B(KEYINPUT39), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n680), .B1(new_n688), .B2(KEYINPUT40), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(KEYINPUT40), .B2(new_n688), .ZN(new_n690));
  AOI22_X1  g504(.A1(new_n610), .A2(new_n244), .B1(new_n355), .B2(new_n356), .ZN(new_n691));
  OR3_X1    g505(.A1(new_n357), .A2(new_n358), .A3(new_n250), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n250), .B1(new_n350), .B2(new_n358), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n692), .A2(new_n693), .A3(KEYINPUT94), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n440), .ZN(new_n695));
  AOI21_X1  g509(.A(KEYINPUT94), .B1(new_n692), .B2(new_n693), .ZN(new_n696));
  OAI21_X1  g510(.A(G472), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT95), .B1(new_n691), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n355), .A2(new_n356), .ZN(new_n699));
  AND4_X1   g513(.A1(KEYINPUT95), .A2(new_n347), .A3(new_n699), .A4(new_n697), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n690), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G143), .ZN(G45));
  AOI211_X1 g516(.A(new_n673), .B(new_n544), .C1(new_n629), .C2(new_n630), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n663), .A2(new_n668), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G146), .ZN(G48));
  INV_X1    g519(.A(new_n243), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n367), .A2(G472), .ZN(new_n707));
  INV_X1    g521(.A(new_n356), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n707), .B1(new_n344), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(KEYINPUT32), .B1(new_n355), .B2(new_n345), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n706), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT96), .ZN(new_n712));
  AOI22_X1  g526(.A1(new_n437), .A2(new_n448), .B1(new_n450), .B2(new_n416), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n712), .B1(new_n713), .B2(new_n238), .ZN(new_n714));
  OAI211_X1 g528(.A(KEYINPUT96), .B(new_n188), .C1(new_n443), .C2(new_n444), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(G469), .A3(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n445), .A2(KEYINPUT81), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n453), .B1(new_n452), .B2(new_n442), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n716), .B(new_n605), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT97), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n681), .A2(KEYINPUT97), .A3(new_n605), .A4(new_n716), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n544), .B1(new_n629), .B2(new_n630), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n603), .A3(new_n639), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n711), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT41), .B(G113), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  NAND4_X1  g542(.A1(new_n369), .A2(new_n652), .A3(new_n721), .A4(new_n722), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  NAND2_X1  g544(.A1(new_n664), .A2(new_n661), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n347), .B2(new_n368), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(new_n639), .A3(new_n721), .A4(new_n722), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G119), .ZN(G21));
  AND2_X1   g548(.A1(new_n352), .A2(new_n337), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n359), .A2(new_n323), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n251), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n346), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n613), .A2(new_n243), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n634), .A2(new_n650), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n640), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n739), .A2(new_n721), .A3(new_n722), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  NAND3_X1  g557(.A1(new_n721), .A2(new_n639), .A3(new_n722), .ZN(new_n744));
  OAI21_X1  g558(.A(G472), .B1(new_n344), .B2(new_n238), .ZN(new_n745));
  INV_X1    g559(.A(new_n738), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n745), .A2(new_n703), .A3(new_n661), .A4(new_n746), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G125), .ZN(G27));
  NAND2_X1  g563(.A1(new_n711), .A2(KEYINPUT99), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT99), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n668), .A2(new_n751), .A3(new_n706), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT98), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n637), .A2(new_n638), .A3(new_n753), .A4(new_n456), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT98), .B1(new_n677), .B2(new_n636), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n686), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n703), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n750), .A2(new_n752), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT42), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n711), .A2(new_n756), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT42), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n762), .A3(new_n703), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G131), .ZN(G33));
  INV_X1    g579(.A(new_n674), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n711), .A2(new_n766), .A3(new_n756), .ZN(new_n767));
  XOR2_X1   g581(.A(KEYINPUT100), .B(G134), .Z(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(G36));
  NOR2_X1   g583(.A1(new_n442), .A2(new_n440), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n684), .A2(KEYINPUT45), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT102), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n442), .B1(new_n439), .B2(new_n773), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(KEYINPUT101), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(KEYINPUT101), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n772), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n777), .A2(KEYINPUT103), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(KEYINPUT103), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n770), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n780), .A2(KEYINPUT46), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n681), .B1(new_n780), .B2(KEYINPUT46), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n605), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n687), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n634), .B1(new_n629), .B2(new_n630), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT104), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT43), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(KEYINPUT43), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n785), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(new_n785), .B2(new_n789), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n614), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n792), .A2(KEYINPUT44), .A3(new_n793), .A4(new_n661), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT44), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n661), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n795), .B1(new_n796), .B2(new_n791), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n755), .A2(new_n754), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT105), .Z(new_n799));
  NAND3_X1  g613(.A1(new_n794), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  OR3_X1    g614(.A1(new_n783), .A2(new_n784), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G137), .ZN(G39));
  OR2_X1    g616(.A1(new_n781), .A2(new_n782), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(KEYINPUT47), .A3(new_n605), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT47), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n783), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NOR4_X1   g621(.A1(new_n668), .A2(new_n757), .A3(new_n798), .A4(new_n706), .ZN(new_n808));
  XOR2_X1   g622(.A(new_n808), .B(KEYINPUT106), .Z(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G140), .ZN(G42));
  NAND4_X1  g625(.A1(new_n785), .A2(new_n706), .A3(new_n605), .A4(new_n456), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(KEYINPUT107), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n681), .A2(new_n716), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT49), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n678), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n813), .B(new_n816), .C1(new_n815), .C2(new_n814), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n698), .A2(new_n700), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n812), .A2(KEYINPUT107), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n723), .A2(new_n798), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n821), .A2(new_n671), .A3(new_n791), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n822), .A2(new_n745), .A3(new_n661), .A4(new_n746), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n821), .A2(new_n243), .A3(new_n671), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n818), .ZN(new_n825));
  OR3_X1    g639(.A1(new_n825), .A2(new_n634), .A3(new_n631), .ZN(new_n826));
  XNOR2_X1  g640(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n792), .A2(new_n599), .A3(new_n739), .ZN(new_n828));
  INV_X1    g642(.A(new_n723), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n636), .A3(new_n678), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n827), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n832));
  OR4_X1    g646(.A1(new_n832), .A2(new_n828), .A3(KEYINPUT50), .A4(new_n830), .ZN(new_n833));
  AND4_X1   g647(.A1(new_n823), .A2(new_n826), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n814), .A2(new_n606), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n804), .A2(new_n806), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n828), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n839), .A2(new_n799), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n840), .B1(new_n836), .B2(new_n837), .ZN(new_n841));
  OAI211_X1 g655(.A(KEYINPUT51), .B(new_n834), .C1(new_n838), .C2(new_n841), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n835), .B(KEYINPUT113), .Z(new_n843));
  OAI21_X1  g657(.A(new_n840), .B1(new_n807), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n834), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT51), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n822), .A2(new_n750), .A3(new_n752), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n848), .B(KEYINPUT48), .Z(new_n849));
  NOR2_X1   g663(.A1(new_n825), .A2(new_n635), .ZN(new_n850));
  OAI211_X1 g664(.A(G952), .B(new_n229), .C1(new_n828), .C2(new_n744), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n842), .A2(new_n847), .A3(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n729), .A2(new_n733), .A3(new_n742), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n745), .A2(new_n686), .A3(new_n610), .A4(new_n706), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n544), .A2(new_n650), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT109), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n603), .A3(new_n639), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n745), .A2(new_n610), .A3(new_n664), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n686), .A2(new_n639), .A3(new_n661), .ZN(new_n860));
  OAI22_X1  g674(.A1(new_n855), .A2(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n726), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n608), .A2(new_n642), .A3(KEYINPUT108), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n608), .A2(new_n642), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT108), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n854), .A2(new_n862), .A3(new_n863), .A4(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT110), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n597), .A2(new_n672), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n869), .B1(new_n647), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n650), .A2(new_n673), .ZN(new_n872));
  INV_X1    g686(.A(new_n645), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n542), .A2(KEYINPUT92), .A3(new_n543), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n872), .A2(new_n875), .A3(KEYINPUT110), .A4(new_n632), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n871), .A2(new_n876), .A3(new_n661), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n877), .B1(new_n709), .B2(new_n710), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n756), .B1(new_n878), .B2(new_n747), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n767), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n760), .A2(new_n880), .A3(new_n763), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT52), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n663), .B(new_n668), .C1(new_n674), .C2(new_n703), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n883), .B1(new_n744), .B2(new_n747), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n740), .A2(new_n661), .A3(new_n673), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n686), .A2(new_n885), .A3(new_n639), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n347), .A2(new_n699), .A3(new_n697), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT95), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n691), .A2(KEYINPUT95), .A3(new_n697), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n882), .B1(new_n884), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n886), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(new_n698), .B2(new_n700), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n894), .A2(KEYINPUT52), .A3(new_n748), .A4(new_n883), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n868), .A2(new_n881), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT53), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n760), .A2(new_n880), .A3(new_n763), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n867), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g715(.A(KEYINPUT111), .B(new_n882), .C1(new_n884), .C2(new_n891), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT111), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n892), .A2(new_n895), .A3(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n901), .A2(KEYINPUT53), .A3(new_n902), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n899), .A2(new_n905), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n906), .A2(KEYINPUT54), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n901), .A2(KEYINPUT53), .A3(new_n896), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n904), .A2(new_n902), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n909), .A2(new_n867), .A3(new_n900), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n910), .B2(KEYINPUT53), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT54), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n907), .A2(new_n912), .A3(KEYINPUT112), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n912), .A2(KEYINPUT112), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n853), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(G952), .A2(G953), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n820), .B1(new_n915), .B2(new_n916), .ZN(G75));
  NOR2_X1   g731(.A1(new_n229), .A2(G952), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT117), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n188), .B1(new_n899), .B2(new_n905), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT56), .B1(new_n921), .B2(new_n497), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n478), .A2(new_n480), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(new_n465), .Z(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT55), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  OR3_X1    g741(.A1(new_n922), .A2(KEYINPUT116), .A3(new_n926), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT116), .B1(new_n922), .B2(new_n926), .ZN(new_n929));
  AOI211_X1 g743(.A(new_n920), .B(new_n927), .C1(new_n928), .C2(new_n929), .ZN(G51));
  INV_X1    g744(.A(KEYINPUT118), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n906), .A2(KEYINPUT54), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n907), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n906), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n770), .B(KEYINPUT57), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n443), .B2(new_n444), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n921), .A2(new_n778), .A3(new_n779), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT119), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n918), .B1(new_n937), .B2(new_n939), .ZN(G54));
  NAND3_X1  g754(.A1(new_n921), .A2(KEYINPUT58), .A3(G475), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n941), .A2(new_n535), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n941), .A2(new_n535), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n942), .A2(new_n943), .A3(new_n918), .ZN(G60));
  NAND2_X1  g758(.A1(new_n617), .A2(new_n621), .ZN(new_n945));
  NAND2_X1  g759(.A1(G478), .A2(G902), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT59), .Z(new_n947));
  NOR2_X1   g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n933), .A2(new_n934), .A3(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n947), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n914), .A2(new_n913), .A3(new_n950), .ZN(new_n951));
  AOI211_X1 g765(.A(new_n920), .B(new_n949), .C1(new_n951), .C2(new_n945), .ZN(G63));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n953));
  XNOR2_X1  g767(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n187), .A2(new_n440), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n829), .A2(new_n369), .A3(new_n641), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n503), .A2(new_n602), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n614), .A2(new_n615), .A3(new_n958), .A4(new_n857), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n957), .A2(new_n665), .A3(new_n959), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n608), .A2(new_n642), .A3(KEYINPUT108), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT108), .B1(new_n608), .B2(new_n642), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n881), .A2(new_n963), .A3(KEYINPUT53), .A4(new_n854), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n964), .A2(new_n909), .ZN(new_n965));
  AOI21_X1  g779(.A(KEYINPUT53), .B1(new_n901), .B2(new_n896), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n956), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n235), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n920), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n659), .B(new_n956), .C1(new_n965), .C2(new_n966), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT121), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n970), .A2(new_n971), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n953), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT123), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT122), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n967), .B2(new_n968), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n920), .A2(new_n953), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n970), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n967), .A2(new_n977), .A3(new_n968), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n976), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n956), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(new_n899), .B2(new_n905), .ZN(new_n985));
  OAI21_X1  g799(.A(KEYINPUT122), .B1(new_n985), .B2(new_n235), .ZN(new_n986));
  INV_X1    g800(.A(new_n979), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n987), .B1(new_n985), .B2(new_n659), .ZN(new_n988));
  AND4_X1   g802(.A1(new_n976), .A2(new_n986), .A3(new_n988), .A4(new_n982), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n975), .B1(new_n983), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(KEYINPUT124), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT124), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n992), .B(new_n975), .C1(new_n983), .C2(new_n989), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n991), .A2(new_n993), .ZN(G66));
  OAI21_X1  g808(.A(G953), .B1(new_n601), .B2(new_n462), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n868), .B2(G953), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n923), .B1(G898), .B2(new_n229), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(G69));
  OAI211_X1 g812(.A(new_n761), .B(new_n687), .C1(new_n724), .C2(new_n857), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT125), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n801), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT126), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n701), .A2(new_n748), .A3(new_n883), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT62), .Z(new_n1005));
  NAND3_X1  g819(.A1(new_n1003), .A2(new_n810), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n326), .B1(KEYINPUT30), .B2(new_n348), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(new_n531), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1006), .A2(new_n229), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n414), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n229), .B1(new_n1010), .B2(G900), .ZN(new_n1011));
  INV_X1    g825(.A(new_n810), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n750), .A2(new_n752), .ZN(new_n1013));
  AOI211_X1 g827(.A(new_n679), .B(new_n1013), .C1(new_n637), .C2(new_n638), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n803), .A2(new_n605), .A3(new_n687), .A4(new_n1014), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n884), .A2(new_n767), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n801), .A2(new_n1015), .A3(new_n764), .A4(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n229), .B1(new_n1012), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1008), .B1(new_n414), .B2(G953), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1011), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1009), .A2(new_n1020), .ZN(G72));
  NAND2_X1  g835(.A1(G472), .A2(G902), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT63), .Z(new_n1023));
  NOR2_X1   g837(.A1(new_n364), .A2(new_n250), .ZN(new_n1024));
  AND2_X1   g838(.A1(new_n1024), .A2(KEYINPUT127), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n339), .B1(new_n1024), .B2(KEYINPUT127), .ZN(new_n1026));
  OAI211_X1 g840(.A(new_n911), .B(new_n1023), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1023), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1028), .B1(new_n1029), .B2(new_n868), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n364), .A2(new_n251), .ZN(new_n1031));
  OAI221_X1 g845(.A(new_n1027), .B1(G952), .B2(new_n229), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g846(.A1(new_n1003), .A2(new_n810), .A3(new_n868), .A4(new_n1005), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n693), .B1(new_n1033), .B2(new_n1023), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n1032), .A2(new_n1034), .ZN(G57));
endmodule


