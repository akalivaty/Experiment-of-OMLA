//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070;
  OR2_X1    g000(.A1(KEYINPUT68), .A2(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT68), .A2(G119), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(G116), .A3(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  INV_X1    g005(.A(G113), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT2), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G113), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n189), .A2(new_n191), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT69), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n189), .A2(new_n196), .A3(KEYINPUT69), .A4(new_n191), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n189), .A2(new_n191), .ZN(new_n202));
  INV_X1    g016(.A(new_n196), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  NOR3_X1   g020(.A1(new_n206), .A2(KEYINPUT3), .A3(G107), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  AND2_X1   g022(.A1(KEYINPUT79), .A2(G104), .ZN(new_n209));
  NOR2_X1   g023(.A1(KEYINPUT79), .A2(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n207), .B1(new_n211), .B2(KEYINPUT3), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT79), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n206), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT79), .A2(G104), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(G107), .A3(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n205), .B1(new_n212), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n201), .A2(new_n204), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT4), .ZN(new_n220));
  INV_X1    g034(.A(new_n207), .ZN(new_n221));
  AOI21_X1  g035(.A(G107), .B1(new_n214), .B2(new_n215), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n221), .B(new_n216), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n220), .B1(new_n224), .B2(G101), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n209), .A2(new_n210), .ZN(new_n226));
  AOI21_X1  g040(.A(G101), .B1(new_n226), .B2(G107), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n212), .A2(KEYINPUT80), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT80), .B1(new_n212), .B2(new_n227), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n225), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n219), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n206), .A2(G107), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n205), .B1(new_n211), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT80), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n216), .A2(new_n205), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n212), .A2(KEYINPUT80), .A3(new_n227), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n233), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT5), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n187), .A2(new_n240), .A3(G116), .A4(new_n188), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n241), .B(KEYINPUT84), .ZN(new_n242));
  INV_X1    g056(.A(new_n191), .ZN(new_n243));
  AND2_X1   g057(.A1(KEYINPUT68), .A2(G119), .ZN(new_n244));
  NOR2_X1   g058(.A1(KEYINPUT68), .A2(G119), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n243), .B1(new_n246), .B2(G116), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n192), .B1(new_n247), .B2(KEYINPUT5), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n242), .A2(new_n248), .B1(new_n199), .B2(new_n200), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n239), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n231), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(G110), .B(G122), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n219), .A2(new_n230), .B1(new_n239), .B2(new_n249), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n252), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(KEYINPUT6), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G143), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT64), .B1(new_n258), .B2(G146), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT64), .ZN(new_n260));
  INV_X1    g074(.A(G146), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(G143), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n258), .A2(G146), .ZN(new_n263));
  INV_X1    g077(.A(G128), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(KEYINPUT1), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n259), .A2(new_n262), .A3(new_n263), .A4(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n261), .A2(G143), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n263), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n264), .B1(new_n267), .B2(KEYINPUT1), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OR2_X1    g085(.A1(new_n271), .A2(G125), .ZN(new_n272));
  NAND2_X1  g086(.A1(KEYINPUT0), .A2(G128), .ZN(new_n273));
  OR2_X1    g087(.A1(KEYINPUT0), .A2(G128), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n268), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n262), .A2(new_n263), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT65), .ZN(new_n278));
  INV_X1    g092(.A(new_n273), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n277), .A2(new_n278), .A3(new_n279), .A4(new_n259), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n259), .A2(new_n262), .A3(new_n279), .A4(new_n263), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT65), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n276), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G125), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n272), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G953), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G224), .ZN(new_n287));
  XOR2_X1   g101(.A(new_n285), .B(new_n287), .Z(new_n288));
  AOI21_X1  g102(.A(new_n252), .B1(new_n231), .B2(new_n250), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT6), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT85), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT85), .ZN(new_n292));
  NOR4_X1   g106(.A1(new_n255), .A2(new_n292), .A3(KEYINPUT6), .A4(new_n252), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n257), .B(new_n288), .C1(new_n291), .C2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n233), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n296), .B1(new_n228), .B2(new_n229), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n189), .A2(KEYINPUT5), .A3(new_n191), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n241), .A2(KEYINPUT84), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n241), .A2(KEYINPUT84), .ZN(new_n300));
  OAI211_X1 g114(.A(G113), .B(new_n298), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n201), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT86), .B1(new_n297), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT86), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n239), .A2(new_n304), .A3(new_n249), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n297), .A2(new_n302), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n252), .B(KEYINPUT8), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n287), .A2(KEYINPUT7), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n285), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n310), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n272), .B(new_n312), .C1(new_n283), .C2(new_n284), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n309), .A2(KEYINPUT87), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n256), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n314), .B1(new_n307), .B2(new_n308), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(KEYINPUT87), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n294), .B(new_n295), .C1(new_n317), .C2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(G210), .B1(G237), .B2(G902), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n321), .B(KEYINPUT88), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  OR2_X1    g137(.A1(new_n318), .A2(KEYINPUT87), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n318), .A2(KEYINPUT87), .B1(new_n252), .B2(new_n255), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n322), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n326), .A2(new_n295), .A3(new_n294), .A4(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT9), .B(G234), .ZN(new_n330));
  OAI21_X1  g144(.A(G221), .B1(new_n330), .B2(G902), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT77), .ZN(new_n332));
  INV_X1    g146(.A(G469), .ZN(new_n333));
  XOR2_X1   g147(.A(G110), .B(G140), .Z(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(KEYINPUT78), .ZN(new_n335));
  AND2_X1   g149(.A1(KEYINPUT70), .A2(G953), .ZN(new_n336));
  NOR2_X1   g150(.A1(KEYINPUT70), .A2(G953), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G227), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n335), .B(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n259), .A2(new_n262), .A3(new_n263), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n266), .B1(new_n344), .B2(new_n270), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n296), .B(new_n345), .C1(new_n228), .C2(new_n229), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT10), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n224), .A2(G101), .A3(new_n218), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n280), .A2(new_n282), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n349), .A2(new_n350), .A3(new_n275), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n230), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT11), .ZN(new_n353));
  INV_X1    g167(.A(G134), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n353), .B1(new_n354), .B2(G137), .ZN(new_n355));
  INV_X1    g169(.A(G137), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(KEYINPUT11), .A3(G134), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n354), .A2(G137), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n355), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G131), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT66), .B(G131), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n361), .A2(new_n355), .A3(new_n357), .A4(new_n358), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n271), .A2(KEYINPUT10), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n239), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n348), .A2(new_n352), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n351), .A2(new_n230), .B1(new_n239), .B2(new_n365), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n364), .B1(new_n369), .B2(new_n348), .ZN(new_n370));
  OAI211_X1 g184(.A(KEYINPUT83), .B(new_n343), .C1(new_n368), .C2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n346), .B1(new_n239), .B2(new_n271), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n364), .A2(KEYINPUT82), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT12), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT12), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n372), .A2(new_n376), .A3(new_n373), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n375), .A2(new_n342), .A3(new_n367), .A4(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n371), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n348), .A2(new_n352), .A3(new_n366), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n363), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n367), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT83), .B1(new_n382), .B2(new_n343), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n333), .B(new_n295), .C1(new_n379), .C2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n333), .A2(new_n295), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n375), .A2(new_n367), .A3(new_n377), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n367), .A2(new_n342), .ZN(new_n387));
  AOI22_X1  g201(.A1(new_n386), .A2(new_n343), .B1(new_n387), .B2(new_n381), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n385), .B1(new_n388), .B2(G469), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n332), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT16), .ZN(new_n391));
  INV_X1    g205(.A(G140), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(G125), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(G125), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n284), .A2(G140), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n393), .B1(new_n396), .B2(new_n391), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n261), .ZN(new_n398));
  OAI211_X1 g212(.A(G146), .B(new_n393), .C1(new_n396), .C2(new_n391), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  OR2_X1    g215(.A1(KEYINPUT70), .A2(G953), .ZN(new_n402));
  INV_X1    g216(.A(G237), .ZN(new_n403));
  NAND2_X1  g217(.A1(KEYINPUT70), .A2(G953), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n402), .A2(G214), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n258), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n338), .A2(G143), .A3(G214), .A4(new_n403), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n361), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT17), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n406), .A2(new_n407), .A3(new_n361), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n361), .B1(new_n406), .B2(new_n407), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT89), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n414), .A2(new_n415), .A3(KEYINPUT17), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n415), .B1(new_n414), .B2(KEYINPUT17), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n401), .B(new_n413), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G113), .B(G122), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(new_n206), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n408), .A2(KEYINPUT18), .A3(G131), .ZN(new_n421));
  NAND2_X1  g235(.A1(KEYINPUT18), .A2(G131), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n406), .A2(new_n407), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n396), .A2(G146), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n394), .A2(new_n395), .A3(new_n261), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n421), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n418), .A2(new_n420), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n420), .B1(new_n418), .B2(new_n427), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n295), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G475), .ZN(new_n432));
  INV_X1    g246(.A(new_n420), .ZN(new_n433));
  INV_X1    g247(.A(new_n427), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n396), .B(KEYINPUT19), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n399), .B1(new_n435), .B2(G146), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(new_n410), .B2(new_n412), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n433), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n428), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(G475), .A2(G902), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n440), .A2(KEYINPUT90), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(KEYINPUT90), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n439), .A2(KEYINPUT91), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n440), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n428), .B2(new_n438), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n446), .B1(new_n442), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n444), .B1(new_n428), .B2(new_n438), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(KEYINPUT91), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n432), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n286), .A2(G952), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(G234), .B2(G237), .ZN(new_n454));
  AOI211_X1 g268(.A(new_n295), .B(new_n338), .C1(G234), .C2(G237), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(G898), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G217), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n330), .A2(new_n458), .A3(G953), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT93), .ZN(new_n461));
  OR2_X1    g275(.A1(KEYINPUT92), .A2(G122), .ZN(new_n462));
  NAND2_X1  g276(.A1(KEYINPUT92), .A2(G122), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n190), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G122), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(G116), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n464), .A2(G107), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n463), .ZN(new_n468));
  NOR2_X1   g282(.A1(KEYINPUT92), .A2(G122), .ZN(new_n469));
  OAI21_X1  g283(.A(G116), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n466), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n208), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n461), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G107), .B1(new_n464), .B2(new_n466), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(new_n208), .A3(new_n471), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(KEYINPUT93), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n258), .A2(G128), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n264), .A2(G143), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n478), .A3(new_n354), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT13), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n481), .B1(new_n264), .B2(G143), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT94), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT94), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n477), .A2(new_n484), .A3(new_n481), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n264), .A2(G143), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT13), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n483), .A2(new_n485), .A3(new_n487), .A4(new_n478), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n480), .B1(new_n488), .B2(G134), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n473), .A2(new_n476), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT14), .B1(new_n465), .B2(G116), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT14), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n190), .A3(G122), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(G107), .B1(new_n464), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n258), .A2(G128), .ZN(new_n496));
  OAI21_X1  g310(.A(G134), .B1(new_n486), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n479), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n495), .A2(new_n475), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT95), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n495), .A2(KEYINPUT95), .A3(new_n498), .A4(new_n475), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n460), .B1(new_n490), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT96), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n473), .A2(new_n476), .A3(new_n489), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n506), .A2(new_n501), .A3(new_n502), .A4(new_n459), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n501), .A3(new_n502), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(KEYINPUT96), .A3(new_n460), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n295), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G478), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n512), .A2(KEYINPUT15), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n513), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n508), .A2(new_n295), .A3(new_n510), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NOR3_X1   g331(.A1(new_n452), .A2(new_n457), .A3(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(G214), .B1(G237), .B2(G902), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n329), .A2(new_n390), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n199), .A2(new_n200), .B1(new_n202), .B2(new_n203), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n281), .A2(KEYINPUT65), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n281), .A2(KEYINPUT65), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n363), .B(new_n275), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT30), .ZN(new_n526));
  INV_X1    g340(.A(G131), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n356), .A2(G134), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n527), .B1(new_n528), .B2(new_n358), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT67), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n530), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n271), .A2(new_n531), .A3(new_n362), .A4(new_n532), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n525), .A2(new_n526), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n526), .B1(new_n525), .B2(new_n533), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n522), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n525), .A2(new_n521), .A3(new_n533), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n338), .A2(G210), .A3(new_n403), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT27), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT26), .B(G101), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n540), .A2(new_n541), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT71), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n536), .A2(new_n537), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT31), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n536), .A2(KEYINPUT31), .A3(new_n537), .A4(new_n544), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n542), .A2(new_n543), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT28), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n537), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n537), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n521), .B1(new_n525), .B2(new_n533), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT28), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n550), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n549), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT32), .ZN(new_n560));
  NOR2_X1   g374(.A1(G472), .A2(G902), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n557), .B1(new_n547), .B2(new_n548), .ZN(new_n563));
  INV_X1    g377(.A(new_n561), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT32), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT29), .ZN(new_n567));
  INV_X1    g381(.A(new_n550), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n553), .B2(new_n556), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n536), .A2(new_n537), .A3(new_n568), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT72), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n556), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n568), .A2(new_n567), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n525), .A2(new_n533), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n522), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n537), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n552), .B1(new_n577), .B2(KEYINPUT28), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n573), .B(new_n574), .C1(new_n578), .C2(new_n572), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n571), .A2(new_n295), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G472), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n566), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G234), .ZN(new_n583));
  OAI21_X1  g397(.A(G217), .B1(new_n583), .B2(G902), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(KEYINPUT73), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT23), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n187), .A2(G128), .A3(new_n188), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n264), .A2(G119), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n187), .A2(new_n188), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT23), .B1(new_n590), .B2(new_n264), .ZN(new_n591));
  OAI21_X1  g405(.A(G110), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n587), .A2(new_n588), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(G110), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(KEYINPUT24), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT24), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G110), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n596), .A2(new_n598), .A3(KEYINPUT74), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT74), .B1(new_n596), .B2(new_n598), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT75), .B1(new_n594), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT75), .ZN(new_n603));
  NOR4_X1   g417(.A1(new_n593), .A2(new_n599), .A3(new_n600), .A4(new_n603), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n592), .B(new_n400), .C1(new_n602), .C2(new_n604), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n399), .A2(new_n425), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n589), .A2(new_n591), .A3(G110), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n594), .A2(new_n601), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n338), .A2(G221), .A3(G234), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT22), .B(G137), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n605), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n612), .B1(new_n605), .B2(new_n609), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(KEYINPUT25), .B1(new_n615), .B2(new_n295), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n605), .A2(new_n609), .ZN(new_n617));
  INV_X1    g431(.A(new_n612), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n605), .A2(new_n609), .A3(new_n612), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n619), .A2(KEYINPUT25), .A3(new_n295), .A4(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n585), .B1(new_n616), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT76), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n619), .A2(new_n295), .A3(new_n620), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT25), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n621), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n629), .A2(KEYINPUT76), .A3(new_n585), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n585), .A2(G902), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n615), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n625), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n582), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n520), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(new_n205), .ZN(G3));
  INV_X1    g451(.A(new_n519), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n323), .B2(new_n328), .ZN(new_n639));
  INV_X1    g453(.A(new_n457), .ZN(new_n640));
  INV_X1    g454(.A(G475), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n418), .A2(new_n427), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n433), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n428), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n641), .B1(new_n644), .B2(new_n295), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n439), .A2(new_n440), .ZN(new_n646));
  AOI22_X1  g460(.A1(new_n646), .A2(KEYINPUT20), .B1(new_n450), .B2(KEYINPUT91), .ZN(new_n647));
  INV_X1    g461(.A(new_n451), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT33), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n507), .A2(new_n505), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n462), .A2(new_n463), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n466), .B1(new_n652), .B2(G116), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n653), .A2(new_n208), .B1(new_n497), .B2(new_n479), .ZN(new_n654));
  AOI21_X1  g468(.A(KEYINPUT95), .B1(new_n654), .B2(new_n495), .ZN(new_n655));
  INV_X1    g469(.A(new_n502), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n459), .B1(new_n657), .B2(new_n506), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n510), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n650), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n509), .A2(KEYINPUT97), .A3(new_n460), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n507), .ZN(new_n663));
  AOI21_X1  g477(.A(KEYINPUT97), .B1(new_n509), .B2(new_n460), .ZN(new_n664));
  OAI21_X1  g478(.A(KEYINPUT33), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n512), .A2(G902), .ZN(new_n667));
  AOI22_X1  g481(.A1(new_n666), .A2(new_n667), .B1(new_n512), .B2(new_n511), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n649), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n639), .A2(new_n640), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT98), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT98), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n639), .A2(new_n672), .A3(new_n640), .A4(new_n669), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(G902), .B1(new_n549), .B2(new_n558), .ZN(new_n675));
  INV_X1    g489(.A(G472), .ZN(new_n676));
  OAI22_X1  g490(.A1(new_n675), .A2(new_n676), .B1(new_n564), .B2(new_n563), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n390), .A2(new_n678), .A3(new_n634), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT34), .B(G104), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G6));
  NOR2_X1   g497(.A1(new_n646), .A2(KEYINPUT20), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n448), .A2(new_n442), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n645), .A2(KEYINPUT99), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n645), .A2(KEYINPUT99), .ZN(new_n688));
  AND4_X1   g502(.A1(new_n517), .A2(new_n686), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n639), .A2(new_n689), .A3(new_n640), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n679), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n208), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT100), .B(KEYINPUT35), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G9));
  OAI21_X1  g508(.A(new_n617), .B1(KEYINPUT36), .B2(new_n618), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT36), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n605), .A2(new_n696), .A3(new_n609), .A4(new_n612), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n695), .A2(new_n631), .A3(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n698), .B(KEYINPUT101), .Z(new_n699));
  NAND3_X1  g513(.A1(new_n625), .A2(new_n630), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n625), .A2(new_n699), .A3(KEYINPUT102), .A4(new_n630), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n678), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n520), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT37), .B(G110), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G12));
  AOI22_X1  g522(.A1(new_n562), .A2(new_n565), .B1(G472), .B2(new_n580), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n709), .B1(new_n702), .B2(new_n703), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n687), .A2(new_n688), .ZN(new_n711));
  INV_X1    g525(.A(new_n517), .ZN(new_n712));
  INV_X1    g526(.A(G900), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n454), .B1(new_n455), .B2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n684), .B2(new_n685), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n711), .A2(new_n712), .A3(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n710), .A2(new_n717), .A3(new_n639), .A4(new_n390), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G128), .ZN(G30));
  XOR2_X1   g533(.A(new_n714), .B(KEYINPUT39), .Z(new_n720));
  AND2_X1   g534(.A1(new_n390), .A2(new_n720), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n721), .A2(KEYINPUT40), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(KEYINPUT40), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT104), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n722), .A2(new_n726), .A3(new_n723), .ZN(new_n727));
  AOI21_X1  g541(.A(KEYINPUT76), .B1(new_n629), .B2(new_n585), .ZN(new_n728));
  INV_X1    g542(.A(new_n585), .ZN(new_n729));
  AOI211_X1 g543(.A(new_n624), .B(new_n729), .C1(new_n628), .C2(new_n621), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT102), .B1(new_n731), .B2(new_n699), .ZN(new_n732));
  INV_X1    g546(.A(new_n703), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n536), .A2(new_n537), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n550), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n295), .B1(new_n577), .B2(new_n550), .ZN(new_n738));
  OAI21_X1  g552(.A(G472), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n566), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n452), .A2(new_n517), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n734), .A2(new_n519), .A3(new_n740), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n323), .A2(new_n328), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n744), .B1(new_n323), .B2(new_n328), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n725), .A2(new_n727), .A3(new_n748), .ZN(new_n749));
  XOR2_X1   g563(.A(KEYINPUT105), .B(G143), .Z(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G45));
  AND2_X1   g565(.A1(new_n662), .A2(new_n507), .ZN(new_n752));
  INV_X1    g566(.A(new_n664), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n650), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT33), .B1(new_n508), .B2(new_n510), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n667), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n511), .A2(new_n512), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n452), .A3(new_n715), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n710), .A2(new_n639), .A3(new_n390), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G146), .ZN(G48));
  OAI21_X1  g576(.A(new_n295), .B1(new_n379), .B2(new_n383), .ZN(new_n763));
  NAND2_X1  g577(.A1(KEYINPUT106), .A2(G469), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n332), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n295), .B(new_n764), .C1(new_n379), .C2(new_n383), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n633), .B1(new_n566), .B2(new_n581), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(new_n671), .B2(new_n673), .ZN(new_n772));
  XOR2_X1   g586(.A(KEYINPUT41), .B(G113), .Z(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(G15));
  AND3_X1   g588(.A1(new_n639), .A2(new_n689), .A3(new_n640), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n776), .A2(new_n709), .A3(new_n633), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G116), .ZN(G18));
  OAI211_X1 g593(.A(new_n582), .B(new_n518), .C1(new_n732), .C2(new_n733), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n329), .A2(new_n519), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n776), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G119), .ZN(G21));
  NAND2_X1  g599(.A1(new_n639), .A2(new_n742), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n573), .B1(new_n578), .B2(new_n572), .ZN(new_n788));
  AOI22_X1  g602(.A1(new_n788), .A2(new_n568), .B1(new_n547), .B2(new_n548), .ZN(new_n789));
  OAI22_X1  g603(.A1(new_n675), .A2(new_n676), .B1(new_n789), .B2(new_n564), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n790), .A2(new_n633), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n766), .A2(new_n767), .A3(new_n640), .A4(new_n768), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n787), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(KEYINPUT107), .B(G122), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(G24));
  AOI21_X1  g610(.A(new_n790), .B1(new_n702), .B2(new_n703), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(new_n639), .A3(new_n760), .A4(new_n769), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G125), .ZN(G27));
  NAND2_X1  g613(.A1(new_n384), .A2(new_n389), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n767), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n323), .A2(new_n519), .A3(new_n328), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(new_n770), .A3(new_n760), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT42), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n803), .A2(KEYINPUT42), .A3(new_n770), .A4(new_n760), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G131), .ZN(G33));
  NOR3_X1   g623(.A1(new_n635), .A2(new_n801), .A3(new_n802), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n717), .ZN(new_n811));
  XNOR2_X1  g625(.A(KEYINPUT108), .B(G134), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n811), .B(new_n812), .ZN(G36));
  NOR2_X1   g627(.A1(new_n734), .A2(new_n678), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n649), .A2(new_n758), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT43), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT43), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n649), .A2(new_n758), .A3(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT44), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n388), .A2(KEYINPUT45), .ZN(new_n823));
  OAI21_X1  g637(.A(G469), .B1(new_n388), .B2(KEYINPUT45), .ZN(new_n824));
  OAI22_X1  g638(.A1(new_n823), .A2(new_n824), .B1(new_n333), .B2(new_n295), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT46), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n384), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n767), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n825), .A2(KEYINPUT46), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n720), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n802), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n814), .A2(KEYINPUT44), .A3(new_n819), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n822), .A2(new_n832), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(G137), .ZN(G39));
  NAND4_X1  g650(.A1(new_n833), .A2(new_n709), .A3(new_n633), .A4(new_n760), .ZN(new_n837));
  NAND2_X1  g651(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT109), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT47), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n829), .A2(new_n830), .A3(new_n838), .A4(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n830), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n839), .B(new_n840), .C1(new_n843), .C2(new_n828), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n837), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(new_n392), .ZN(G42));
  INV_X1    g660(.A(new_n768), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n343), .B1(new_n368), .B2(new_n370), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT83), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n378), .A3(new_n371), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n764), .B1(new_n851), .B2(new_n295), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT49), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n634), .A2(new_n519), .A3(new_n767), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n855), .A2(new_n740), .A3(new_n815), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n854), .A2(new_n747), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n819), .A2(KEYINPUT113), .A3(new_n454), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n816), .A2(new_n454), .A3(new_n818), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT113), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n776), .A2(new_n802), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n797), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n454), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n740), .A2(new_n633), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n864), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT115), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT115), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n867), .A2(new_n870), .A3(new_n864), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n869), .A2(new_n649), .A3(new_n668), .A4(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n791), .B1(new_n859), .B2(new_n862), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT114), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT50), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n638), .B1(KEYINPUT114), .B2(KEYINPUT50), .ZN(new_n877));
  NOR4_X1   g691(.A1(new_n745), .A2(new_n746), .A3(new_n776), .A4(new_n877), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n873), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n876), .B1(new_n873), .B2(new_n878), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n865), .B(new_n872), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n873), .A2(new_n833), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n853), .A2(new_n332), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n842), .A2(new_n844), .A3(new_n883), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n858), .B1(new_n881), .B2(new_n885), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n879), .A2(new_n880), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n884), .A2(KEYINPUT116), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT116), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n842), .A2(new_n844), .A3(new_n889), .A4(new_n883), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n882), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n872), .A2(new_n865), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n887), .A2(new_n891), .A3(KEYINPUT51), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n873), .A2(new_n783), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT117), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n873), .A2(new_n896), .A3(new_n783), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n863), .A2(new_n770), .A3(new_n864), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT48), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT48), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n863), .A2(new_n901), .A3(new_n770), .A4(new_n864), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n869), .A2(new_n871), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n453), .B1(new_n904), .B2(new_n669), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n898), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n886), .A2(new_n893), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT53), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n741), .A2(new_n700), .A3(new_n714), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(new_n639), .A3(new_n390), .A4(new_n740), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n718), .A2(new_n761), .A3(new_n798), .A4(new_n910), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT52), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n769), .A2(new_n639), .ZN(new_n913));
  OAI22_X1  g727(.A1(new_n913), .A2(new_n780), .B1(new_n771), .B2(new_n690), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n790), .A2(new_n633), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n853), .A2(new_n915), .A3(new_n767), .A4(new_n640), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n517), .B(new_n432), .C1(new_n449), .C2(new_n451), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(new_n649), .B2(new_n668), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n329), .A2(new_n918), .A3(new_n519), .A4(new_n640), .ZN(new_n919));
  OAI22_X1  g733(.A1(new_n916), .A2(new_n786), .B1(new_n679), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n520), .B1(new_n705), .B2(new_n635), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n914), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n674), .A2(new_n777), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n797), .A2(new_n760), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n711), .A2(new_n517), .A3(new_n716), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n704), .A2(new_n925), .A3(new_n582), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  AOI22_X1  g741(.A1(new_n927), .A2(new_n803), .B1(new_n810), .B2(new_n717), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n922), .A2(new_n923), .A3(new_n808), .A4(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n908), .B1(new_n912), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT111), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XOR2_X1   g746(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n933));
  INV_X1    g747(.A(new_n921), .ZN(new_n934));
  INV_X1    g748(.A(new_n920), .ZN(new_n935));
  AOI22_X1  g749(.A1(new_n781), .A2(new_n783), .B1(new_n775), .B2(new_n777), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n923), .A2(new_n934), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n928), .A2(new_n808), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n582), .B1(new_n732), .B2(new_n733), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n639), .A2(new_n390), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI211_X1 g756(.A(new_n790), .B(new_n759), .C1(new_n702), .C2(new_n703), .ZN(new_n943));
  AOI22_X1  g757(.A1(new_n942), .A2(new_n717), .B1(new_n943), .B2(new_n783), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n944), .A2(KEYINPUT52), .A3(new_n761), .A4(new_n910), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT110), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT52), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n911), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  OR3_X1    g763(.A1(new_n911), .A2(new_n946), .A3(new_n947), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n939), .A2(new_n949), .A3(KEYINPUT53), .A4(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(KEYINPUT111), .B(new_n908), .C1(new_n912), .C2(new_n929), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n932), .A2(new_n933), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n911), .A2(new_n946), .A3(new_n947), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n929), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT53), .B1(new_n955), .B2(new_n949), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n945), .A2(new_n948), .ZN(new_n957));
  INV_X1    g771(.A(new_n937), .ZN(new_n958));
  INV_X1    g772(.A(new_n938), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n960), .A2(new_n908), .ZN(new_n961));
  OAI21_X1  g775(.A(KEYINPUT54), .B1(new_n956), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n907), .A2(new_n953), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT118), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OR2_X1    g779(.A1(G952), .A2(G953), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(new_n963), .B2(new_n964), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n857), .B1(new_n965), .B2(new_n967), .ZN(G75));
  NAND3_X1  g782(.A1(new_n932), .A2(new_n951), .A3(new_n952), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n969), .A2(G902), .A3(new_n322), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT56), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n257), .B1(new_n291), .B2(new_n293), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(new_n288), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT55), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n970), .A2(new_n971), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n970), .B2(new_n971), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n338), .A2(G952), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(G51));
  INV_X1    g792(.A(new_n933), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n952), .A2(new_n951), .ZN(new_n980));
  AOI21_X1  g794(.A(KEYINPUT111), .B1(new_n960), .B2(new_n908), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n979), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n953), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n385), .B(KEYINPUT57), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n851), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n823), .A2(new_n824), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n969), .A2(G902), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n977), .B1(new_n986), .B2(new_n988), .ZN(G54));
  NAND4_X1  g803(.A1(new_n969), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n990));
  INV_X1    g804(.A(new_n439), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n990), .A2(new_n991), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n992), .A2(new_n993), .A3(new_n977), .ZN(G60));
  XNOR2_X1  g808(.A(new_n666), .B(KEYINPUT119), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n953), .A2(new_n962), .ZN(new_n996));
  NAND2_X1  g810(.A1(G478), .A2(G902), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT59), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n995), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n995), .A2(new_n998), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n1000), .B1(new_n982), .B2(new_n953), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n999), .A2(new_n977), .A3(new_n1001), .ZN(G63));
  NAND2_X1  g816(.A1(G217), .A2(G902), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(KEYINPUT121), .ZN(new_n1004));
  XNOR2_X1  g818(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1006), .B1(new_n980), .B2(new_n981), .ZN(new_n1007));
  INV_X1    g821(.A(new_n615), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n969), .A2(new_n697), .A3(new_n695), .A4(new_n1006), .ZN(new_n1010));
  INV_X1    g824(.A(new_n977), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT61), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1009), .A2(new_n1010), .A3(KEYINPUT61), .A4(new_n1011), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(G66));
  INV_X1    g830(.A(G224), .ZN(new_n1017));
  OAI21_X1  g831(.A(G953), .B1(new_n456), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1018), .B(KEYINPUT122), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1019), .B1(new_n958), .B2(new_n339), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n972), .B1(G898), .B2(new_n338), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1020), .B(new_n1021), .ZN(G69));
  OAI21_X1  g836(.A(new_n339), .B1(new_n340), .B2(new_n713), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1023), .A2(KEYINPUT125), .ZN(new_n1024));
  XOR2_X1   g838(.A(new_n1024), .B(KEYINPUT126), .Z(new_n1025));
  INV_X1    g839(.A(new_n1025), .ZN(new_n1026));
  OR2_X1    g840(.A1(new_n534), .A2(new_n535), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1027), .B(new_n435), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1028), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n338), .A2(G900), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n787), .A2(new_n770), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n811), .B1(new_n831), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1032), .B1(new_n806), .B2(new_n807), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n718), .A2(new_n761), .A3(new_n798), .ZN(new_n1034));
  XNOR2_X1  g848(.A(new_n1034), .B(KEYINPUT123), .ZN(new_n1035));
  INV_X1    g849(.A(new_n845), .ZN(new_n1036));
  NAND4_X1  g850(.A1(new_n1033), .A2(new_n1035), .A3(new_n835), .A4(new_n1036), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1030), .B1(new_n1037), .B2(new_n338), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1029), .B1(new_n1038), .B2(KEYINPUT124), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1039), .B1(KEYINPUT124), .B2(new_n1038), .ZN(new_n1040));
  NAND4_X1  g854(.A1(new_n721), .A2(new_n833), .A3(new_n770), .A4(new_n918), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n835), .A2(new_n1036), .A3(new_n1041), .ZN(new_n1042));
  AND2_X1   g856(.A1(new_n1035), .A2(new_n749), .ZN(new_n1043));
  INV_X1    g857(.A(KEYINPUT62), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1035), .A2(new_n749), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1046), .A2(KEYINPUT62), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n339), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  OAI22_X1  g862(.A1(new_n1048), .A2(new_n1029), .B1(KEYINPUT125), .B2(new_n1023), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1026), .B1(new_n1040), .B2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g864(.A1(new_n1023), .A2(KEYINPUT125), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1052), .A2(new_n338), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1051), .B1(new_n1053), .B2(new_n1028), .ZN(new_n1054));
  OR2_X1    g868(.A1(new_n1038), .A2(KEYINPUT124), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1038), .A2(KEYINPUT124), .ZN(new_n1056));
  NAND3_X1  g870(.A1(new_n1055), .A2(new_n1056), .A3(new_n1029), .ZN(new_n1057));
  NAND3_X1  g871(.A1(new_n1054), .A2(new_n1025), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n1050), .A2(new_n1058), .ZN(G72));
  NAND3_X1  g873(.A1(new_n1045), .A2(new_n958), .A3(new_n1047), .ZN(new_n1060));
  NAND2_X1  g874(.A1(G472), .A2(G902), .ZN(new_n1061));
  XOR2_X1   g875(.A(new_n1061), .B(KEYINPUT63), .Z(new_n1062));
  AOI21_X1  g876(.A(new_n736), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g877(.A1(new_n956), .A2(new_n961), .ZN(new_n1064));
  INV_X1    g878(.A(new_n570), .ZN(new_n1065));
  NAND3_X1  g879(.A1(new_n1065), .A2(new_n736), .A3(new_n1062), .ZN(new_n1066));
  XOR2_X1   g880(.A(new_n1066), .B(KEYINPUT127), .Z(new_n1067));
  NOR2_X1   g881(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g882(.A(new_n1062), .B1(new_n1037), .B2(new_n937), .ZN(new_n1069));
  AND2_X1   g883(.A1(new_n1069), .A2(new_n570), .ZN(new_n1070));
  NOR4_X1   g884(.A1(new_n1063), .A2(new_n1068), .A3(new_n1070), .A4(new_n977), .ZN(G57));
endmodule


