

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592;

  XNOR2_X1 U325 ( .A(n346), .B(n312), .ZN(n508) );
  XNOR2_X1 U326 ( .A(n309), .B(n308), .ZN(n311) );
  AND2_X1 U327 ( .A1(G227GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U328 ( .A(KEYINPUT40), .B(n509), .Z(n294) );
  XNOR2_X1 U329 ( .A(n366), .B(n365), .ZN(n373) );
  XNOR2_X1 U330 ( .A(n435), .B(n293), .ZN(n308) );
  XOR2_X1 U331 ( .A(G120GAT), .B(G71GAT), .Z(n416) );
  XNOR2_X1 U332 ( .A(n373), .B(n407), .ZN(n374) );
  NOR2_X1 U333 ( .A1(n432), .A2(n431), .ZN(n433) );
  INV_X1 U334 ( .A(n499), .ZN(n500) );
  XOR2_X1 U335 ( .A(KEYINPUT48), .B(n433), .Z(n557) );
  XNOR2_X1 U336 ( .A(n502), .B(KEYINPUT106), .ZN(n503) );
  XNOR2_X1 U337 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U338 ( .A(n463), .B(n462), .ZN(G1349GAT) );
  XOR2_X1 U339 ( .A(KEYINPUT17), .B(G183GAT), .Z(n296) );
  XNOR2_X1 U340 ( .A(KEYINPUT84), .B(KEYINPUT86), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U342 ( .A(n297), .B(KEYINPUT19), .Z(n299) );
  XNOR2_X1 U343 ( .A(KEYINPUT85), .B(KEYINPUT18), .ZN(n298) );
  XNOR2_X1 U344 ( .A(n299), .B(n298), .ZN(n346) );
  XOR2_X1 U345 ( .A(KEYINPUT87), .B(KEYINPUT20), .Z(n301) );
  XNOR2_X1 U346 ( .A(G176GAT), .B(KEYINPUT83), .ZN(n300) );
  XNOR2_X1 U347 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U348 ( .A(G99GAT), .B(n416), .Z(n303) );
  XOR2_X1 U349 ( .A(G190GAT), .B(G134GAT), .Z(n375) );
  XNOR2_X1 U350 ( .A(G43GAT), .B(n375), .ZN(n302) );
  XNOR2_X1 U351 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U352 ( .A(n305), .B(n304), .Z(n309) );
  XOR2_X1 U353 ( .A(G127GAT), .B(KEYINPUT0), .Z(n307) );
  XNOR2_X1 U354 ( .A(G113GAT), .B(KEYINPUT82), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n435) );
  XNOR2_X1 U356 ( .A(G169GAT), .B(G15GAT), .ZN(n310) );
  XNOR2_X1 U357 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U358 ( .A(G218GAT), .B(G162GAT), .Z(n366) );
  XOR2_X1 U359 ( .A(G211GAT), .B(KEYINPUT21), .Z(n314) );
  XNOR2_X1 U360 ( .A(G197GAT), .B(KEYINPUT89), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n314), .B(n313), .ZN(n335) );
  XOR2_X1 U362 ( .A(n366), .B(n335), .Z(n316) );
  NAND2_X1 U363 ( .A1(G228GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n316), .B(n315), .ZN(n328) );
  XOR2_X1 U365 ( .A(KEYINPUT93), .B(KEYINPUT88), .Z(n318) );
  XNOR2_X1 U366 ( .A(KEYINPUT24), .B(KEYINPUT92), .ZN(n317) );
  XNOR2_X1 U367 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U368 ( .A(n319), .B(G106GAT), .Z(n321) );
  XOR2_X1 U369 ( .A(G141GAT), .B(G22GAT), .Z(n398) );
  XNOR2_X1 U370 ( .A(G50GAT), .B(n398), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U372 ( .A(n322), .B(KEYINPUT22), .Z(n326) );
  XOR2_X1 U373 ( .A(G78GAT), .B(G148GAT), .Z(n324) );
  XNOR2_X1 U374 ( .A(KEYINPUT74), .B(G204GAT), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n410) );
  XNOR2_X1 U376 ( .A(n410), .B(KEYINPUT23), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U379 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n330) );
  XNOR2_X1 U380 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U382 ( .A(KEYINPUT3), .B(n331), .ZN(n450) );
  XNOR2_X1 U383 ( .A(n332), .B(n450), .ZN(n477) );
  XOR2_X1 U384 ( .A(G169GAT), .B(G8GAT), .Z(n395) );
  XNOR2_X1 U385 ( .A(n395), .B(G218GAT), .ZN(n334) );
  XNOR2_X1 U386 ( .A(G176GAT), .B(G64GAT), .ZN(n333) );
  XNOR2_X1 U387 ( .A(n333), .B(KEYINPUT75), .ZN(n409) );
  XNOR2_X1 U388 ( .A(n334), .B(n409), .ZN(n339) );
  XOR2_X1 U389 ( .A(n335), .B(KEYINPUT99), .Z(n337) );
  NAND2_X1 U390 ( .A1(G226GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U391 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U392 ( .A(n339), .B(n338), .Z(n344) );
  XOR2_X1 U393 ( .A(KEYINPUT100), .B(G92GAT), .Z(n341) );
  XNOR2_X1 U394 ( .A(G190GAT), .B(G204GAT), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U396 ( .A(G36GAT), .B(n342), .ZN(n343) );
  XNOR2_X1 U397 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n506) );
  INV_X1 U399 ( .A(n506), .ZN(n532) );
  XNOR2_X1 U400 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n347) );
  XNOR2_X1 U401 ( .A(n347), .B(KEYINPUT72), .ZN(n408) );
  XOR2_X1 U402 ( .A(n408), .B(KEYINPUT81), .Z(n349) );
  NAND2_X1 U403 ( .A1(G231GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U404 ( .A(n349), .B(n348), .ZN(n364) );
  XOR2_X1 U405 ( .A(KEYINPUT80), .B(G64GAT), .Z(n351) );
  XNOR2_X1 U406 ( .A(G8GAT), .B(G211GAT), .ZN(n350) );
  XNOR2_X1 U407 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U408 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n353) );
  XNOR2_X1 U409 ( .A(KEYINPUT79), .B(KEYINPUT14), .ZN(n352) );
  XNOR2_X1 U410 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U411 ( .A(n355), .B(n354), .ZN(n362) );
  XOR2_X1 U412 ( .A(G155GAT), .B(G71GAT), .Z(n357) );
  XNOR2_X1 U413 ( .A(G183GAT), .B(G127GAT), .ZN(n356) );
  XNOR2_X1 U414 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U415 ( .A(n358), .B(G78GAT), .Z(n360) );
  XOR2_X1 U416 ( .A(G15GAT), .B(G1GAT), .Z(n394) );
  XNOR2_X1 U417 ( .A(G22GAT), .B(n394), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U419 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U420 ( .A(n364), .B(n363), .ZN(n482) );
  INV_X1 U421 ( .A(KEYINPUT36), .ZN(n388) );
  AND2_X1 U422 ( .A1(G232GAT), .A2(G233GAT), .ZN(n365) );
  INV_X1 U423 ( .A(G85GAT), .ZN(n367) );
  NAND2_X1 U424 ( .A1(G92GAT), .A2(n367), .ZN(n370) );
  INV_X1 U425 ( .A(G92GAT), .ZN(n368) );
  NAND2_X1 U426 ( .A1(n368), .A2(G85GAT), .ZN(n369) );
  NAND2_X1 U427 ( .A1(n370), .A2(n369), .ZN(n372) );
  XNOR2_X1 U428 ( .A(G99GAT), .B(G106GAT), .ZN(n371) );
  XNOR2_X1 U429 ( .A(n372), .B(n371), .ZN(n407) );
  XOR2_X1 U430 ( .A(KEYINPUT10), .B(n374), .Z(n377) );
  XNOR2_X1 U431 ( .A(n375), .B(KEYINPUT76), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n377), .B(n376), .ZN(n387) );
  XOR2_X1 U433 ( .A(G43GAT), .B(G29GAT), .Z(n379) );
  XNOR2_X1 U434 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U436 ( .A(n380), .B(KEYINPUT69), .Z(n382) );
  XNOR2_X1 U437 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n382), .B(n381), .ZN(n393) );
  XOR2_X1 U439 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n384) );
  XNOR2_X1 U440 ( .A(KEYINPUT77), .B(KEYINPUT64), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U442 ( .A(n393), .B(n385), .Z(n386) );
  XNOR2_X1 U443 ( .A(n387), .B(n386), .ZN(n569) );
  XOR2_X2 U444 ( .A(KEYINPUT78), .B(n569), .Z(n575) );
  XNOR2_X1 U445 ( .A(n388), .B(n575), .ZN(n497) );
  NOR2_X1 U446 ( .A1(n482), .A2(n497), .ZN(n389) );
  XNOR2_X1 U447 ( .A(KEYINPUT45), .B(n389), .ZN(n423) );
  XOR2_X1 U448 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n391) );
  XNOR2_X1 U449 ( .A(KEYINPUT70), .B(KEYINPUT67), .ZN(n390) );
  XNOR2_X1 U450 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n393), .B(n392), .ZN(n406) );
  XOR2_X1 U452 ( .A(G197GAT), .B(G113GAT), .Z(n397) );
  XNOR2_X1 U453 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n399) );
  XOR2_X1 U455 ( .A(n399), .B(n398), .Z(n404) );
  XOR2_X1 U456 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n401) );
  NAND2_X1 U457 ( .A1(G229GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U459 ( .A(KEYINPUT65), .B(n402), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n513) );
  XNOR2_X1 U462 ( .A(KEYINPUT71), .B(n513), .ZN(n572) );
  XOR2_X1 U463 ( .A(n408), .B(n407), .Z(n412) );
  XNOR2_X1 U464 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U465 ( .A(n412), .B(n411), .ZN(n420) );
  XOR2_X1 U466 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n414) );
  XNOR2_X1 U467 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n413) );
  XNOR2_X1 U468 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U469 ( .A(n416), .B(n415), .Z(n418) );
  NAND2_X1 U470 ( .A1(G230GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U471 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U472 ( .A(n420), .B(n419), .Z(n585) );
  INV_X1 U473 ( .A(n585), .ZN(n421) );
  NOR2_X1 U474 ( .A1(n572), .A2(n421), .ZN(n422) );
  AND2_X1 U475 ( .A1(n423), .A2(n422), .ZN(n424) );
  XOR2_X1 U476 ( .A(n424), .B(KEYINPUT117), .Z(n432) );
  INV_X1 U477 ( .A(n482), .ZN(n589) );
  XOR2_X1 U478 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n426) );
  XNOR2_X1 U479 ( .A(n585), .B(KEYINPUT41), .ZN(n561) );
  INV_X1 U480 ( .A(n513), .ZN(n580) );
  NAND2_X1 U481 ( .A1(n561), .A2(n580), .ZN(n425) );
  XOR2_X1 U482 ( .A(n426), .B(n425), .Z(n427) );
  NOR2_X1 U483 ( .A1(n589), .A2(n427), .ZN(n428) );
  NAND2_X1 U484 ( .A1(n569), .A2(n428), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n429), .B(KEYINPUT116), .ZN(n430) );
  XNOR2_X1 U486 ( .A(KEYINPUT47), .B(n430), .ZN(n431) );
  AND2_X1 U487 ( .A1(n532), .A2(n557), .ZN(n434) );
  XNOR2_X1 U488 ( .A(KEYINPUT54), .B(n434), .ZN(n457) );
  XOR2_X1 U489 ( .A(G162GAT), .B(n435), .Z(n437) );
  NAND2_X1 U490 ( .A1(G225GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n456) );
  XOR2_X1 U492 ( .A(KEYINPUT1), .B(G57GAT), .Z(n439) );
  XNOR2_X1 U493 ( .A(G141GAT), .B(G1GAT), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U495 ( .A(G85GAT), .B(G148GAT), .Z(n441) );
  XNOR2_X1 U496 ( .A(G134GAT), .B(G120GAT), .ZN(n440) );
  XNOR2_X1 U497 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n453) );
  XOR2_X1 U499 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n445) );
  XNOR2_X1 U500 ( .A(KEYINPUT97), .B(KEYINPUT4), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U502 ( .A(KEYINPUT98), .B(KEYINPUT94), .Z(n447) );
  XNOR2_X1 U503 ( .A(KEYINPUT6), .B(KEYINPUT5), .ZN(n446) );
  XNOR2_X1 U504 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U505 ( .A(n449), .B(n448), .ZN(n451) );
  XNOR2_X1 U506 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U507 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U508 ( .A(G29GAT), .B(n454), .Z(n455) );
  XNOR2_X1 U509 ( .A(n456), .B(n455), .ZN(n559) );
  NAND2_X1 U510 ( .A1(n457), .A2(n559), .ZN(n465) );
  NOR2_X1 U511 ( .A1(n477), .A2(n465), .ZN(n458) );
  XNOR2_X1 U512 ( .A(n458), .B(KEYINPUT55), .ZN(n459) );
  NOR2_X2 U513 ( .A1(n508), .A2(n459), .ZN(n576) );
  NAND2_X1 U514 ( .A1(n576), .A2(n561), .ZN(n463) );
  XOR2_X1 U515 ( .A(KEYINPUT56), .B(KEYINPUT124), .Z(n461) );
  XNOR2_X1 U516 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n460) );
  INV_X1 U517 ( .A(G218GAT), .ZN(n468) );
  NAND2_X1 U518 ( .A1(n477), .A2(n508), .ZN(n464) );
  XNOR2_X1 U519 ( .A(n464), .B(KEYINPUT26), .ZN(n472) );
  NOR2_X1 U520 ( .A1(n472), .A2(n465), .ZN(n590) );
  INV_X1 U521 ( .A(n590), .ZN(n586) );
  NOR2_X1 U522 ( .A1(n497), .A2(n586), .ZN(n466) );
  XNOR2_X1 U523 ( .A(KEYINPUT62), .B(n466), .ZN(n467) );
  XNOR2_X1 U524 ( .A(n468), .B(n467), .ZN(G1355GAT) );
  XNOR2_X1 U525 ( .A(G1GAT), .B(KEYINPUT103), .ZN(n469) );
  XNOR2_X1 U526 ( .A(n469), .B(KEYINPUT34), .ZN(n470) );
  XOR2_X1 U527 ( .A(KEYINPUT102), .B(n470), .Z(n487) );
  NAND2_X1 U528 ( .A1(n585), .A2(n572), .ZN(n499) );
  XOR2_X1 U529 ( .A(KEYINPUT27), .B(n506), .Z(n478) );
  INV_X1 U530 ( .A(n478), .ZN(n471) );
  NOR2_X1 U531 ( .A1(n472), .A2(n471), .ZN(n556) );
  NOR2_X1 U532 ( .A1(n508), .A2(n506), .ZN(n473) );
  NOR2_X1 U533 ( .A1(n477), .A2(n473), .ZN(n474) );
  XOR2_X1 U534 ( .A(KEYINPUT25), .B(n474), .Z(n475) );
  NOR2_X1 U535 ( .A1(n556), .A2(n475), .ZN(n476) );
  INV_X1 U536 ( .A(n559), .ZN(n529) );
  NOR2_X1 U537 ( .A1(n476), .A2(n529), .ZN(n481) );
  INV_X1 U538 ( .A(n508), .ZN(n541) );
  XNOR2_X1 U539 ( .A(KEYINPUT28), .B(n477), .ZN(n535) );
  NOR2_X1 U540 ( .A1(n559), .A2(n535), .ZN(n479) );
  NAND2_X1 U541 ( .A1(n479), .A2(n478), .ZN(n543) );
  NOR2_X1 U542 ( .A1(n541), .A2(n543), .ZN(n480) );
  NOR2_X1 U543 ( .A1(n481), .A2(n480), .ZN(n494) );
  NOR2_X1 U544 ( .A1(n482), .A2(n575), .ZN(n483) );
  XOR2_X1 U545 ( .A(KEYINPUT16), .B(n483), .Z(n484) );
  NOR2_X1 U546 ( .A1(n494), .A2(n484), .ZN(n485) );
  XNOR2_X1 U547 ( .A(KEYINPUT101), .B(n485), .ZN(n514) );
  NOR2_X1 U548 ( .A1(n499), .A2(n514), .ZN(n492) );
  NAND2_X1 U549 ( .A1(n492), .A2(n529), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n487), .B(n486), .ZN(G1324GAT) );
  NAND2_X1 U551 ( .A1(n492), .A2(n532), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n488), .B(KEYINPUT104), .ZN(n489) );
  XNOR2_X1 U553 ( .A(G8GAT), .B(n489), .ZN(G1325GAT) );
  XOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT35), .Z(n491) );
  NAND2_X1 U555 ( .A1(n492), .A2(n541), .ZN(n490) );
  XNOR2_X1 U556 ( .A(n491), .B(n490), .ZN(G1326GAT) );
  NAND2_X1 U557 ( .A1(n492), .A2(n535), .ZN(n493) );
  XNOR2_X1 U558 ( .A(n493), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U559 ( .A1(n494), .A2(n589), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n495), .B(KEYINPUT105), .ZN(n496) );
  NOR2_X1 U561 ( .A1(n497), .A2(n496), .ZN(n498) );
  XNOR2_X1 U562 ( .A(KEYINPUT37), .B(n498), .ZN(n527) );
  INV_X1 U563 ( .A(n527), .ZN(n501) );
  NAND2_X1 U564 ( .A1(n501), .A2(n500), .ZN(n502) );
  XNOR2_X1 U565 ( .A(KEYINPUT38), .B(n503), .ZN(n510) );
  NOR2_X1 U566 ( .A1(n559), .A2(n510), .ZN(n505) );
  XNOR2_X1 U567 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  NOR2_X1 U569 ( .A1(n506), .A2(n510), .ZN(n507) );
  XOR2_X1 U570 ( .A(G36GAT), .B(n507), .Z(G1329GAT) );
  NOR2_X1 U571 ( .A1(n508), .A2(n510), .ZN(n509) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(n294), .ZN(G1330GAT) );
  INV_X1 U573 ( .A(n535), .ZN(n511) );
  NOR2_X1 U574 ( .A1(n511), .A2(n510), .ZN(n512) );
  XOR2_X1 U575 ( .A(G50GAT), .B(n512), .Z(G1331GAT) );
  XNOR2_X1 U576 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n516) );
  NAND2_X1 U577 ( .A1(n513), .A2(n561), .ZN(n526) );
  NOR2_X1 U578 ( .A1(n526), .A2(n514), .ZN(n521) );
  NAND2_X1 U579 ( .A1(n521), .A2(n529), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(G1332GAT) );
  NAND2_X1 U581 ( .A1(n521), .A2(n532), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n517), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n519) );
  NAND2_X1 U584 ( .A1(n521), .A2(n541), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G71GAT), .B(n520), .ZN(G1334GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n523) );
  NAND2_X1 U588 ( .A1(n521), .A2(n535), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(n525) );
  XOR2_X1 U590 ( .A(G78GAT), .B(KEYINPUT110), .Z(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(G1335GAT) );
  XNOR2_X1 U592 ( .A(G85GAT), .B(KEYINPUT112), .ZN(n531) );
  NOR2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U594 ( .A(KEYINPUT111), .B(n528), .Z(n536) );
  NAND2_X1 U595 ( .A1(n536), .A2(n529), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(G1336GAT) );
  NAND2_X1 U597 ( .A1(n532), .A2(n536), .ZN(n533) );
  XNOR2_X1 U598 ( .A(G92GAT), .B(n533), .ZN(G1337GAT) );
  NAND2_X1 U599 ( .A1(n536), .A2(n541), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n534), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(KEYINPUT113), .ZN(n540) );
  XOR2_X1 U602 ( .A(KEYINPUT114), .B(KEYINPUT44), .Z(n538) );
  NAND2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(G1339GAT) );
  NAND2_X1 U606 ( .A1(n541), .A2(n557), .ZN(n542) );
  NOR2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n551) );
  NAND2_X1 U608 ( .A1(n551), .A2(n572), .ZN(n544) );
  XNOR2_X1 U609 ( .A(G113GAT), .B(n544), .ZN(G1340GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n546) );
  NAND2_X1 U611 ( .A1(n551), .A2(n561), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G120GAT), .B(n547), .ZN(G1341GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT119), .B(KEYINPUT50), .Z(n549) );
  NAND2_X1 U615 ( .A1(n551), .A2(n589), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(G127GAT), .B(n550), .ZN(G1342GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT121), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U619 ( .A1(n551), .A2(n575), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n555) );
  XOR2_X1 U621 ( .A(G134GAT), .B(KEYINPUT120), .Z(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1343GAT) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n567) );
  NAND2_X1 U625 ( .A1(n580), .A2(n567), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n563) );
  NAND2_X1 U628 ( .A1(n567), .A2(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G148GAT), .B(n564), .ZN(G1345GAT) );
  NAND2_X1 U631 ( .A1(n567), .A2(n589), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(KEYINPUT122), .ZN(n566) );
  XNOR2_X1 U633 ( .A(G155GAT), .B(n566), .ZN(G1346GAT) );
  INV_X1 U634 ( .A(n567), .ZN(n568) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G162GAT), .B(KEYINPUT123), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1347GAT) );
  NAND2_X1 U638 ( .A1(n576), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(G169GAT), .B(n573), .ZN(G1348GAT) );
  NAND2_X1 U640 ( .A1(n576), .A2(n589), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n574), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n578) );
  XOR2_X1 U643 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n579), .B(G190GAT), .ZN(G1351GAT) );
  NAND2_X1 U646 ( .A1(n580), .A2(n590), .ZN(n584) );
  XOR2_X1 U647 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n582) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n581) );
  XNOR2_X1 U649 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U651 ( .A(G204GAT), .B(KEYINPUT61), .Z(n588) );
  OR2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1353GAT) );
  XOR2_X1 U654 ( .A(G211GAT), .B(KEYINPUT127), .Z(n592) );
  NAND2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n592), .B(n591), .ZN(G1354GAT) );
endmodule

