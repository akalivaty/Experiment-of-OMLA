

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754;

  AND2_X1 U380 ( .A1(n381), .A2(n379), .ZN(n378) );
  XNOR2_X1 U381 ( .A(n583), .B(n582), .ZN(n754) );
  XNOR2_X1 U382 ( .A(n740), .B(n411), .ZN(n718) );
  XNOR2_X1 U383 ( .A(G113), .B(G143), .ZN(n476) );
  INV_X1 U384 ( .A(KEYINPUT3), .ZN(n446) );
  INV_X1 U385 ( .A(G953), .ZN(n746) );
  NAND2_X1 U386 ( .A1(n369), .A2(n707), .ZN(n703) );
  XNOR2_X2 U387 ( .A(n599), .B(KEYINPUT45), .ZN(n707) );
  NOR2_X2 U388 ( .A1(n611), .A2(n728), .ZN(n613) );
  NOR2_X2 U389 ( .A1(n632), .A2(n728), .ZN(n635) );
  NOR2_X2 U390 ( .A1(n640), .A2(n728), .ZN(n641) );
  INV_X1 U391 ( .A(n554), .ZN(n430) );
  AND2_X1 U392 ( .A1(n555), .A2(n430), .ZN(n591) );
  XNOR2_X2 U393 ( .A(n493), .B(n400), .ZN(n455) );
  NOR2_X1 U394 ( .A1(n385), .A2(KEYINPUT69), .ZN(n588) );
  INV_X1 U395 ( .A(n668), .ZN(n589) );
  INV_X1 U396 ( .A(n528), .ZN(n668) );
  NAND2_X1 U397 ( .A1(n704), .A2(n708), .ZN(n367) );
  NOR2_X1 U398 ( .A1(n377), .A2(KEYINPUT44), .ZN(n376) );
  XNOR2_X1 U399 ( .A(n389), .B(KEYINPUT65), .ZN(n724) );
  XNOR2_X1 U400 ( .A(n389), .B(KEYINPUT65), .ZN(n361) );
  NAND2_X2 U401 ( .A1(n368), .A2(n367), .ZN(n389) );
  AND2_X1 U402 ( .A1(n605), .A2(n604), .ZN(n369) );
  XNOR2_X1 U403 ( .A(n553), .B(KEYINPUT83), .ZN(n709) );
  NAND2_X1 U404 ( .A1(n378), .A2(n374), .ZN(n599) );
  NAND2_X1 U405 ( .A1(n376), .A2(n375), .ZN(n374) );
  AND2_X1 U406 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U407 ( .A(n403), .B(G137), .ZN(n416) );
  XNOR2_X1 U408 ( .A(G116), .B(G113), .ZN(n447) );
  BUF_X1 U409 ( .A(n373), .Z(n359) );
  XNOR2_X1 U410 ( .A(n389), .B(KEYINPUT65), .ZN(n360) );
  INV_X1 U411 ( .A(n586), .ZN(n362) );
  XNOR2_X1 U412 ( .A(n432), .B(n431), .ZN(n373) );
  XNOR2_X1 U413 ( .A(n429), .B(n428), .ZN(n531) );
  NOR2_X1 U414 ( .A1(n607), .A2(G902), .ZN(n429) );
  XNOR2_X2 U415 ( .A(n388), .B(n404), .ZN(n740) );
  NOR2_X2 U416 ( .A1(n699), .A2(n592), .ZN(n566) );
  XNOR2_X2 U417 ( .A(n557), .B(n556), .ZN(n699) );
  AND2_X1 U418 ( .A1(n522), .A2(n622), .ZN(n391) );
  NAND2_X1 U419 ( .A1(n382), .A2(KEYINPUT44), .ZN(n381) );
  XNOR2_X1 U420 ( .A(n387), .B(KEYINPUT1), .ZN(n555) );
  XNOR2_X1 U421 ( .A(G119), .B(G110), .ZN(n417) );
  XNOR2_X1 U422 ( .A(KEYINPUT88), .B(KEYINPUT15), .ZN(n412) );
  XNOR2_X1 U423 ( .A(n505), .B(KEYINPUT28), .ZN(n396) );
  AND2_X1 U424 ( .A1(n392), .A2(n391), .ZN(n390) );
  AND2_X1 U425 ( .A1(n517), .A2(KEYINPUT47), .ZN(n394) );
  XNOR2_X1 U426 ( .A(n380), .B(KEYINPUT101), .ZN(n379) );
  NAND2_X1 U427 ( .A1(n642), .A2(n598), .ZN(n380) );
  XNOR2_X1 U428 ( .A(G101), .B(G146), .ZN(n442) );
  XOR2_X1 U429 ( .A(G137), .B(KEYINPUT5), .Z(n443) );
  XNOR2_X1 U430 ( .A(G131), .B(G104), .ZN(n475) );
  INV_X1 U431 ( .A(KEYINPUT70), .ZN(n403) );
  BUF_X1 U432 ( .A(n707), .Z(n729) );
  XNOR2_X1 U433 ( .A(G107), .B(G104), .ZN(n405) );
  INV_X1 U434 ( .A(KEYINPUT4), .ZN(n400) );
  AND2_X1 U435 ( .A1(n395), .A2(n507), .ZN(n515) );
  XNOR2_X1 U436 ( .A(n504), .B(n396), .ZN(n395) );
  XNOR2_X1 U437 ( .A(n366), .B(KEYINPUT75), .ZN(n397) );
  NAND2_X1 U438 ( .A1(n373), .A2(n441), .ZN(n366) );
  INV_X1 U439 ( .A(KEYINPUT32), .ZN(n582) );
  INV_X1 U440 ( .A(G122), .ZN(n384) );
  XOR2_X1 U441 ( .A(G128), .B(KEYINPUT23), .Z(n363) );
  AND2_X1 U442 ( .A1(n454), .A2(n685), .ZN(n364) );
  XNOR2_X2 U443 ( .A(n365), .B(KEYINPUT39), .ZN(n499) );
  NAND2_X1 U444 ( .A1(n397), .A2(n364), .ZN(n365) );
  NAND2_X1 U445 ( .A1(n709), .A2(n707), .ZN(n704) );
  AND2_X2 U446 ( .A1(n703), .A2(n606), .ZN(n368) );
  NAND2_X1 U447 ( .A1(n541), .A2(n370), .ZN(n543) );
  XNOR2_X1 U448 ( .A(n371), .B(n513), .ZN(n370) );
  NAND2_X1 U449 ( .A1(n626), .A2(n623), .ZN(n371) );
  XNOR2_X1 U450 ( .A(n372), .B(n501), .ZN(n626) );
  NAND2_X1 U451 ( .A1(n499), .A2(n654), .ZN(n372) );
  NAND2_X1 U452 ( .A1(n359), .A2(n589), .ZN(n590) );
  XNOR2_X1 U453 ( .A(n385), .B(KEYINPUT69), .ZN(n375) );
  XNOR2_X2 U454 ( .A(n570), .B(n569), .ZN(n385) );
  INV_X1 U455 ( .A(n383), .ZN(n377) );
  NAND2_X1 U456 ( .A1(n588), .A2(n383), .ZN(n382) );
  NOR2_X2 U457 ( .A1(n650), .A2(n754), .ZN(n383) );
  XNOR2_X1 U458 ( .A(n385), .B(n384), .ZN(G24) );
  XNOR2_X2 U459 ( .A(n386), .B(G469), .ZN(n387) );
  OR2_X2 U460 ( .A1(n718), .A2(G902), .ZN(n386) );
  NAND2_X1 U461 ( .A1(n387), .A2(n430), .ZN(n432) );
  XNOR2_X1 U462 ( .A(n387), .B(n506), .ZN(n507) );
  INV_X1 U463 ( .A(n499), .ZN(n551) );
  XNOR2_X1 U464 ( .A(n450), .B(n388), .ZN(n614) );
  XNOR2_X2 U465 ( .A(n455), .B(n402), .ZN(n388) );
  NAND2_X1 U466 ( .A1(n393), .A2(n390), .ZN(n540) );
  NAND2_X1 U467 ( .A1(n655), .A2(n520), .ZN(n392) );
  XNOR2_X1 U468 ( .A(n394), .B(KEYINPUT81), .ZN(n393) );
  XNOR2_X2 U469 ( .A(n399), .B(G128), .ZN(n493) );
  NAND2_X1 U470 ( .A1(n515), .A2(n562), .ZN(n516) );
  AND2_X1 U471 ( .A1(n397), .A2(n454), .ZN(n527) );
  AND2_X1 U472 ( .A1(n471), .A2(G210), .ZN(n398) );
  NAND2_X1 U473 ( .A1(G234), .A2(n746), .ZN(n421) );
  INV_X1 U474 ( .A(n664), .ZN(n571) );
  XNOR2_X1 U475 ( .A(n449), .B(n466), .ZN(n450) );
  BUF_X1 U476 ( .A(n709), .Z(n745) );
  INV_X1 U477 ( .A(n728), .ZN(n618) );
  XNOR2_X1 U478 ( .A(KEYINPUT84), .B(KEYINPUT35), .ZN(n569) );
  INV_X1 U479 ( .A(KEYINPUT125), .ZN(n612) );
  XNOR2_X2 U480 ( .A(G143), .B(KEYINPUT64), .ZN(n399) );
  XNOR2_X1 U481 ( .A(G134), .B(G131), .ZN(n401) );
  XNOR2_X1 U482 ( .A(n401), .B(KEYINPUT71), .ZN(n402) );
  XNOR2_X1 U483 ( .A(n416), .B(KEYINPUT92), .ZN(n404) );
  XNOR2_X1 U484 ( .A(n405), .B(G110), .ZN(n407) );
  XNOR2_X1 U485 ( .A(G101), .B(KEYINPUT89), .ZN(n406) );
  XNOR2_X1 U486 ( .A(n407), .B(n406), .ZN(n467) );
  XOR2_X1 U487 ( .A(G146), .B(G140), .Z(n409) );
  NAND2_X1 U488 ( .A1(G227), .A2(n746), .ZN(n408) );
  XNOR2_X1 U489 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U490 ( .A(n467), .B(n410), .ZN(n411) );
  XNOR2_X1 U491 ( .A(n412), .B(G902), .ZN(n470) );
  NAND2_X1 U492 ( .A1(n470), .A2(G234), .ZN(n413) );
  XNOR2_X1 U493 ( .A(KEYINPUT20), .B(n413), .ZN(n425) );
  NAND2_X1 U494 ( .A1(G221), .A2(n425), .ZN(n414) );
  XNOR2_X1 U495 ( .A(n414), .B(KEYINPUT21), .ZN(n665) );
  XNOR2_X1 U496 ( .A(n665), .B(KEYINPUT93), .ZN(n576) );
  XNOR2_X1 U497 ( .A(G146), .B(G125), .ZN(n457) );
  XOR2_X1 U498 ( .A(KEYINPUT10), .B(G140), .Z(n415) );
  XNOR2_X1 U499 ( .A(n457), .B(n415), .ZN(n741) );
  XNOR2_X1 U500 ( .A(n417), .B(n416), .ZN(n420) );
  XOR2_X1 U501 ( .A(KEYINPUT24), .B(KEYINPUT72), .Z(n418) );
  XNOR2_X1 U502 ( .A(n418), .B(n363), .ZN(n419) );
  XNOR2_X1 U503 ( .A(n420), .B(n419), .ZN(n423) );
  XOR2_X1 U504 ( .A(KEYINPUT8), .B(n421), .Z(n491) );
  NAND2_X1 U505 ( .A1(G221), .A2(n491), .ZN(n422) );
  XNOR2_X1 U506 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U507 ( .A(n741), .B(n424), .ZN(n607) );
  XOR2_X1 U508 ( .A(KEYINPUT76), .B(KEYINPUT25), .Z(n427) );
  NAND2_X1 U509 ( .A1(G217), .A2(n425), .ZN(n426) );
  XOR2_X1 U510 ( .A(n427), .B(n426), .Z(n428) );
  NAND2_X1 U511 ( .A1(n576), .A2(n531), .ZN(n554) );
  INV_X1 U512 ( .A(KEYINPUT94), .ZN(n431) );
  NAND2_X1 U513 ( .A1(G234), .A2(G237), .ZN(n433) );
  XNOR2_X1 U514 ( .A(KEYINPUT14), .B(n433), .ZN(n437) );
  AND2_X1 U515 ( .A1(G953), .A2(G902), .ZN(n434) );
  NAND2_X1 U516 ( .A1(n437), .A2(n434), .ZN(n558) );
  XNOR2_X1 U517 ( .A(n558), .B(KEYINPUT103), .ZN(n436) );
  INV_X1 U518 ( .A(G900), .ZN(n435) );
  NAND2_X1 U519 ( .A1(n436), .A2(n435), .ZN(n440) );
  NAND2_X1 U520 ( .A1(G952), .A2(n437), .ZN(n696) );
  NOR2_X1 U521 ( .A1(n696), .A2(G953), .ZN(n439) );
  INV_X1 U522 ( .A(KEYINPUT90), .ZN(n438) );
  XNOR2_X1 U523 ( .A(n439), .B(n438), .ZN(n560) );
  AND2_X1 U524 ( .A1(n440), .A2(n560), .ZN(n502) );
  INV_X1 U525 ( .A(n502), .ZN(n441) );
  XNOR2_X1 U526 ( .A(n443), .B(n442), .ZN(n445) );
  NOR2_X1 U527 ( .A1(G953), .A2(G237), .ZN(n473) );
  NAND2_X1 U528 ( .A1(n473), .A2(G210), .ZN(n444) );
  XNOR2_X1 U529 ( .A(n445), .B(n444), .ZN(n449) );
  XNOR2_X1 U530 ( .A(n446), .B(G119), .ZN(n448) );
  XNOR2_X1 U531 ( .A(n448), .B(n447), .ZN(n466) );
  NOR2_X1 U532 ( .A1(n614), .A2(G902), .ZN(n451) );
  XNOR2_X1 U533 ( .A(G472), .B(n451), .ZN(n528) );
  INV_X1 U534 ( .A(G902), .ZN(n496) );
  INV_X1 U535 ( .A(G237), .ZN(n452) );
  NAND2_X1 U536 ( .A1(n496), .A2(n452), .ZN(n471) );
  NAND2_X1 U537 ( .A1(n471), .A2(G214), .ZN(n684) );
  INV_X1 U538 ( .A(n684), .ZN(n508) );
  NOR2_X1 U539 ( .A1(n589), .A2(n508), .ZN(n453) );
  XNOR2_X1 U540 ( .A(n453), .B(KEYINPUT30), .ZN(n454) );
  INV_X1 U541 ( .A(n455), .ZN(n462) );
  XNOR2_X1 U542 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n456) );
  XNOR2_X1 U543 ( .A(n457), .B(n456), .ZN(n460) );
  NAND2_X1 U544 ( .A1(n746), .A2(G224), .ZN(n458) );
  XNOR2_X1 U545 ( .A(n458), .B(KEYINPUT77), .ZN(n459) );
  XNOR2_X1 U546 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U547 ( .A(n462), .B(n461), .ZN(n469) );
  XNOR2_X1 U548 ( .A(KEYINPUT74), .B(KEYINPUT16), .ZN(n464) );
  XNOR2_X1 U549 ( .A(G122), .B(KEYINPUT73), .ZN(n463) );
  XNOR2_X1 U550 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U551 ( .A(n466), .B(n465), .ZN(n468) );
  XNOR2_X1 U552 ( .A(n468), .B(n467), .ZN(n734) );
  XNOR2_X1 U553 ( .A(n469), .B(n734), .ZN(n637) );
  INV_X1 U554 ( .A(n470), .ZN(n606) );
  OR2_X1 U555 ( .A1(n637), .A2(n606), .ZN(n472) );
  XNOR2_X2 U556 ( .A(n472), .B(n398), .ZN(n525) );
  INV_X1 U557 ( .A(n525), .ZN(n547) );
  XNOR2_X1 U558 ( .A(n547), .B(KEYINPUT38), .ZN(n685) );
  NAND2_X1 U559 ( .A1(G214), .A2(n473), .ZN(n474) );
  XNOR2_X1 U560 ( .A(n741), .B(n474), .ZN(n481) );
  XNOR2_X1 U561 ( .A(n475), .B(KEYINPUT12), .ZN(n479) );
  XOR2_X1 U562 ( .A(KEYINPUT11), .B(G122), .Z(n477) );
  XNOR2_X1 U563 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U564 ( .A(n479), .B(n478), .Z(n480) );
  XNOR2_X1 U565 ( .A(n481), .B(n480), .ZN(n629) );
  NOR2_X1 U566 ( .A1(G902), .A2(n629), .ZN(n483) );
  XNOR2_X1 U567 ( .A(KEYINPUT13), .B(KEYINPUT96), .ZN(n482) );
  XNOR2_X1 U568 ( .A(n483), .B(n482), .ZN(n485) );
  XNOR2_X1 U569 ( .A(KEYINPUT95), .B(G475), .ZN(n484) );
  XNOR2_X1 U570 ( .A(n485), .B(n484), .ZN(n524) );
  XOR2_X1 U571 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n487) );
  XNOR2_X1 U572 ( .A(G116), .B(G134), .ZN(n486) );
  XNOR2_X1 U573 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U574 ( .A(n488), .B(KEYINPUT97), .Z(n490) );
  XNOR2_X1 U575 ( .A(G107), .B(G122), .ZN(n489) );
  XNOR2_X1 U576 ( .A(n490), .B(n489), .ZN(n495) );
  NAND2_X1 U577 ( .A1(G217), .A2(n491), .ZN(n492) );
  XNOR2_X1 U578 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U579 ( .A(n495), .B(n494), .ZN(n726) );
  NAND2_X1 U580 ( .A1(n726), .A2(n496), .ZN(n498) );
  XNOR2_X1 U581 ( .A(KEYINPUT98), .B(G478), .ZN(n497) );
  XNOR2_X1 U582 ( .A(n498), .B(n497), .ZN(n518) );
  OR2_X1 U583 ( .A1(n524), .A2(n518), .ZN(n658) );
  INV_X1 U584 ( .A(KEYINPUT107), .ZN(n500) );
  XNOR2_X1 U585 ( .A(n500), .B(KEYINPUT40), .ZN(n501) );
  NOR2_X1 U586 ( .A1(n665), .A2(n502), .ZN(n529) );
  NOR2_X1 U587 ( .A1(n528), .A2(n531), .ZN(n503) );
  NAND2_X1 U588 ( .A1(n529), .A2(n503), .ZN(n504) );
  INV_X1 U589 ( .A(KEYINPUT106), .ZN(n505) );
  INV_X1 U590 ( .A(KEYINPUT105), .ZN(n506) );
  INV_X1 U591 ( .A(n518), .ZN(n523) );
  NAND2_X1 U592 ( .A1(n524), .A2(n523), .ZN(n686) );
  NOR2_X1 U593 ( .A1(n686), .A2(n508), .ZN(n509) );
  NAND2_X1 U594 ( .A1(n509), .A2(n685), .ZN(n510) );
  XNOR2_X1 U595 ( .A(n510), .B(KEYINPUT41), .ZN(n697) );
  NAND2_X1 U596 ( .A1(n515), .A2(n697), .ZN(n512) );
  XNOR2_X1 U597 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n511) );
  XNOR2_X1 U598 ( .A(n512), .B(n511), .ZN(n623) );
  XNOR2_X1 U599 ( .A(KEYINPUT85), .B(KEYINPUT46), .ZN(n513) );
  NAND2_X1 U600 ( .A1(n525), .A2(n684), .ZN(n514) );
  XNOR2_X1 U601 ( .A(n514), .B(KEYINPUT19), .ZN(n562) );
  XOR2_X1 U602 ( .A(n516), .B(KEYINPUT79), .Z(n517) );
  INV_X1 U603 ( .A(n517), .ZN(n655) );
  AND2_X1 U604 ( .A1(n524), .A2(n518), .ZN(n651) );
  INV_X1 U605 ( .A(n658), .ZN(n654) );
  NOR2_X1 U606 ( .A1(n651), .A2(n654), .ZN(n519) );
  XNOR2_X1 U607 ( .A(KEYINPUT99), .B(n519), .ZN(n681) );
  INV_X1 U608 ( .A(n681), .ZN(n521) );
  NOR2_X1 U609 ( .A1(n521), .A2(KEYINPUT47), .ZN(n520) );
  NAND2_X1 U610 ( .A1(n521), .A2(KEYINPUT47), .ZN(n522) );
  NOR2_X1 U611 ( .A1(n524), .A2(n523), .ZN(n567) );
  AND2_X1 U612 ( .A1(n567), .A2(n525), .ZN(n526) );
  NAND2_X1 U613 ( .A1(n527), .A2(n526), .ZN(n622) );
  XOR2_X1 U614 ( .A(n528), .B(KEYINPUT6), .Z(n596) );
  NAND2_X1 U615 ( .A1(n529), .A2(n684), .ZN(n530) );
  NOR2_X1 U616 ( .A1(n596), .A2(n530), .ZN(n533) );
  NOR2_X1 U617 ( .A1(n362), .A2(n658), .ZN(n532) );
  NAND2_X1 U618 ( .A1(n533), .A2(n532), .ZN(n544) );
  NOR2_X1 U619 ( .A1(n544), .A2(n547), .ZN(n534) );
  XNOR2_X1 U620 ( .A(n534), .B(KEYINPUT36), .ZN(n536) );
  BUF_X2 U621 ( .A(n555), .Z(n584) );
  INV_X1 U622 ( .A(KEYINPUT87), .ZN(n535) );
  XNOR2_X1 U623 ( .A(n584), .B(n535), .ZN(n574) );
  NAND2_X1 U624 ( .A1(n536), .A2(n574), .ZN(n538) );
  INV_X1 U625 ( .A(KEYINPUT109), .ZN(n537) );
  XNOR2_X1 U626 ( .A(n538), .B(n537), .ZN(n752) );
  INV_X1 U627 ( .A(n752), .ZN(n539) );
  NOR2_X1 U628 ( .A1(n540), .A2(n539), .ZN(n541) );
  INV_X1 U629 ( .A(KEYINPUT48), .ZN(n542) );
  XNOR2_X1 U630 ( .A(n543), .B(n542), .ZN(n601) );
  NOR2_X1 U631 ( .A1(n544), .A2(n584), .ZN(n546) );
  INV_X1 U632 ( .A(KEYINPUT43), .ZN(n545) );
  XNOR2_X1 U633 ( .A(n546), .B(n545), .ZN(n548) );
  NAND2_X1 U634 ( .A1(n548), .A2(n547), .ZN(n550) );
  INV_X1 U635 ( .A(KEYINPUT104), .ZN(n549) );
  XNOR2_X1 U636 ( .A(n550), .B(n549), .ZN(n753) );
  INV_X1 U637 ( .A(n753), .ZN(n600) );
  INV_X1 U638 ( .A(n651), .ZN(n661) );
  OR2_X1 U639 ( .A1(n551), .A2(n661), .ZN(n625) );
  AND2_X1 U640 ( .A1(n600), .A2(n625), .ZN(n552) );
  NAND2_X1 U641 ( .A1(n601), .A2(n552), .ZN(n553) );
  INV_X1 U642 ( .A(n596), .ZN(n572) );
  NAND2_X1 U643 ( .A1(n591), .A2(n572), .ZN(n557) );
  XOR2_X1 U644 ( .A(KEYINPUT102), .B(KEYINPUT33), .Z(n556) );
  NOR2_X1 U645 ( .A1(G898), .A2(n558), .ZN(n559) );
  XNOR2_X1 U646 ( .A(KEYINPUT91), .B(n559), .ZN(n561) );
  NAND2_X1 U647 ( .A1(n561), .A2(n560), .ZN(n563) );
  AND2_X1 U648 ( .A1(n563), .A2(n562), .ZN(n565) );
  XOR2_X1 U649 ( .A(KEYINPUT86), .B(KEYINPUT0), .Z(n564) );
  XNOR2_X1 U650 ( .A(n565), .B(n564), .ZN(n592) );
  XNOR2_X1 U651 ( .A(n566), .B(KEYINPUT34), .ZN(n568) );
  NAND2_X1 U652 ( .A1(n568), .A2(n567), .ZN(n570) );
  XOR2_X1 U653 ( .A(KEYINPUT100), .B(n362), .Z(n664) );
  NOR2_X1 U654 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U655 ( .A(KEYINPUT78), .B(n575), .ZN(n581) );
  INV_X1 U656 ( .A(n686), .ZN(n577) );
  NAND2_X1 U657 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U658 ( .A1(n592), .A2(n578), .ZN(n580) );
  XNOR2_X1 U659 ( .A(KEYINPUT22), .B(KEYINPUT66), .ZN(n579) );
  XNOR2_X1 U660 ( .A(n580), .B(n579), .ZN(n585) );
  NAND2_X1 U661 ( .A1(n581), .A2(n585), .ZN(n583) );
  INV_X1 U662 ( .A(n584), .ZN(n670) );
  NAND2_X1 U663 ( .A1(n585), .A2(n670), .ZN(n595) );
  INV_X1 U664 ( .A(n531), .ZN(n586) );
  NAND2_X1 U665 ( .A1(n589), .A2(n586), .ZN(n587) );
  NOR2_X1 U666 ( .A1(n595), .A2(n587), .ZN(n650) );
  OR2_X1 U667 ( .A1(n592), .A2(n590), .ZN(n646) );
  NAND2_X1 U668 ( .A1(n668), .A2(n591), .ZN(n675) );
  NOR2_X1 U669 ( .A1(n675), .A2(n592), .ZN(n593) );
  XNOR2_X1 U670 ( .A(n593), .B(KEYINPUT31), .ZN(n660) );
  NAND2_X1 U671 ( .A1(n646), .A2(n660), .ZN(n594) );
  NAND2_X1 U672 ( .A1(n594), .A2(n681), .ZN(n598) );
  NOR2_X1 U673 ( .A1(n664), .A2(n595), .ZN(n597) );
  NAND2_X1 U674 ( .A1(n597), .A2(n596), .ZN(n642) );
  INV_X1 U675 ( .A(KEYINPUT2), .ZN(n708) );
  AND2_X1 U676 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U677 ( .A1(n625), .A2(KEYINPUT2), .ZN(n603) );
  INV_X1 U678 ( .A(KEYINPUT80), .ZN(n602) );
  XNOR2_X1 U679 ( .A(n603), .B(n602), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n361), .A2(G217), .ZN(n609) );
  XNOR2_X1 U681 ( .A(n607), .B(KEYINPUT124), .ZN(n608) );
  XNOR2_X1 U682 ( .A(n609), .B(n608), .ZN(n611) );
  INV_X1 U683 ( .A(G952), .ZN(n610) );
  AND2_X1 U684 ( .A1(n610), .A2(G953), .ZN(n728) );
  XNOR2_X1 U685 ( .A(n613), .B(n612), .ZN(G66) );
  NAND2_X1 U686 ( .A1(n360), .A2(G472), .ZN(n616) );
  XNOR2_X1 U687 ( .A(n614), .B(KEYINPUT62), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n616), .B(n615), .ZN(n617) );
  INV_X1 U689 ( .A(n617), .ZN(n619) );
  NAND2_X1 U690 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U691 ( .A(n620), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U692 ( .A(G143), .B(KEYINPUT112), .ZN(n621) );
  XNOR2_X1 U693 ( .A(n622), .B(n621), .ZN(G45) );
  XNOR2_X1 U694 ( .A(n623), .B(G137), .ZN(G39) );
  XOR2_X1 U695 ( .A(G134), .B(KEYINPUT115), .Z(n624) );
  XNOR2_X1 U696 ( .A(n625), .B(n624), .ZN(G36) );
  BUF_X1 U697 ( .A(n626), .Z(n627) );
  XNOR2_X1 U698 ( .A(n627), .B(G131), .ZN(G33) );
  NAND2_X1 U699 ( .A1(n724), .A2(G475), .ZN(n631) );
  XNOR2_X1 U700 ( .A(KEYINPUT67), .B(KEYINPUT59), .ZN(n628) );
  XNOR2_X1 U701 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U702 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U703 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n633) );
  XOR2_X1 U704 ( .A(n633), .B(KEYINPUT68), .Z(n634) );
  XNOR2_X1 U705 ( .A(n635), .B(n634), .ZN(G60) );
  NAND2_X1 U706 ( .A1(n724), .A2(G210), .ZN(n639) );
  XOR2_X1 U707 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n636) );
  XNOR2_X1 U708 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U709 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U710 ( .A(n641), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U711 ( .A(G101), .B(n642), .ZN(G3) );
  NOR2_X1 U712 ( .A1(n658), .A2(n646), .ZN(n644) );
  XNOR2_X1 U713 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U715 ( .A(G104), .B(n645), .ZN(G6) );
  NOR2_X1 U716 ( .A1(n661), .A2(n646), .ZN(n648) );
  XNOR2_X1 U717 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U719 ( .A(G107), .B(n649), .ZN(G9) );
  XOR2_X1 U720 ( .A(G110), .B(n650), .Z(G12) );
  XOR2_X1 U721 ( .A(G128), .B(KEYINPUT29), .Z(n653) );
  NAND2_X1 U722 ( .A1(n655), .A2(n651), .ZN(n652) );
  XNOR2_X1 U723 ( .A(n653), .B(n652), .ZN(G30) );
  XOR2_X1 U724 ( .A(G146), .B(KEYINPUT113), .Z(n657) );
  NAND2_X1 U725 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U726 ( .A(n657), .B(n656), .ZN(G48) );
  NOR2_X1 U727 ( .A1(n658), .A2(n660), .ZN(n659) );
  XOR2_X1 U728 ( .A(G113), .B(n659), .Z(G15) );
  NOR2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U730 ( .A(KEYINPUT114), .B(n662), .Z(n663) );
  XNOR2_X1 U731 ( .A(G116), .B(n663), .ZN(G18) );
  NAND2_X1 U732 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U733 ( .A(KEYINPUT49), .B(n666), .ZN(n667) );
  NOR2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U735 ( .A(n669), .B(KEYINPUT116), .ZN(n674) );
  XOR2_X1 U736 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n672) );
  NAND2_X1 U737 ( .A1(n670), .A2(n554), .ZN(n671) );
  XNOR2_X1 U738 ( .A(n672), .B(n671), .ZN(n673) );
  NAND2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n676) );
  NAND2_X1 U740 ( .A1(n676), .A2(n675), .ZN(n678) );
  XOR2_X1 U741 ( .A(KEYINPUT51), .B(KEYINPUT118), .Z(n677) );
  XNOR2_X1 U742 ( .A(n678), .B(n677), .ZN(n679) );
  NAND2_X1 U743 ( .A1(n679), .A2(n697), .ZN(n680) );
  XNOR2_X1 U744 ( .A(n680), .B(KEYINPUT119), .ZN(n692) );
  NAND2_X1 U745 ( .A1(n681), .A2(n684), .ZN(n683) );
  INV_X1 U746 ( .A(n685), .ZN(n682) );
  NOR2_X1 U747 ( .A1(n683), .A2(n682), .ZN(n689) );
  NOR2_X1 U748 ( .A1(n685), .A2(n684), .ZN(n687) );
  NOR2_X1 U749 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U750 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U751 ( .A1(n699), .A2(n690), .ZN(n691) );
  NOR2_X1 U752 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U753 ( .A(n693), .B(KEYINPUT52), .ZN(n694) );
  XNOR2_X1 U754 ( .A(KEYINPUT120), .B(n694), .ZN(n695) );
  NOR2_X1 U755 ( .A1(n696), .A2(n695), .ZN(n701) );
  INV_X1 U756 ( .A(n697), .ZN(n698) );
  NOR2_X1 U757 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U758 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U759 ( .A(n702), .B(KEYINPUT121), .ZN(n715) );
  AND2_X1 U760 ( .A1(n708), .A2(KEYINPUT82), .ZN(n705) );
  NAND2_X1 U761 ( .A1(n704), .A2(n705), .ZN(n706) );
  NAND2_X1 U762 ( .A1(n703), .A2(n706), .ZN(n713) );
  NAND2_X1 U763 ( .A1(n729), .A2(n708), .ZN(n710) );
  NOR2_X1 U764 ( .A1(n710), .A2(n745), .ZN(n711) );
  NOR2_X1 U765 ( .A1(KEYINPUT82), .A2(n711), .ZN(n712) );
  NOR2_X1 U766 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U767 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U768 ( .A1(n746), .A2(n716), .ZN(n717) );
  XOR2_X1 U769 ( .A(KEYINPUT53), .B(n717), .Z(G75) );
  NAND2_X1 U770 ( .A1(n360), .A2(G469), .ZN(n722) );
  XNOR2_X1 U771 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n719) );
  XOR2_X1 U772 ( .A(n719), .B(KEYINPUT57), .Z(n720) );
  XNOR2_X1 U773 ( .A(n718), .B(n720), .ZN(n721) );
  XNOR2_X1 U774 ( .A(n722), .B(n721), .ZN(n723) );
  NOR2_X1 U775 ( .A1(n728), .A2(n723), .ZN(G54) );
  NAND2_X1 U776 ( .A1(n361), .A2(G478), .ZN(n725) );
  XOR2_X1 U777 ( .A(n726), .B(n725), .Z(n727) );
  NOR2_X1 U778 ( .A1(n728), .A2(n727), .ZN(G63) );
  NAND2_X1 U779 ( .A1(n746), .A2(n729), .ZN(n733) );
  NAND2_X1 U780 ( .A1(G953), .A2(G224), .ZN(n730) );
  XNOR2_X1 U781 ( .A(KEYINPUT61), .B(n730), .ZN(n731) );
  NAND2_X1 U782 ( .A1(n731), .A2(G898), .ZN(n732) );
  NAND2_X1 U783 ( .A1(n733), .A2(n732), .ZN(n738) );
  INV_X1 U784 ( .A(n734), .ZN(n736) );
  NOR2_X1 U785 ( .A1(G898), .A2(n746), .ZN(n735) );
  NOR2_X1 U786 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U787 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U788 ( .A(KEYINPUT126), .B(n739), .ZN(G69) );
  XOR2_X1 U789 ( .A(n740), .B(n741), .Z(n744) );
  XOR2_X1 U790 ( .A(G227), .B(n744), .Z(n742) );
  NOR2_X1 U791 ( .A1(n746), .A2(n742), .ZN(n743) );
  NAND2_X1 U792 ( .A1(n743), .A2(G900), .ZN(n749) );
  XNOR2_X1 U793 ( .A(n745), .B(n744), .ZN(n747) );
  NAND2_X1 U794 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U795 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U796 ( .A(n750), .B(KEYINPUT127), .ZN(G72) );
  XOR2_X1 U797 ( .A(G125), .B(KEYINPUT37), .Z(n751) );
  XNOR2_X1 U798 ( .A(n752), .B(n751), .ZN(G27) );
  XOR2_X1 U799 ( .A(G140), .B(n753), .Z(G42) );
  XOR2_X1 U800 ( .A(G119), .B(n754), .Z(G21) );
endmodule

