

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U550 ( .A(n691), .B(KEYINPUT64), .ZN(n709) );
  NOR2_X1 U551 ( .A1(n967), .A2(n704), .ZN(n703) );
  XNOR2_X1 U552 ( .A(n756), .B(KEYINPUT103), .ZN(n759) );
  XOR2_X1 U553 ( .A(KEYINPUT102), .B(n736), .Z(n513) );
  XOR2_X1 U554 ( .A(n721), .B(KEYINPUT29), .Z(n514) );
  INV_X1 U555 ( .A(KEYINPUT28), .ZN(n702) );
  INV_X1 U556 ( .A(n709), .ZN(n737) );
  NOR2_X1 U557 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U558 ( .A1(G651), .A2(n622), .ZN(n638) );
  NOR2_X2 U559 ( .A1(n515), .A2(G2105), .ZN(n890) );
  INV_X1 U560 ( .A(G2104), .ZN(n515) );
  NAND2_X1 U561 ( .A1(G101), .A2(n890), .ZN(n517) );
  XOR2_X1 U562 ( .A(KEYINPUT66), .B(KEYINPUT23), .Z(n516) );
  XNOR2_X1 U563 ( .A(n517), .B(n516), .ZN(n519) );
  AND2_X1 U564 ( .A1(n515), .A2(G2105), .ZN(n884) );
  NAND2_X1 U565 ( .A1(n884), .A2(G125), .ZN(n518) );
  NAND2_X1 U566 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U567 ( .A(n520), .B(KEYINPUT67), .ZN(n679) );
  NOR2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n521) );
  XOR2_X2 U569 ( .A(KEYINPUT17), .B(n521), .Z(n891) );
  NAND2_X1 U570 ( .A1(G137), .A2(n891), .ZN(n676) );
  AND2_X1 U571 ( .A1(n679), .A2(n676), .ZN(n523) );
  AND2_X1 U572 ( .A1(G2104), .A2(G2105), .ZN(n885) );
  NAND2_X1 U573 ( .A1(G113), .A2(n885), .ZN(n522) );
  XNOR2_X1 U574 ( .A(KEYINPUT68), .B(n522), .ZN(n675) );
  AND2_X1 U575 ( .A1(n523), .A2(n675), .ZN(G160) );
  XOR2_X1 U576 ( .A(G543), .B(KEYINPUT0), .Z(n622) );
  NAND2_X1 U577 ( .A1(G47), .A2(n638), .ZN(n526) );
  INV_X1 U578 ( .A(G651), .ZN(n527) );
  NOR2_X1 U579 ( .A1(G543), .A2(n527), .ZN(n524) );
  XOR2_X1 U580 ( .A(KEYINPUT1), .B(n524), .Z(n639) );
  NAND2_X1 U581 ( .A1(G60), .A2(n639), .ZN(n525) );
  NAND2_X1 U582 ( .A1(n526), .A2(n525), .ZN(n531) );
  NOR2_X1 U583 ( .A1(G543), .A2(G651), .ZN(n642) );
  NAND2_X1 U584 ( .A1(G85), .A2(n642), .ZN(n529) );
  NOR2_X1 U585 ( .A1(n622), .A2(n527), .ZN(n636) );
  NAND2_X1 U586 ( .A1(G72), .A2(n636), .ZN(n528) );
  NAND2_X1 U587 ( .A1(n529), .A2(n528), .ZN(n530) );
  OR2_X1 U588 ( .A1(n531), .A2(n530), .ZN(G290) );
  NAND2_X1 U589 ( .A1(G90), .A2(n642), .ZN(n533) );
  NAND2_X1 U590 ( .A1(G77), .A2(n636), .ZN(n532) );
  NAND2_X1 U591 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U592 ( .A(n534), .B(KEYINPUT9), .ZN(n536) );
  NAND2_X1 U593 ( .A1(G64), .A2(n639), .ZN(n535) );
  NAND2_X1 U594 ( .A1(n536), .A2(n535), .ZN(n539) );
  NAND2_X1 U595 ( .A1(G52), .A2(n638), .ZN(n537) );
  XNOR2_X1 U596 ( .A(KEYINPUT69), .B(n537), .ZN(n538) );
  NOR2_X1 U597 ( .A1(n539), .A2(n538), .ZN(G171) );
  AND2_X1 U598 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U599 ( .A(G132), .ZN(G219) );
  INV_X1 U600 ( .A(G82), .ZN(G220) );
  INV_X1 U601 ( .A(G57), .ZN(G237) );
  INV_X1 U602 ( .A(G120), .ZN(G236) );
  INV_X1 U603 ( .A(G69), .ZN(G235) );
  AND2_X1 U604 ( .A1(n891), .A2(G138), .ZN(n544) );
  NAND2_X1 U605 ( .A1(G126), .A2(n884), .ZN(n541) );
  NAND2_X1 U606 ( .A1(G114), .A2(n885), .ZN(n540) );
  AND2_X1 U607 ( .A1(n541), .A2(n540), .ZN(n543) );
  NAND2_X1 U608 ( .A1(G102), .A2(n890), .ZN(n542) );
  NAND2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n681) );
  NOR2_X1 U610 ( .A1(n544), .A2(n681), .ZN(G164) );
  XOR2_X1 U611 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n546) );
  NAND2_X1 U612 ( .A1(G7), .A2(G661), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G223) );
  XOR2_X1 U614 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n548) );
  INV_X1 U615 ( .A(G223), .ZN(n826) );
  NAND2_X1 U616 ( .A1(G567), .A2(n826), .ZN(n547) );
  XNOR2_X1 U617 ( .A(n548), .B(n547), .ZN(G234) );
  NAND2_X1 U618 ( .A1(n638), .A2(G43), .ZN(n549) );
  XNOR2_X1 U619 ( .A(KEYINPUT74), .B(n549), .ZN(n559) );
  NAND2_X1 U620 ( .A1(n639), .A2(G56), .ZN(n550) );
  XNOR2_X1 U621 ( .A(KEYINPUT14), .B(n550), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n642), .A2(G81), .ZN(n551) );
  XNOR2_X1 U623 ( .A(n551), .B(KEYINPUT12), .ZN(n553) );
  NAND2_X1 U624 ( .A1(G68), .A2(n636), .ZN(n552) );
  NAND2_X1 U625 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U626 ( .A(KEYINPUT13), .B(n554), .ZN(n555) );
  NAND2_X1 U627 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U628 ( .A(KEYINPUT73), .B(n557), .ZN(n558) );
  NAND2_X1 U629 ( .A1(n559), .A2(n558), .ZN(n974) );
  INV_X1 U630 ( .A(G860), .ZN(n612) );
  OR2_X1 U631 ( .A1(n974), .A2(n612), .ZN(G153) );
  XNOR2_X1 U632 ( .A(G171), .B(KEYINPUT75), .ZN(G301) );
  NAND2_X1 U633 ( .A1(G868), .A2(G301), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n639), .A2(G66), .ZN(n566) );
  NAND2_X1 U635 ( .A1(G92), .A2(n642), .ZN(n561) );
  NAND2_X1 U636 ( .A1(G79), .A2(n636), .ZN(n560) );
  NAND2_X1 U637 ( .A1(n561), .A2(n560), .ZN(n564) );
  NAND2_X1 U638 ( .A1(n638), .A2(G54), .ZN(n562) );
  XOR2_X1 U639 ( .A(KEYINPUT76), .B(n562), .Z(n563) );
  NOR2_X1 U640 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U641 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U642 ( .A(KEYINPUT15), .B(n567), .Z(n966) );
  INV_X1 U643 ( .A(G868), .ZN(n595) );
  NAND2_X1 U644 ( .A1(n966), .A2(n595), .ZN(n568) );
  NAND2_X1 U645 ( .A1(n569), .A2(n568), .ZN(G284) );
  NAND2_X1 U646 ( .A1(G51), .A2(n638), .ZN(n571) );
  NAND2_X1 U647 ( .A1(G63), .A2(n639), .ZN(n570) );
  NAND2_X1 U648 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U649 ( .A(KEYINPUT6), .B(n572), .ZN(n579) );
  NAND2_X1 U650 ( .A1(n642), .A2(G89), .ZN(n573) );
  XNOR2_X1 U651 ( .A(n573), .B(KEYINPUT4), .ZN(n575) );
  NAND2_X1 U652 ( .A1(G76), .A2(n636), .ZN(n574) );
  NAND2_X1 U653 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U654 ( .A(KEYINPUT77), .B(n576), .ZN(n577) );
  XNOR2_X1 U655 ( .A(KEYINPUT5), .B(n577), .ZN(n578) );
  NOR2_X1 U656 ( .A1(n579), .A2(n578), .ZN(n581) );
  XOR2_X1 U657 ( .A(KEYINPUT7), .B(KEYINPUT78), .Z(n580) );
  XNOR2_X1 U658 ( .A(n581), .B(n580), .ZN(G168) );
  XOR2_X1 U659 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U660 ( .A1(G91), .A2(n642), .ZN(n583) );
  NAND2_X1 U661 ( .A1(G78), .A2(n636), .ZN(n582) );
  NAND2_X1 U662 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U663 ( .A(KEYINPUT70), .B(n584), .Z(n588) );
  NAND2_X1 U664 ( .A1(G53), .A2(n638), .ZN(n586) );
  NAND2_X1 U665 ( .A1(G65), .A2(n639), .ZN(n585) );
  AND2_X1 U666 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U667 ( .A1(n588), .A2(n587), .ZN(G299) );
  NOR2_X1 U668 ( .A1(G286), .A2(n595), .ZN(n589) );
  XOR2_X1 U669 ( .A(KEYINPUT79), .B(n589), .Z(n591) );
  NOR2_X1 U670 ( .A1(G868), .A2(G299), .ZN(n590) );
  NOR2_X1 U671 ( .A1(n591), .A2(n590), .ZN(G297) );
  NAND2_X1 U672 ( .A1(G559), .A2(n612), .ZN(n592) );
  XNOR2_X1 U673 ( .A(KEYINPUT80), .B(n592), .ZN(n593) );
  INV_X1 U674 ( .A(n966), .ZN(n610) );
  NAND2_X1 U675 ( .A1(n593), .A2(n610), .ZN(n594) );
  XNOR2_X1 U676 ( .A(KEYINPUT16), .B(n594), .ZN(G148) );
  NOR2_X1 U677 ( .A1(G559), .A2(n595), .ZN(n596) );
  NAND2_X1 U678 ( .A1(n610), .A2(n596), .ZN(n597) );
  XNOR2_X1 U679 ( .A(n597), .B(KEYINPUT81), .ZN(n599) );
  NOR2_X1 U680 ( .A1(n974), .A2(G868), .ZN(n598) );
  NOR2_X1 U681 ( .A1(n599), .A2(n598), .ZN(G282) );
  NAND2_X1 U682 ( .A1(G135), .A2(n891), .ZN(n600) );
  XNOR2_X1 U683 ( .A(n600), .B(KEYINPUT82), .ZN(n607) );
  NAND2_X1 U684 ( .A1(G99), .A2(n890), .ZN(n602) );
  NAND2_X1 U685 ( .A1(G111), .A2(n885), .ZN(n601) );
  NAND2_X1 U686 ( .A1(n602), .A2(n601), .ZN(n605) );
  NAND2_X1 U687 ( .A1(n884), .A2(G123), .ZN(n603) );
  XOR2_X1 U688 ( .A(KEYINPUT18), .B(n603), .Z(n604) );
  NOR2_X1 U689 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U690 ( .A1(n607), .A2(n606), .ZN(n923) );
  XOR2_X1 U691 ( .A(n923), .B(G2096), .Z(n609) );
  XNOR2_X1 U692 ( .A(G2100), .B(KEYINPUT83), .ZN(n608) );
  NAND2_X1 U693 ( .A1(n609), .A2(n608), .ZN(G156) );
  NAND2_X1 U694 ( .A1(G559), .A2(n610), .ZN(n611) );
  XOR2_X1 U695 ( .A(n974), .B(n611), .Z(n655) );
  NAND2_X1 U696 ( .A1(n612), .A2(n655), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G93), .A2(n642), .ZN(n614) );
  NAND2_X1 U698 ( .A1(G80), .A2(n636), .ZN(n613) );
  NAND2_X1 U699 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U700 ( .A(KEYINPUT84), .B(n615), .Z(n617) );
  NAND2_X1 U701 ( .A1(n639), .A2(G67), .ZN(n616) );
  NAND2_X1 U702 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U703 ( .A1(G55), .A2(n638), .ZN(n618) );
  XNOR2_X1 U704 ( .A(KEYINPUT85), .B(n618), .ZN(n619) );
  NOR2_X1 U705 ( .A1(n620), .A2(n619), .ZN(n657) );
  XOR2_X1 U706 ( .A(n621), .B(n657), .Z(G145) );
  NAND2_X1 U707 ( .A1(G87), .A2(n622), .ZN(n623) );
  XNOR2_X1 U708 ( .A(n623), .B(KEYINPUT86), .ZN(n628) );
  NAND2_X1 U709 ( .A1(G49), .A2(n638), .ZN(n625) );
  NAND2_X1 U710 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U711 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U712 ( .A1(n639), .A2(n626), .ZN(n627) );
  NAND2_X1 U713 ( .A1(n628), .A2(n627), .ZN(G288) );
  NAND2_X1 U714 ( .A1(G50), .A2(n638), .ZN(n630) );
  NAND2_X1 U715 ( .A1(G62), .A2(n639), .ZN(n629) );
  NAND2_X1 U716 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U717 ( .A1(G88), .A2(n642), .ZN(n632) );
  NAND2_X1 U718 ( .A1(G75), .A2(n636), .ZN(n631) );
  NAND2_X1 U719 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U720 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U721 ( .A(KEYINPUT88), .B(n635), .Z(G303) );
  NAND2_X1 U722 ( .A1(G73), .A2(n636), .ZN(n637) );
  XNOR2_X1 U723 ( .A(n637), .B(KEYINPUT2), .ZN(n647) );
  NAND2_X1 U724 ( .A1(G48), .A2(n638), .ZN(n641) );
  NAND2_X1 U725 ( .A1(G61), .A2(n639), .ZN(n640) );
  NAND2_X1 U726 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U727 ( .A1(G86), .A2(n642), .ZN(n643) );
  XNOR2_X1 U728 ( .A(KEYINPUT87), .B(n643), .ZN(n644) );
  NOR2_X1 U729 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U730 ( .A1(n647), .A2(n646), .ZN(G305) );
  XOR2_X1 U731 ( .A(KEYINPUT89), .B(KEYINPUT19), .Z(n648) );
  XNOR2_X1 U732 ( .A(G288), .B(n648), .ZN(n649) );
  XOR2_X1 U733 ( .A(n649), .B(n657), .Z(n651) );
  INV_X1 U734 ( .A(G299), .ZN(n967) );
  XNOR2_X1 U735 ( .A(n967), .B(G303), .ZN(n650) );
  XNOR2_X1 U736 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U737 ( .A(n652), .B(G305), .ZN(n653) );
  XNOR2_X1 U738 ( .A(n653), .B(G290), .ZN(n851) );
  XOR2_X1 U739 ( .A(n851), .B(KEYINPUT90), .Z(n654) );
  XNOR2_X1 U740 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U741 ( .A1(n656), .A2(G868), .ZN(n659) );
  OR2_X1 U742 ( .A1(G868), .A2(n657), .ZN(n658) );
  NAND2_X1 U743 ( .A1(n659), .A2(n658), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2084), .A2(G2078), .ZN(n660) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(n660), .Z(n661) );
  NAND2_X1 U746 ( .A1(G2090), .A2(n661), .ZN(n662) );
  XNOR2_X1 U747 ( .A(KEYINPUT21), .B(n662), .ZN(n663) );
  NAND2_X1 U748 ( .A1(n663), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U750 ( .A1(G483), .A2(G661), .ZN(n672) );
  NOR2_X1 U751 ( .A1(G235), .A2(G236), .ZN(n664) );
  NAND2_X1 U752 ( .A1(G108), .A2(n664), .ZN(n665) );
  NOR2_X1 U753 ( .A1(n665), .A2(G237), .ZN(n666) );
  XNOR2_X1 U754 ( .A(n666), .B(KEYINPUT91), .ZN(n830) );
  NAND2_X1 U755 ( .A1(n830), .A2(G567), .ZN(n671) );
  NOR2_X1 U756 ( .A1(G220), .A2(G219), .ZN(n667) );
  XOR2_X1 U757 ( .A(KEYINPUT22), .B(n667), .Z(n668) );
  NOR2_X1 U758 ( .A1(G218), .A2(n668), .ZN(n669) );
  NAND2_X1 U759 ( .A1(G96), .A2(n669), .ZN(n831) );
  NAND2_X1 U760 ( .A1(n831), .A2(G2106), .ZN(n670) );
  NAND2_X1 U761 ( .A1(n671), .A2(n670), .ZN(n832) );
  NOR2_X1 U762 ( .A1(n672), .A2(n832), .ZN(n673) );
  XNOR2_X1 U763 ( .A(n673), .B(KEYINPUT92), .ZN(n829) );
  NAND2_X1 U764 ( .A1(n829), .A2(G36), .ZN(n674) );
  XOR2_X1 U765 ( .A(KEYINPUT93), .B(n674), .Z(G176) );
  XNOR2_X1 U766 ( .A(G1986), .B(G290), .ZN(n959) );
  AND2_X1 U767 ( .A1(G40), .A2(n675), .ZN(n677) );
  AND2_X1 U768 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U769 ( .A1(n679), .A2(n678), .ZN(n690) );
  INV_X1 U770 ( .A(G1384), .ZN(n682) );
  AND2_X1 U771 ( .A1(G138), .A2(n682), .ZN(n680) );
  NAND2_X1 U772 ( .A1(n891), .A2(n680), .ZN(n684) );
  NAND2_X1 U773 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U774 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U775 ( .A(n685), .B(KEYINPUT65), .ZN(n689) );
  INV_X1 U776 ( .A(n689), .ZN(n686) );
  NOR2_X1 U777 ( .A1(n690), .A2(n686), .ZN(n687) );
  XOR2_X1 U778 ( .A(n687), .B(KEYINPUT94), .Z(n783) );
  INV_X1 U779 ( .A(n783), .ZN(n811) );
  NAND2_X1 U780 ( .A1(n959), .A2(n811), .ZN(n800) );
  XOR2_X1 U781 ( .A(KEYINPUT105), .B(G1981), .Z(n688) );
  XNOR2_X1 U782 ( .A(G305), .B(n688), .ZN(n978) );
  NOR2_X1 U783 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U784 ( .A1(n737), .A2(G8), .ZN(n762) );
  NOR2_X1 U785 ( .A1(G1976), .A2(G288), .ZN(n963) );
  NAND2_X1 U786 ( .A1(n963), .A2(KEYINPUT33), .ZN(n692) );
  NOR2_X1 U787 ( .A1(n762), .A2(n692), .ZN(n693) );
  XNOR2_X1 U788 ( .A(n693), .B(KEYINPUT104), .ZN(n694) );
  NOR2_X1 U789 ( .A1(n978), .A2(n694), .ZN(n757) );
  NAND2_X1 U790 ( .A1(n757), .A2(KEYINPUT33), .ZN(n751) );
  NOR2_X1 U791 ( .A1(G1966), .A2(n762), .ZN(n732) );
  XNOR2_X1 U792 ( .A(G2078), .B(KEYINPUT25), .ZN(n937) );
  NAND2_X1 U793 ( .A1(n709), .A2(n937), .ZN(n696) );
  INV_X1 U794 ( .A(G1961), .ZN(n984) );
  NAND2_X1 U795 ( .A1(n737), .A2(n984), .ZN(n695) );
  NAND2_X1 U796 ( .A1(n696), .A2(n695), .ZN(n726) );
  NAND2_X1 U797 ( .A1(n726), .A2(G171), .ZN(n722) );
  NAND2_X1 U798 ( .A1(G2072), .A2(n709), .ZN(n697) );
  XNOR2_X1 U799 ( .A(KEYINPUT27), .B(n697), .ZN(n701) );
  INV_X1 U800 ( .A(KEYINPUT101), .ZN(n699) );
  XOR2_X1 U801 ( .A(G1956), .B(KEYINPUT100), .Z(n985) );
  NOR2_X1 U802 ( .A1(n985), .A2(n709), .ZN(n698) );
  XNOR2_X1 U803 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U804 ( .A1(n701), .A2(n700), .ZN(n704) );
  XNOR2_X1 U805 ( .A(n703), .B(n702), .ZN(n720) );
  NAND2_X1 U806 ( .A1(n967), .A2(n704), .ZN(n718) );
  NAND2_X1 U807 ( .A1(n709), .A2(G1996), .ZN(n705) );
  XNOR2_X1 U808 ( .A(n705), .B(KEYINPUT26), .ZN(n707) );
  NAND2_X1 U809 ( .A1(n737), .A2(G1341), .ZN(n706) );
  NAND2_X1 U810 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U811 ( .A1(n974), .A2(n708), .ZN(n713) );
  NAND2_X1 U812 ( .A1(G2067), .A2(n709), .ZN(n711) );
  NAND2_X1 U813 ( .A1(n737), .A2(G1348), .ZN(n710) );
  NAND2_X1 U814 ( .A1(n711), .A2(n710), .ZN(n714) );
  NOR2_X1 U815 ( .A1(n966), .A2(n714), .ZN(n712) );
  OR2_X1 U816 ( .A1(n713), .A2(n712), .ZN(n716) );
  NAND2_X1 U817 ( .A1(n966), .A2(n714), .ZN(n715) );
  NAND2_X1 U818 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U819 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U820 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U821 ( .A1(n722), .A2(n514), .ZN(n731) );
  NOR2_X1 U822 ( .A1(n737), .A2(G2084), .ZN(n733) );
  NOR2_X1 U823 ( .A1(n732), .A2(n733), .ZN(n723) );
  NAND2_X1 U824 ( .A1(G8), .A2(n723), .ZN(n724) );
  XNOR2_X1 U825 ( .A(KEYINPUT30), .B(n724), .ZN(n725) );
  NOR2_X1 U826 ( .A1(G168), .A2(n725), .ZN(n728) );
  NOR2_X1 U827 ( .A1(G171), .A2(n726), .ZN(n727) );
  NOR2_X1 U828 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U829 ( .A(KEYINPUT31), .B(n729), .Z(n730) );
  NAND2_X1 U830 ( .A1(n731), .A2(n730), .ZN(n736) );
  NOR2_X1 U831 ( .A1(n732), .A2(n513), .ZN(n735) );
  NAND2_X1 U832 ( .A1(G8), .A2(n733), .ZN(n734) );
  NAND2_X1 U833 ( .A1(n735), .A2(n734), .ZN(n746) );
  NAND2_X1 U834 ( .A1(n736), .A2(G286), .ZN(n742) );
  NOR2_X1 U835 ( .A1(G1971), .A2(n762), .ZN(n739) );
  NOR2_X1 U836 ( .A1(n737), .A2(G2090), .ZN(n738) );
  NOR2_X1 U837 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U838 ( .A1(G303), .A2(n740), .ZN(n741) );
  NAND2_X1 U839 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U840 ( .A1(n743), .A2(G8), .ZN(n744) );
  XNOR2_X1 U841 ( .A(KEYINPUT32), .B(n744), .ZN(n745) );
  NAND2_X1 U842 ( .A1(n746), .A2(n745), .ZN(n755) );
  NOR2_X1 U843 ( .A1(G2090), .A2(G303), .ZN(n747) );
  NAND2_X1 U844 ( .A1(G8), .A2(n747), .ZN(n748) );
  NAND2_X1 U845 ( .A1(n755), .A2(n748), .ZN(n749) );
  NAND2_X1 U846 ( .A1(n749), .A2(n762), .ZN(n750) );
  NAND2_X1 U847 ( .A1(n751), .A2(n750), .ZN(n765) );
  NOR2_X1 U848 ( .A1(G1981), .A2(G305), .ZN(n752) );
  XNOR2_X1 U849 ( .A(KEYINPUT24), .B(n752), .ZN(n761) );
  NOR2_X1 U850 ( .A1(G303), .A2(G1971), .ZN(n753) );
  NOR2_X1 U851 ( .A1(n963), .A2(n753), .ZN(n754) );
  NAND2_X1 U852 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n958) );
  NAND2_X1 U854 ( .A1(n757), .A2(n958), .ZN(n758) );
  NOR2_X1 U855 ( .A1(n761), .A2(n760), .ZN(n763) );
  NOR2_X1 U856 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U857 ( .A1(n765), .A2(n764), .ZN(n798) );
  NAND2_X1 U858 ( .A1(G119), .A2(n884), .ZN(n767) );
  NAND2_X1 U859 ( .A1(G107), .A2(n885), .ZN(n766) );
  NAND2_X1 U860 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U861 ( .A(KEYINPUT98), .B(n768), .ZN(n772) );
  NAND2_X1 U862 ( .A1(G95), .A2(n890), .ZN(n770) );
  NAND2_X1 U863 ( .A1(G131), .A2(n891), .ZN(n769) );
  NAND2_X1 U864 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n881) );
  INV_X1 U866 ( .A(G1991), .ZN(n942) );
  NOR2_X1 U867 ( .A1(n881), .A2(n942), .ZN(n782) );
  NAND2_X1 U868 ( .A1(G105), .A2(n890), .ZN(n773) );
  XNOR2_X1 U869 ( .A(n773), .B(KEYINPUT38), .ZN(n780) );
  NAND2_X1 U870 ( .A1(G117), .A2(n885), .ZN(n775) );
  NAND2_X1 U871 ( .A1(G141), .A2(n891), .ZN(n774) );
  NAND2_X1 U872 ( .A1(n775), .A2(n774), .ZN(n778) );
  NAND2_X1 U873 ( .A1(G129), .A2(n884), .ZN(n776) );
  XNOR2_X1 U874 ( .A(KEYINPUT99), .B(n776), .ZN(n777) );
  NOR2_X1 U875 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U876 ( .A1(n780), .A2(n779), .ZN(n875) );
  AND2_X1 U877 ( .A1(G1996), .A2(n875), .ZN(n781) );
  NOR2_X1 U878 ( .A1(n782), .A2(n781), .ZN(n911) );
  NOR2_X1 U879 ( .A1(n911), .A2(n783), .ZN(n804) );
  INV_X1 U880 ( .A(n804), .ZN(n796) );
  NAND2_X1 U881 ( .A1(G104), .A2(n890), .ZN(n785) );
  NAND2_X1 U882 ( .A1(G140), .A2(n891), .ZN(n784) );
  NAND2_X1 U883 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U884 ( .A(KEYINPUT34), .B(n786), .ZN(n792) );
  NAND2_X1 U885 ( .A1(n885), .A2(G116), .ZN(n787) );
  XOR2_X1 U886 ( .A(KEYINPUT95), .B(n787), .Z(n789) );
  NAND2_X1 U887 ( .A1(n884), .A2(G128), .ZN(n788) );
  NAND2_X1 U888 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U889 ( .A(n790), .B(KEYINPUT35), .Z(n791) );
  NOR2_X1 U890 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U891 ( .A(KEYINPUT36), .B(n793), .Z(n794) );
  XOR2_X1 U892 ( .A(KEYINPUT96), .B(n794), .Z(n880) );
  XNOR2_X1 U893 ( .A(G2067), .B(KEYINPUT37), .ZN(n809) );
  OR2_X1 U894 ( .A1(n880), .A2(n809), .ZN(n795) );
  XNOR2_X1 U895 ( .A(n795), .B(KEYINPUT97), .ZN(n927) );
  NAND2_X1 U896 ( .A1(n927), .A2(n811), .ZN(n807) );
  NAND2_X1 U897 ( .A1(n796), .A2(n807), .ZN(n797) );
  NOR2_X1 U898 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U899 ( .A1(n800), .A2(n799), .ZN(n814) );
  NOR2_X1 U900 ( .A1(G1996), .A2(n875), .ZN(n908) );
  AND2_X1 U901 ( .A1(n942), .A2(n881), .ZN(n922) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n801) );
  XNOR2_X1 U903 ( .A(KEYINPUT106), .B(n801), .ZN(n802) );
  NOR2_X1 U904 ( .A1(n922), .A2(n802), .ZN(n803) );
  NOR2_X1 U905 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U906 ( .A1(n908), .A2(n805), .ZN(n806) );
  XNOR2_X1 U907 ( .A(n806), .B(KEYINPUT39), .ZN(n808) );
  NAND2_X1 U908 ( .A1(n808), .A2(n807), .ZN(n810) );
  NAND2_X1 U909 ( .A1(n880), .A2(n809), .ZN(n919) );
  NAND2_X1 U910 ( .A1(n810), .A2(n919), .ZN(n812) );
  NAND2_X1 U911 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U912 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U913 ( .A(KEYINPUT40), .B(n815), .ZN(G329) );
  XOR2_X1 U914 ( .A(G2454), .B(G2430), .Z(n817) );
  XNOR2_X1 U915 ( .A(G2451), .B(G2446), .ZN(n816) );
  XNOR2_X1 U916 ( .A(n817), .B(n816), .ZN(n824) );
  XOR2_X1 U917 ( .A(G2443), .B(G2427), .Z(n819) );
  XNOR2_X1 U918 ( .A(G2438), .B(KEYINPUT107), .ZN(n818) );
  XNOR2_X1 U919 ( .A(n819), .B(n818), .ZN(n820) );
  XOR2_X1 U920 ( .A(n820), .B(G2435), .Z(n822) );
  XNOR2_X1 U921 ( .A(G1341), .B(G1348), .ZN(n821) );
  XNOR2_X1 U922 ( .A(n822), .B(n821), .ZN(n823) );
  XNOR2_X1 U923 ( .A(n824), .B(n823), .ZN(n825) );
  NAND2_X1 U924 ( .A1(n825), .A2(G14), .ZN(n901) );
  XOR2_X1 U925 ( .A(KEYINPUT108), .B(n901), .Z(G401) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n826), .ZN(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U928 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U930 ( .A1(n829), .A2(n828), .ZN(G188) );
  NOR2_X1 U931 ( .A1(n831), .A2(n830), .ZN(G325) );
  XNOR2_X1 U932 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  XNOR2_X1 U933 ( .A(G108), .B(KEYINPUT117), .ZN(G238) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  INV_X1 U936 ( .A(n832), .ZN(G319) );
  XOR2_X1 U937 ( .A(G1981), .B(G1956), .Z(n834) );
  XNOR2_X1 U938 ( .A(G1966), .B(G1961), .ZN(n833) );
  XNOR2_X1 U939 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U940 ( .A(n835), .B(G2474), .Z(n837) );
  XNOR2_X1 U941 ( .A(G1996), .B(G1991), .ZN(n836) );
  XNOR2_X1 U942 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U943 ( .A(KEYINPUT41), .B(G1986), .Z(n839) );
  XNOR2_X1 U944 ( .A(G1971), .B(G1976), .ZN(n838) );
  XNOR2_X1 U945 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U946 ( .A(n841), .B(n840), .ZN(G229) );
  XOR2_X1 U947 ( .A(G2096), .B(KEYINPUT110), .Z(n843) );
  XNOR2_X1 U948 ( .A(G2067), .B(KEYINPUT43), .ZN(n842) );
  XNOR2_X1 U949 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U950 ( .A(n844), .B(KEYINPUT42), .Z(n846) );
  XNOR2_X1 U951 ( .A(G2072), .B(G2090), .ZN(n845) );
  XNOR2_X1 U952 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U953 ( .A(G2678), .B(G2100), .Z(n848) );
  XNOR2_X1 U954 ( .A(G2084), .B(G2078), .ZN(n847) );
  XNOR2_X1 U955 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U956 ( .A(n850), .B(n849), .ZN(G227) );
  XNOR2_X1 U957 ( .A(n851), .B(G286), .ZN(n854) );
  XNOR2_X1 U958 ( .A(G171), .B(KEYINPUT115), .ZN(n852) );
  XNOR2_X1 U959 ( .A(n852), .B(n966), .ZN(n853) );
  XNOR2_X1 U960 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U961 ( .A(n855), .B(n974), .Z(n856) );
  NOR2_X1 U962 ( .A1(G37), .A2(n856), .ZN(n857) );
  XNOR2_X1 U963 ( .A(KEYINPUT116), .B(n857), .ZN(G397) );
  NAND2_X1 U964 ( .A1(n884), .A2(G124), .ZN(n858) );
  XNOR2_X1 U965 ( .A(n858), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U966 ( .A1(G112), .A2(n885), .ZN(n859) );
  NAND2_X1 U967 ( .A1(n860), .A2(n859), .ZN(n864) );
  NAND2_X1 U968 ( .A1(G100), .A2(n890), .ZN(n862) );
  NAND2_X1 U969 ( .A1(G136), .A2(n891), .ZN(n861) );
  NAND2_X1 U970 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U971 ( .A1(n864), .A2(n863), .ZN(G162) );
  NAND2_X1 U972 ( .A1(G130), .A2(n884), .ZN(n866) );
  NAND2_X1 U973 ( .A1(G118), .A2(n885), .ZN(n865) );
  NAND2_X1 U974 ( .A1(n866), .A2(n865), .ZN(n871) );
  NAND2_X1 U975 ( .A1(G106), .A2(n890), .ZN(n868) );
  NAND2_X1 U976 ( .A1(G142), .A2(n891), .ZN(n867) );
  NAND2_X1 U977 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U978 ( .A(n869), .B(KEYINPUT45), .Z(n870) );
  NOR2_X1 U979 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U980 ( .A(n872), .B(n923), .ZN(n879) );
  XNOR2_X1 U981 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n873) );
  XNOR2_X1 U982 ( .A(n873), .B(KEYINPUT46), .ZN(n874) );
  XOR2_X1 U983 ( .A(n874), .B(G162), .Z(n877) );
  XOR2_X1 U984 ( .A(G164), .B(n875), .Z(n876) );
  XNOR2_X1 U985 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U986 ( .A(n879), .B(n878), .Z(n883) );
  XNOR2_X1 U987 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U988 ( .A(n883), .B(n882), .ZN(n898) );
  NAND2_X1 U989 ( .A1(G127), .A2(n884), .ZN(n887) );
  NAND2_X1 U990 ( .A1(G115), .A2(n885), .ZN(n886) );
  NAND2_X1 U991 ( .A1(n887), .A2(n886), .ZN(n889) );
  XOR2_X1 U992 ( .A(KEYINPUT112), .B(KEYINPUT47), .Z(n888) );
  XNOR2_X1 U993 ( .A(n889), .B(n888), .ZN(n896) );
  NAND2_X1 U994 ( .A1(G103), .A2(n890), .ZN(n893) );
  NAND2_X1 U995 ( .A1(G139), .A2(n891), .ZN(n892) );
  NAND2_X1 U996 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U997 ( .A(KEYINPUT111), .B(n894), .Z(n895) );
  NOR2_X1 U998 ( .A1(n896), .A2(n895), .ZN(n912) );
  XNOR2_X1 U999 ( .A(n912), .B(G160), .ZN(n897) );
  XNOR2_X1 U1000 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n899), .ZN(n900) );
  XNOR2_X1 U1002 ( .A(KEYINPUT114), .B(n900), .ZN(G395) );
  NAND2_X1 U1003 ( .A1(G319), .A2(n901), .ZN(n904) );
  NOR2_X1 U1004 ( .A1(G229), .A2(G227), .ZN(n902) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n902), .ZN(n903) );
  NOR2_X1 U1006 ( .A1(n904), .A2(n903), .ZN(n906) );
  NOR2_X1 U1007 ( .A1(G397), .A2(G395), .ZN(n905) );
  NAND2_X1 U1008 ( .A1(n906), .A2(n905), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(G303), .ZN(G166) );
  XOR2_X1 U1011 ( .A(G2090), .B(G162), .Z(n907) );
  NOR2_X1 U1012 ( .A1(n908), .A2(n907), .ZN(n909) );
  XOR2_X1 U1013 ( .A(KEYINPUT51), .B(n909), .Z(n910) );
  NAND2_X1 U1014 ( .A1(n911), .A2(n910), .ZN(n918) );
  XOR2_X1 U1015 ( .A(G2072), .B(n912), .Z(n914) );
  XOR2_X1 U1016 ( .A(G164), .B(G2078), .Z(n913) );
  NOR2_X1 U1017 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1018 ( .A(KEYINPUT50), .B(n915), .Z(n916) );
  XNOR2_X1 U1019 ( .A(KEYINPUT120), .B(n916), .ZN(n917) );
  NOR2_X1 U1020 ( .A1(n918), .A2(n917), .ZN(n920) );
  NAND2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n930) );
  XOR2_X1 U1022 ( .A(G2084), .B(G160), .Z(n921) );
  NOR2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n924) );
  NAND2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(KEYINPUT118), .B(n925), .ZN(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(KEYINPUT119), .B(n928), .ZN(n929) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(KEYINPUT52), .B(n931), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n954) );
  NAND2_X1 U1031 ( .A1(n932), .A2(n954), .ZN(n933) );
  NAND2_X1 U1032 ( .A1(n933), .A2(G29), .ZN(n1015) );
  XNOR2_X1 U1033 ( .A(G2084), .B(G34), .ZN(n934) );
  XNOR2_X1 U1034 ( .A(n934), .B(KEYINPUT54), .ZN(n949) );
  XNOR2_X1 U1035 ( .A(G1996), .B(G32), .ZN(n936) );
  XNOR2_X1 U1036 ( .A(G2072), .B(G33), .ZN(n935) );
  NOR2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n941) );
  XOR2_X1 U1038 ( .A(n937), .B(G27), .Z(n939) );
  XNOR2_X1 U1039 ( .A(G2067), .B(G26), .ZN(n938) );
  NOR2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1041 ( .A1(n941), .A2(n940), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(G25), .B(n942), .ZN(n943) );
  NAND2_X1 U1043 ( .A1(n943), .A2(G28), .ZN(n944) );
  XOR2_X1 U1044 ( .A(KEYINPUT123), .B(n944), .Z(n945) );
  NOR2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1046 ( .A(n947), .B(KEYINPUT53), .ZN(n948) );
  NOR2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n952) );
  XOR2_X1 U1048 ( .A(G2090), .B(KEYINPUT122), .Z(n950) );
  XNOR2_X1 U1049 ( .A(G35), .B(n950), .ZN(n951) );
  NAND2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(n954), .B(n953), .ZN(n956) );
  INV_X1 U1052 ( .A(G29), .ZN(n955) );
  NAND2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1054 ( .A1(G11), .A2(n957), .ZN(n1013) );
  XNOR2_X1 U1055 ( .A(KEYINPUT56), .B(G16), .ZN(n983) );
  XNOR2_X1 U1056 ( .A(G1971), .B(G166), .ZN(n962) );
  INV_X1 U1057 ( .A(n958), .ZN(n960) );
  NOR2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(KEYINPUT124), .B(n963), .ZN(n964) );
  NOR2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n973) );
  XOR2_X1 U1062 ( .A(n966), .B(G1348), .Z(n969) );
  XNOR2_X1 U1063 ( .A(n967), .B(G1956), .ZN(n968) );
  NAND2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n971) );
  XOR2_X1 U1065 ( .A(G171), .B(G1961), .Z(n970) );
  NOR2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(G1341), .B(n974), .ZN(n975) );
  NOR2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n981) );
  XOR2_X1 U1070 ( .A(G168), .B(G1966), .Z(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1072 ( .A(KEYINPUT57), .B(n979), .Z(n980) );
  NAND2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n1011) );
  XNOR2_X1 U1075 ( .A(G5), .B(n984), .ZN(n1004) );
  XNOR2_X1 U1076 ( .A(n985), .B(G20), .ZN(n993) );
  XOR2_X1 U1077 ( .A(G1981), .B(G6), .Z(n988) );
  XOR2_X1 U1078 ( .A(G19), .B(KEYINPUT126), .Z(n986) );
  XNOR2_X1 U1079 ( .A(G1341), .B(n986), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n991) );
  XOR2_X1 U1081 ( .A(KEYINPUT59), .B(G1348), .Z(n989) );
  XNOR2_X1 U1082 ( .A(G4), .B(n989), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(n994), .B(KEYINPUT60), .ZN(n1002) );
  XNOR2_X1 U1086 ( .A(G1971), .B(G22), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(G1986), .B(G24), .ZN(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(G1976), .B(KEYINPUT127), .ZN(n997) );
  XNOR2_X1 U1090 ( .A(n997), .B(G23), .ZN(n998) );
  NAND2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1092 ( .A(KEYINPUT58), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(G21), .B(G1966), .ZN(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(n1007), .B(KEYINPUT61), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(G16), .B(KEYINPUT125), .ZN(n1008) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(KEYINPUT62), .B(n1016), .Z(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

