//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT68), .B1(new_n189), .B2(G116), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT68), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G119), .ZN(new_n193));
  AOI22_X1  g007(.A1(new_n190), .A2(new_n193), .B1(G116), .B2(new_n189), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n196));
  INV_X1    g010(.A(G113), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n199));
  AOI22_X1  g013(.A1(new_n198), .A2(new_n199), .B1(KEYINPUT2), .B2(G113), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT69), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n194), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n201), .B1(new_n194), .B2(new_n200), .ZN(new_n204));
  OAI22_X1  g018(.A1(new_n203), .A2(new_n204), .B1(new_n200), .B2(new_n194), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT30), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G128), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT0), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G128), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n218), .B1(new_n207), .B2(G146), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n209), .A2(KEYINPUT64), .A3(G143), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G128), .A4(new_n208), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n217), .B1(new_n221), .B2(new_n214), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT70), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT11), .ZN(new_n225));
  INV_X1    g039(.A(G134), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(G137), .ZN(new_n227));
  INV_X1    g041(.A(G137), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT11), .A3(G134), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n226), .A2(G137), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G131), .ZN(new_n232));
  INV_X1    g046(.A(G131), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n227), .A2(new_n229), .A3(new_n233), .A4(new_n230), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n217), .B(KEYINPUT70), .C1(new_n221), .C2(new_n214), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n224), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n226), .A2(G137), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n228), .A2(G134), .ZN(new_n239));
  OAI21_X1  g053(.A(G131), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n211), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n210), .ZN(new_n248));
  OR2_X1    g062(.A1(KEYINPUT66), .A2(G128), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT66), .A2(G128), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n242), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n221), .A2(new_n247), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n241), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n206), .B1(new_n237), .B2(new_n254), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n219), .A2(new_n208), .A3(new_n220), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(KEYINPUT0), .A3(G128), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n235), .A2(new_n257), .A3(new_n217), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n254), .A2(new_n258), .A3(new_n206), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n205), .B1(new_n255), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n205), .A2(new_n261), .ZN(new_n262));
  OAI221_X1 g076(.A(KEYINPUT71), .B1(new_n200), .B2(new_n194), .C1(new_n203), .C2(new_n204), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n262), .A2(new_n263), .A3(new_n237), .A4(new_n254), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT72), .B(G237), .ZN(new_n265));
  INV_X1    g079(.A(G953), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(G210), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n267), .B(KEYINPUT27), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT26), .B(G101), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n260), .A2(KEYINPUT73), .A3(new_n264), .A4(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(KEYINPUT31), .ZN(new_n272));
  XOR2_X1   g086(.A(new_n270), .B(KEYINPUT74), .Z(new_n273));
  NAND2_X1  g087(.A1(new_n254), .A2(new_n258), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n205), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT75), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n205), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n264), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT28), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT28), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n264), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n273), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n187), .B(new_n188), .C1(new_n272), .C2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT76), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT32), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT31), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n271), .B(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n280), .A2(new_n282), .ZN(new_n290));
  INV_X1    g104(.A(new_n273), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n293), .A2(KEYINPUT76), .A3(new_n187), .A4(new_n188), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n286), .A2(new_n287), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n284), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT32), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n280), .A2(new_n273), .A3(new_n282), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT29), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n260), .A2(new_n264), .ZN(new_n300));
  INV_X1    g114(.A(new_n270), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n298), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT77), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n298), .A2(KEYINPUT77), .A3(new_n299), .A4(new_n302), .ZN(new_n306));
  INV_X1    g120(.A(new_n282), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n262), .A2(new_n263), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n237), .A2(new_n254), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n264), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n307), .B1(KEYINPUT28), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n301), .A2(new_n299), .ZN(new_n313));
  AOI21_X1  g127(.A(G902), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n305), .A2(new_n306), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G472), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n295), .A2(new_n297), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G110), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT23), .B1(new_n212), .B2(G119), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n319), .B1(new_n189), .B2(G128), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n249), .A2(KEYINPUT23), .A3(G119), .A4(new_n250), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OR2_X1    g136(.A1(new_n322), .A2(KEYINPUT78), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(KEYINPUT78), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n318), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT16), .ZN(new_n326));
  INV_X1    g140(.A(G140), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(G125), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(G125), .ZN(new_n329));
  INV_X1    g143(.A(G125), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G140), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n328), .B1(new_n332), .B2(new_n326), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n209), .ZN(new_n334));
  OAI211_X1 g148(.A(G146), .B(new_n328), .C1(new_n332), .C2(new_n326), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n249), .A2(new_n250), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G119), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n189), .A2(G128), .ZN(new_n339));
  XOR2_X1   g153(.A(KEYINPUT24), .B(G110), .Z(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  OR2_X1    g156(.A1(new_n325), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n329), .A2(new_n331), .A3(new_n209), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n340), .B1(new_n338), .B2(new_n339), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n322), .A2(G110), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n335), .B(new_n345), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n343), .A2(new_n344), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n266), .A2(G221), .A3(G234), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(KEYINPUT79), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT22), .B(G137), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n351), .B(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n348), .B1(new_n325), .B2(new_n342), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n353), .B1(new_n354), .B2(KEYINPUT80), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n343), .A2(new_n344), .A3(new_n353), .A4(new_n348), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G217), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n359), .B1(G234), .B2(new_n188), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(G902), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT25), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n358), .A2(new_n363), .A3(new_n188), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n360), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n363), .B1(new_n358), .B2(new_n188), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n362), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT94), .ZN(new_n369));
  AND2_X1   g183(.A1(KEYINPUT72), .A2(G237), .ZN(new_n370));
  NOR2_X1   g184(.A1(KEYINPUT72), .A2(G237), .ZN(new_n371));
  OAI211_X1 g185(.A(G214), .B(new_n266), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n207), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n265), .A2(G143), .A3(G214), .A4(new_n266), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n233), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT18), .ZN(new_n376));
  NAND2_X1  g190(.A1(KEYINPUT18), .A2(G131), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n373), .A2(new_n374), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT90), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n209), .B1(new_n329), .B2(new_n331), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(new_n345), .A3(KEYINPUT89), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT89), .ZN(new_n384));
  INV_X1    g198(.A(new_n345), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n384), .B1(new_n385), .B2(new_n381), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT90), .A4(new_n377), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n376), .A2(new_n380), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT91), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n375), .A2(KEYINPUT18), .B1(new_n383), .B2(new_n386), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT91), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n391), .A2(new_n392), .A3(new_n380), .A4(new_n388), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(G113), .B(G122), .ZN(new_n395));
  INV_X1    g209(.A(G104), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n395), .B(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n336), .B1(KEYINPUT17), .B2(new_n375), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n373), .A2(new_n374), .A3(new_n233), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n399), .A2(new_n375), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n398), .B1(new_n400), .B2(KEYINPUT17), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n394), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n335), .ZN(new_n403));
  AOI21_X1  g217(.A(KEYINPUT93), .B1(new_n332), .B2(KEYINPUT19), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n332), .A2(new_n405), .ZN(new_n406));
  MUX2_X1   g220(.A(new_n404), .B(KEYINPUT93), .S(new_n406), .Z(new_n407));
  AOI21_X1  g221(.A(new_n403), .B1(new_n407), .B2(new_n209), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n400), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n397), .B1(new_n394), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n369), .B1(new_n402), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(G475), .A2(G902), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n394), .A2(new_n397), .A3(new_n401), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n390), .A2(new_n393), .B1(new_n408), .B2(new_n400), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n413), .B(KEYINPUT94), .C1(new_n397), .C2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT20), .ZN(new_n417));
  NOR3_X1   g231(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n418), .B1(new_n402), .B2(new_n410), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n394), .A2(new_n401), .ZN(new_n421));
  INV_X1    g235(.A(new_n397), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(G902), .B1(new_n423), .B2(new_n413), .ZN(new_n424));
  INV_X1    g238(.A(G475), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n212), .A2(G143), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n428), .B1(new_n337), .B2(G143), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n429), .A2(new_n226), .ZN(new_n430));
  INV_X1    g244(.A(new_n428), .ZN(new_n431));
  OAI21_X1  g245(.A(G134), .B1(new_n431), .B2(KEYINPUT13), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n432), .B1(new_n429), .B2(KEYINPUT13), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n192), .A2(G122), .ZN(new_n434));
  INV_X1    g248(.A(G122), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(G116), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(G107), .ZN(new_n438));
  OR3_X1    g252(.A1(new_n430), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G107), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n429), .A2(new_n226), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n441), .B1(new_n430), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n434), .A2(KEYINPUT14), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT95), .B1(new_n444), .B2(new_n436), .ZN(new_n445));
  INV_X1    g259(.A(new_n436), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n445), .B1(KEYINPUT14), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT14), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n436), .A2(KEYINPUT95), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n440), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n439), .B1(new_n443), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT9), .B(G234), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n452), .A2(new_n359), .A3(G953), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n439), .B(new_n453), .C1(new_n443), .C2(new_n450), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT15), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G478), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(new_n188), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n459), .B1(new_n457), .B2(new_n188), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n266), .A2(G952), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(G234), .B2(G237), .ZN(new_n465));
  XOR2_X1   g279(.A(KEYINPUT21), .B(G898), .Z(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT96), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(G234), .A2(G237), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(G902), .A3(G953), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n465), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n420), .A2(new_n427), .A3(new_n463), .A4(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(G214), .B1(G237), .B2(G902), .ZN(new_n476));
  XOR2_X1   g290(.A(new_n476), .B(KEYINPUT84), .Z(new_n477));
  OR2_X1    g291(.A1(new_n221), .A2(new_n247), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n245), .A2(new_n246), .B1(G143), .B2(new_n209), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n211), .B1(new_n479), .B2(new_n337), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(new_n330), .A3(new_n480), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n481), .A2(KEYINPUT86), .B1(G125), .B2(new_n222), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n222), .A2(G125), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT86), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G224), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(G953), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n483), .A2(KEYINPUT7), .A3(new_n487), .A4(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT3), .B1(new_n396), .B2(G107), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT3), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(new_n440), .A3(G104), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n396), .A2(G107), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(G101), .ZN(new_n497));
  INV_X1    g311(.A(G101), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n492), .A2(new_n494), .A3(new_n498), .A4(new_n495), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(KEYINPUT4), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT4), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n496), .A2(new_n501), .A3(G101), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n205), .A2(new_n503), .ZN(new_n504));
  OR3_X1    g318(.A1(new_n192), .A2(KEYINPUT5), .A3(G119), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G113), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n506), .B1(new_n194), .B2(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n194), .A2(new_n200), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT69), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n507), .B1(new_n509), .B2(new_n202), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n440), .A2(G104), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n396), .A2(G107), .ZN(new_n512));
  OAI21_X1  g326(.A(G101), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n499), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT82), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n499), .A2(new_n513), .A3(KEYINPUT82), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(G110), .B(G122), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n504), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n490), .A2(KEYINPUT7), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n482), .B2(new_n486), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n491), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n203), .A2(new_n204), .ZN(new_n525));
  OAI211_X1 g339(.A(KEYINPUT87), .B(new_n514), .C1(new_n525), .C2(new_n507), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT87), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n499), .A2(new_n513), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n527), .B1(new_n510), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n526), .A2(new_n529), .A3(new_n519), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n520), .B(KEYINPUT8), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n530), .A2(KEYINPUT88), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT88), .B1(new_n530), .B2(new_n531), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n524), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n483), .A2(new_n487), .A3(new_n490), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n489), .B1(new_n482), .B2(new_n486), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n504), .A2(new_n519), .ZN(new_n538));
  INV_X1    g352(.A(new_n520), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(KEYINPUT6), .A3(new_n521), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n520), .B1(new_n504), .B2(new_n519), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT85), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT6), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n543), .B1(new_n542), .B2(new_n544), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n537), .B(new_n541), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n534), .A2(new_n547), .A3(new_n188), .ZN(new_n548));
  OAI21_X1  g362(.A(G210), .B1(G237), .B2(G902), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n534), .A2(new_n547), .A3(new_n188), .A4(new_n549), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n477), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(G221), .B1(new_n452), .B2(G902), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n554), .B(KEYINPUT81), .Z(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G469), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n224), .A2(new_n236), .A3(new_n502), .A4(new_n500), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n247), .A2(new_n210), .B1(new_n249), .B2(new_n250), .ZN(new_n559));
  OAI22_X1  g373(.A1(new_n559), .A2(new_n242), .B1(new_n221), .B2(new_n247), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT82), .B1(new_n499), .B2(new_n513), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n499), .A2(new_n513), .A3(KEYINPUT82), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n560), .B(KEYINPUT10), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n212), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n564));
  OAI22_X1  g378(.A1(new_n256), .A2(new_n564), .B1(new_n221), .B2(new_n247), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n528), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT10), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n235), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n558), .A2(new_n563), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(G110), .B(G140), .ZN(new_n571));
  INV_X1    g385(.A(G227), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(G953), .ZN(new_n573));
  XOR2_X1   g387(.A(new_n571), .B(new_n573), .Z(new_n574));
  NAND2_X1  g388(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n516), .A2(new_n480), .A3(new_n478), .A4(new_n517), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n566), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT12), .B1(new_n577), .B2(new_n235), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT12), .ZN(new_n580));
  AOI211_X1 g394(.A(new_n580), .B(new_n569), .C1(new_n576), .C2(new_n566), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n575), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n558), .A2(new_n563), .A3(new_n568), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n235), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n574), .B1(new_n585), .B2(new_n570), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n557), .B(new_n188), .C1(new_n583), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT83), .ZN(new_n588));
  INV_X1    g402(.A(new_n574), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n567), .B1(new_n478), .B2(new_n480), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n590), .A2(new_n518), .B1(new_n566), .B2(new_n567), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n569), .B1(new_n591), .B2(new_n558), .ZN(new_n592));
  AND4_X1   g406(.A1(new_n569), .A2(new_n558), .A3(new_n563), .A4(new_n568), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n589), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n574), .B(new_n570), .C1(new_n578), .C2(new_n581), .ZN(new_n595));
  AOI21_X1  g409(.A(G902), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT83), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n597), .A3(new_n557), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n588), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(G469), .A2(G902), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n570), .B1(new_n578), .B2(new_n581), .ZN(new_n601));
  INV_X1    g415(.A(new_n575), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n601), .A2(new_n589), .B1(new_n602), .B2(new_n585), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(G469), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n599), .A2(new_n600), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n553), .A2(new_n556), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n317), .A2(new_n368), .A3(new_n475), .A4(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G101), .ZN(G3));
  NAND2_X1  g423(.A1(new_n553), .A2(new_n473), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n457), .A2(new_n188), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(G478), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n457), .A2(KEYINPUT33), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n455), .B2(new_n456), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n188), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n612), .B1(new_n616), .B2(G478), .ZN(new_n617));
  INV_X1    g431(.A(new_n419), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n416), .B2(KEYINPUT20), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n617), .B1(new_n619), .B2(new_n426), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n610), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n188), .B1(new_n272), .B2(new_n283), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(G472), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n286), .A2(new_n294), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n368), .A2(new_n605), .A3(new_n556), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n621), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT97), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT34), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT98), .B(G104), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  NAND3_X1  g445(.A1(new_n411), .A2(new_n415), .A3(new_n418), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(KEYINPUT99), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n411), .A2(new_n634), .A3(new_n415), .A4(new_n418), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n417), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n463), .A2(new_n426), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n610), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(new_n625), .A3(new_n626), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  NOR2_X1   g456(.A1(new_n353), .A2(KEYINPUT36), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n354), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n361), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n645), .B1(new_n365), .B2(new_n366), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n607), .A2(new_n625), .A3(new_n475), .A4(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT37), .B(G110), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G12));
  NAND2_X1  g463(.A1(new_n553), .A2(new_n646), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n465), .B(KEYINPUT100), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n651), .B1(G900), .B2(new_n470), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n650), .A2(new_n638), .A3(new_n653), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n605), .A2(new_n556), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n317), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  XNOR2_X1  g471(.A(new_n652), .B(KEYINPUT39), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n291), .A2(KEYINPUT101), .A3(new_n311), .ZN(new_n662));
  AOI21_X1  g476(.A(KEYINPUT101), .B1(new_n291), .B2(new_n311), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n300), .A2(new_n301), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(G472), .B1(new_n665), .B2(G902), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n295), .A2(new_n666), .A3(new_n297), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n420), .A2(new_n427), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n551), .A2(new_n552), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT38), .ZN(new_n670));
  INV_X1    g484(.A(new_n646), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n463), .A2(new_n477), .ZN(new_n672));
  AND4_X1   g486(.A1(new_n668), .A2(new_n670), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n661), .A2(new_n667), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G143), .ZN(G45));
  OAI211_X1 g489(.A(new_n617), .B(new_n652), .C1(new_n619), .C2(new_n426), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n650), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n317), .A2(new_n677), .A3(new_n655), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  OR2_X1    g493(.A1(new_n596), .A2(new_n557), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n594), .A2(new_n595), .ZN(new_n681));
  AND4_X1   g495(.A1(new_n597), .A2(new_n681), .A3(new_n557), .A4(new_n188), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n597), .B1(new_n596), .B2(new_n557), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n556), .B(new_n680), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT103), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n599), .A2(new_n686), .A3(new_n556), .A4(new_n680), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n317), .A2(new_n621), .A3(new_n368), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT41), .B(G113), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G15));
  NAND4_X1  g506(.A1(new_n317), .A2(new_n639), .A3(new_n368), .A4(new_n689), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT104), .B(G116), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G18));
  NAND4_X1  g509(.A1(new_n685), .A2(new_n553), .A3(new_n646), .A4(new_n687), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n474), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n317), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n697), .A2(KEYINPUT105), .A3(new_n317), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G119), .ZN(G21));
  NAND3_X1  g517(.A1(new_n668), .A2(new_n669), .A3(new_n672), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n271), .A2(new_n288), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n271), .A2(new_n288), .ZN(new_n707));
  OAI22_X1  g521(.A1(new_n706), .A2(new_n707), .B1(new_n312), .B2(new_n273), .ZN(new_n708));
  NOR2_X1   g522(.A1(G472), .A2(G902), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(G902), .B1(new_n289), .B2(new_n292), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n710), .B1(new_n711), .B2(new_n187), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n367), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n705), .A2(new_n473), .A3(new_n689), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G122), .ZN(G24));
  AND3_X1   g529(.A1(new_n685), .A2(new_n553), .A3(new_n687), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n676), .A2(new_n712), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n716), .A2(new_n717), .A3(KEYINPUT106), .A4(new_n646), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n719));
  AOI22_X1  g533(.A1(new_n622), .A2(G472), .B1(new_n708), .B2(new_n709), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n668), .A2(new_n720), .A3(new_n617), .A4(new_n652), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n719), .B1(new_n721), .B2(new_n696), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT107), .B(G125), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G27));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n726));
  INV_X1    g540(.A(new_n477), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n551), .A2(new_n727), .A3(new_n552), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n600), .B(KEYINPUT108), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n730), .B1(new_n603), .B2(G469), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n555), .B1(new_n599), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n728), .A2(KEYINPUT109), .A3(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n731), .B1(new_n682), .B2(new_n683), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n556), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n551), .A2(new_n727), .A3(new_n552), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n317), .A3(new_n368), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n726), .B1(new_n740), .B2(new_n676), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n316), .A2(new_n297), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n284), .A2(new_n287), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n367), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n676), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n744), .A2(KEYINPUT42), .A3(new_n745), .A4(new_n739), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n741), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G131), .ZN(G33));
  NOR2_X1   g562(.A1(new_n638), .A2(new_n653), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n739), .A2(new_n317), .A3(new_n368), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n604), .B1(new_n752), .B2(new_n557), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n753), .A2(KEYINPUT110), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(KEYINPUT110), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n603), .A2(KEYINPUT45), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(KEYINPUT46), .A3(new_n729), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n599), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT46), .B1(new_n757), .B2(new_n729), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n556), .B(new_n658), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n737), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n619), .A2(new_n426), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n617), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT43), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(KEYINPUT44), .A3(new_n624), .A4(new_n646), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n624), .A3(new_n646), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n769), .A2(new_n771), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT111), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n768), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n228), .ZN(G39));
  NAND3_X1  g590(.A1(new_n745), .A2(new_n367), .A3(new_n728), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n317), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n556), .B1(new_n759), .B2(new_n760), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT47), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(KEYINPUT47), .B(new_n556), .C1(new_n759), .C2(new_n760), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n779), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(new_n327), .ZN(G42));
  AND4_X1   g599(.A1(new_n553), .A2(new_n685), .A3(new_n646), .A4(new_n687), .ZN(new_n786));
  AND4_X1   g600(.A1(KEYINPUT105), .A2(new_n786), .A3(new_n317), .A4(new_n475), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT105), .B1(new_n697), .B2(new_n317), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n693), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n690), .A2(new_n714), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n792));
  INV_X1    g606(.A(new_n462), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n460), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n427), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n792), .B1(new_n795), .B2(new_n619), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n420), .A2(new_n637), .A3(KEYINPUT112), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n610), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n798), .A2(new_n625), .A3(new_n799), .A4(new_n626), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n608), .A2(new_n627), .A3(new_n800), .A4(new_n647), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n801), .B1(new_n741), .B2(new_n746), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n646), .A2(new_n551), .A3(new_n727), .A4(new_n552), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n794), .A2(new_n426), .A3(new_n653), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n636), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n803), .B1(new_n805), .B2(KEYINPUT113), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n636), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n806), .A2(new_n317), .A3(new_n655), .A4(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n712), .A2(new_n671), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n739), .A2(new_n745), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n750), .A2(new_n809), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n750), .A2(new_n809), .A3(new_n811), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT114), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n791), .A2(new_n802), .A3(new_n813), .A4(new_n815), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n736), .A2(new_n646), .A3(new_n653), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n705), .A2(new_n667), .A3(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n723), .A2(new_n656), .A3(new_n678), .A4(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT52), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT53), .B1(new_n816), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n815), .A2(new_n813), .ZN(new_n822));
  INV_X1    g636(.A(new_n790), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n702), .A2(new_n823), .A3(new_n693), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n317), .A2(new_n655), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n827), .A2(new_n654), .B1(new_n718), .B2(new_n722), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(KEYINPUT52), .A3(new_n678), .A4(new_n818), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n819), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n825), .A2(new_n826), .A3(new_n832), .A4(new_n802), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT54), .B1(new_n821), .B2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n825), .A2(new_n832), .A3(new_n802), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT53), .B1(new_n832), .B2(KEYINPUT115), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT54), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n836), .A2(new_n837), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n651), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n766), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n713), .ZN(new_n846));
  OR3_X1    g660(.A1(new_n670), .A2(new_n727), .A3(new_n688), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT50), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n846), .A2(new_n737), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n782), .A2(new_n783), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n599), .A2(new_n680), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n556), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n850), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n688), .A2(new_n737), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n845), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n667), .ZN(new_n858));
  AND4_X1   g672(.A1(new_n368), .A2(new_n858), .A3(new_n465), .A4(new_n855), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n668), .A2(new_n617), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n857), .A2(new_n810), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n849), .A2(new_n854), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT51), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n863), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n859), .A2(new_n668), .A3(new_n617), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n464), .B(KEYINPUT117), .Z(new_n867));
  INV_X1    g681(.A(new_n716), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n866), .B(new_n867), .C1(new_n846), .C2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT118), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  INV_X1    g686(.A(new_n744), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n856), .A2(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n874), .A2(KEYINPUT48), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(KEYINPUT48), .ZN(new_n876));
  NOR4_X1   g690(.A1(new_n871), .A2(new_n872), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n864), .A2(new_n865), .A3(new_n877), .ZN(new_n878));
  OAI22_X1  g692(.A1(new_n843), .A2(new_n878), .B1(G952), .B2(G953), .ZN(new_n879));
  NOR4_X1   g693(.A1(new_n670), .A2(new_n367), .A3(new_n477), .A4(new_n555), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n852), .B(KEYINPUT49), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n881), .A2(new_n764), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n880), .A2(new_n858), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n879), .A2(new_n883), .ZN(G75));
  NOR2_X1   g698(.A1(new_n266), .A2(G952), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n541), .B1(new_n545), .B2(new_n546), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(new_n537), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT55), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n821), .A2(new_n833), .A3(G902), .A4(new_n550), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT56), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n821), .A2(G902), .A3(new_n833), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT119), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n821), .A2(new_n833), .A3(new_n894), .A4(G902), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n893), .A2(new_n550), .A3(new_n895), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n888), .A2(new_n890), .ZN(new_n897));
  AOI211_X1 g711(.A(new_n885), .B(new_n891), .C1(new_n896), .C2(new_n897), .ZN(G51));
  XOR2_X1   g712(.A(new_n729), .B(KEYINPUT57), .Z(new_n899));
  AND3_X1   g713(.A1(new_n821), .A2(KEYINPUT54), .A3(new_n833), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n899), .B1(new_n900), .B2(new_n834), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT120), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n903), .B(new_n899), .C1(new_n900), .C2(new_n834), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n902), .A2(new_n681), .A3(new_n904), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n893), .A2(new_n895), .ZN(new_n906));
  INV_X1    g720(.A(new_n757), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n885), .B1(new_n905), .B2(new_n908), .ZN(G54));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n411), .A2(new_n415), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(KEYINPUT58), .A2(G475), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n906), .A2(new_n910), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n893), .A2(new_n895), .A3(new_n913), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT121), .B1(new_n915), .B2(new_n911), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n885), .B1(new_n915), .B2(new_n911), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n914), .A2(new_n916), .A3(new_n917), .ZN(G60));
  NAND2_X1  g732(.A1(G478), .A2(G902), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT59), .ZN(new_n920));
  OAI221_X1 g734(.A(new_n920), .B1(new_n615), .B2(new_n613), .C1(new_n900), .C2(new_n834), .ZN(new_n921));
  INV_X1    g735(.A(new_n885), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n843), .A2(new_n920), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n613), .A2(new_n615), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(G63));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT60), .Z(new_n928));
  NAND4_X1  g742(.A1(new_n821), .A2(new_n833), .A3(new_n644), .A4(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n922), .ZN(new_n930));
  OAI21_X1  g744(.A(KEYINPUT61), .B1(new_n930), .B2(KEYINPUT122), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n821), .A2(new_n833), .A3(new_n928), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n922), .B(new_n929), .C1(new_n932), .C2(new_n358), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n931), .B(new_n933), .ZN(G66));
  OAI21_X1  g748(.A(G953), .B1(new_n468), .B2(new_n488), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n824), .A2(new_n801), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(G953), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n886), .B1(G898), .B2(new_n266), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G69));
  NAND3_X1  g753(.A1(new_n723), .A2(new_n656), .A3(new_n678), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT124), .Z(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n674), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT62), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n317), .A2(new_n368), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n798), .B1(new_n668), .B2(new_n617), .ZN(new_n946));
  NOR4_X1   g760(.A1(new_n945), .A2(new_n946), .A3(new_n659), .A4(new_n737), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n775), .A2(new_n784), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n944), .A2(new_n266), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n407), .B(KEYINPUT123), .Z(new_n951));
  NOR2_X1   g765(.A1(new_n255), .A2(new_n259), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n951), .B(new_n952), .Z(new_n953));
  NAND3_X1  g767(.A1(new_n949), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n784), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n761), .A2(new_n873), .A3(new_n704), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n955), .A2(new_n957), .A3(new_n750), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n958), .A2(new_n775), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n959), .A2(KEYINPUT125), .A3(new_n747), .A4(new_n941), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n774), .A2(new_n772), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n961), .A2(new_n767), .A3(new_n762), .ZN(new_n962));
  INV_X1    g776(.A(new_n750), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n784), .A2(new_n963), .A3(new_n956), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n962), .A2(new_n941), .A3(new_n964), .A4(new_n747), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT125), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(G953), .B1(new_n960), .B2(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n572), .A2(G900), .A3(G953), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n953), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n954), .B1(new_n968), .B2(new_n970), .ZN(G72));
  NAND2_X1  g785(.A1(new_n300), .A2(new_n270), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n944), .A2(new_n936), .A3(new_n948), .ZN(new_n973));
  NAND2_X1  g787(.A1(G472), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT63), .Z(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT126), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n972), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n260), .A2(new_n264), .A3(new_n301), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n960), .A2(new_n936), .A3(new_n967), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n978), .B1(new_n979), .B2(new_n976), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n840), .A2(new_n841), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n302), .B(KEYINPUT127), .Z(new_n982));
  OAI21_X1  g796(.A(new_n975), .B1(new_n982), .B2(new_n664), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NOR4_X1   g798(.A1(new_n977), .A2(new_n980), .A3(new_n885), .A4(new_n984), .ZN(G57));
endmodule


