//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G120gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G113gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(KEYINPUT69), .B(G113gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(new_n205), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT70), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n211));
  INV_X1    g010(.A(G127gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G134gat), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n212), .A2(G134gat), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n210), .A2(new_n211), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n206), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n205), .A2(G113gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n211), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(KEYINPUT67), .B(G134gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n219), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n213), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT68), .B1(new_n219), .B2(G127gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n218), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n215), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT71), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT25), .ZN(new_n226));
  XOR2_X1   g025(.A(KEYINPUT65), .B(G176gat), .Z(new_n227));
  INV_X1    g026(.A(G169gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(KEYINPUT23), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n230));
  INV_X1    g029(.A(G183gat), .ZN(new_n231));
  INV_X1    g030(.A(G190gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G176gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n228), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n228), .A2(new_n236), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT23), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n229), .A2(new_n235), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n237), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n226), .B1(new_n242), .B2(KEYINPUT23), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n243), .A2(new_n240), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n234), .A2(KEYINPUT66), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n234), .A2(KEYINPUT66), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n233), .A3(new_n246), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n226), .A2(new_n241), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT27), .B(G183gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n232), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT28), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n237), .B1(new_n238), .B2(KEYINPUT26), .ZN(new_n252));
  OR2_X1    g051(.A1(new_n237), .A2(KEYINPUT26), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(new_n231), .B2(new_n232), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n224), .B(new_n225), .C1(new_n248), .C2(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n215), .A2(new_n223), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n248), .A2(new_n256), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT71), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n258), .A2(new_n259), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G227gat), .ZN(new_n263));
  INV_X1    g062(.A(G233gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n265), .B(KEYINPUT64), .Z(new_n266));
  NAND2_X1  g065(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT33), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n204), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(KEYINPUT32), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI221_X1 g070(.A(new_n257), .B1(new_n263), .B2(new_n264), .C1(new_n260), .C2(new_n261), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT34), .ZN(new_n273));
  INV_X1    g072(.A(new_n262), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n266), .A2(KEYINPUT34), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n267), .B(KEYINPUT32), .C1(new_n268), .C2(new_n204), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n271), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n271), .A2(new_n277), .A3(KEYINPUT72), .A4(new_n278), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n271), .A2(new_n278), .ZN(new_n284));
  INV_X1    g083(.A(new_n277), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G204gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G197gat), .ZN(new_n288));
  INV_X1    g087(.A(G197gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G204gat), .ZN(new_n290));
  INV_X1    g089(.A(G211gat), .ZN(new_n291));
  INV_X1    g090(.A(G218gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n288), .B(new_n290), .C1(new_n293), .C2(KEYINPUT22), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT73), .ZN(new_n295));
  XNOR2_X1  g094(.A(G211gat), .B(G218gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G155gat), .B(G162gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G141gat), .B(G148gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT2), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT77), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n299), .B(new_n306), .ZN(new_n307));
  XOR2_X1   g106(.A(KEYINPUT78), .B(KEYINPUT2), .Z(new_n308));
  AOI21_X1  g107(.A(new_n301), .B1(new_n308), .B2(new_n303), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n305), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n310), .A2(KEYINPUT3), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n298), .B1(KEYINPUT29), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n310), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT29), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT3), .B1(new_n297), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n312), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G228gat), .A2(G233gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n317), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT79), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n310), .B(new_n320), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n312), .B(new_n319), .C1(new_n321), .C2(new_n315), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G22gat), .ZN(new_n324));
  INV_X1    g123(.A(G22gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n318), .A2(new_n325), .A3(new_n322), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G78gat), .B(G106gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT31), .B(G50gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT83), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n330), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n327), .B(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n283), .A2(new_n286), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT81), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n215), .A2(new_n223), .A3(new_n313), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n335), .B1(new_n336), .B2(KEYINPUT4), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(KEYINPUT4), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n336), .A2(new_n335), .A3(KEYINPUT4), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G225gat), .A2(G233gat), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n311), .B1(new_n215), .B2(new_n223), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n343), .B1(new_n344), .B2(new_n321), .ZN(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n341), .A2(new_n342), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n336), .B1(new_n258), .B2(new_n321), .ZN(new_n348));
  INV_X1    g147(.A(new_n342), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n346), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(new_n336), .B(KEYINPUT4), .Z(new_n351));
  NAND2_X1  g150(.A1(new_n345), .A2(new_n342), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G1gat), .B(G29gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT0), .ZN(new_n356));
  XNOR2_X1  g155(.A(G57gat), .B(G85gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT6), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n347), .A2(new_n358), .A3(new_n353), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n354), .A2(KEYINPUT6), .A3(new_n359), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AND2_X1   g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  OR3_X1    g166(.A1(new_n259), .A2(KEYINPUT74), .A3(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n259), .A2(new_n367), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n314), .B1(new_n248), .B2(new_n256), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT74), .B1(new_n370), .B2(new_n367), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n368), .B(new_n297), .C1(new_n369), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n367), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(new_n259), .B2(new_n367), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n298), .ZN(new_n375));
  XOR2_X1   g174(.A(G8gat), .B(G36gat), .Z(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT75), .ZN(new_n377));
  XOR2_X1   g176(.A(G64gat), .B(G92gat), .Z(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n372), .A2(new_n375), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT30), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n380), .B1(new_n372), .B2(new_n375), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n381), .A2(KEYINPUT76), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT76), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n372), .A2(new_n375), .A3(new_n387), .A4(new_n380), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n382), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT35), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n365), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n334), .A2(new_n393), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n281), .A2(new_n282), .B1(new_n285), .B2(new_n284), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT82), .ZN(new_n396));
  AOI211_X1 g195(.A(new_n396), .B(new_n390), .C1(new_n364), .C2(new_n363), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT82), .B1(new_n365), .B2(new_n391), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n395), .B(new_n333), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n394), .B1(new_n399), .B2(KEYINPUT35), .ZN(new_n400));
  INV_X1    g199(.A(new_n333), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n401), .B1(new_n397), .B2(new_n398), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT37), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n403), .B1(new_n374), .B2(new_n297), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n368), .B1(new_n369), .B2(new_n371), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n404), .B1(new_n297), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT38), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n372), .A2(new_n375), .A3(new_n403), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .A4(new_n379), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n409), .A2(new_n386), .A3(new_n388), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n379), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n403), .B1(new_n372), .B2(new_n375), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT38), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n363), .A2(new_n410), .A3(new_n364), .A4(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n342), .B1(new_n341), .B2(new_n345), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT39), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT39), .B1(new_n348), .B2(new_n349), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n358), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT40), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  OR2_X1    g220(.A1(new_n415), .A2(new_n419), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT40), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n422), .A2(new_n423), .A3(new_n358), .A4(new_n417), .ZN(new_n424));
  AND2_X1   g223(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n390), .A2(new_n360), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n414), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n333), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n283), .A2(new_n286), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT36), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n395), .A2(KEYINPUT36), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n402), .A2(new_n428), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n400), .A2(new_n433), .ZN(new_n434));
  OR2_X1    g233(.A1(G71gat), .A2(G78gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(G71gat), .A2(G78gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G64gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(G57gat), .ZN(new_n439));
  INV_X1    g238(.A(G57gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(G64gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n437), .B1(KEYINPUT9), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT94), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n435), .A2(new_n444), .A3(new_n436), .ZN(new_n445));
  AND2_X1   g244(.A1(G71gat), .A2(G78gat), .ZN(new_n446));
  NOR2_X1   g245(.A1(G71gat), .A2(G78gat), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT94), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT93), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n438), .B1(new_n451), .B2(G57gat), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n438), .A3(G57gat), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT9), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n453), .A2(new_n454), .B1(new_n455), .B2(new_n436), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n443), .B1(new_n450), .B2(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n457), .A2(KEYINPUT21), .ZN(new_n458));
  NAND2_X1  g257(.A1(G231gat), .A2(G233gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n458), .B(new_n459), .ZN(new_n460));
  XOR2_X1   g259(.A(KEYINPUT95), .B(KEYINPUT19), .Z(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(G127gat), .B(G155gat), .Z(new_n463));
  XNOR2_X1  g262(.A(new_n463), .B(KEYINPUT20), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n462), .B(new_n464), .ZN(new_n465));
  XOR2_X1   g264(.A(G183gat), .B(G211gat), .Z(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(G15gat), .B(G22gat), .ZN(new_n468));
  OR2_X1    g267(.A1(new_n468), .A2(G1gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT89), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT16), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n468), .B1(new_n471), .B2(G1gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(new_n473), .A3(G8gat), .ZN(new_n474));
  INV_X1    g273(.A(G8gat), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n469), .B(new_n472), .C1(KEYINPUT89), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G57gat), .B(G64gat), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n436), .B(new_n435), .C1(new_n478), .C2(new_n455), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n436), .A2(new_n455), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n440), .A2(KEYINPUT93), .A3(G64gat), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n480), .B1(new_n452), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n479), .B1(new_n449), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT96), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n477), .B1(new_n485), .B2(KEYINPUT21), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT97), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n487), .B(KEYINPUT98), .Z(new_n488));
  XNOR2_X1  g287(.A(new_n467), .B(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT88), .ZN(new_n490));
  INV_X1    g289(.A(G43gat), .ZN(new_n491));
  INV_X1    g290(.A(G50gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT85), .ZN(new_n494));
  NAND2_X1  g293(.A1(G43gat), .A2(G50gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT15), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT15), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n493), .A2(new_n494), .A3(new_n498), .A4(new_n495), .ZN(new_n499));
  NAND2_X1  g298(.A1(G29gat), .A2(G36gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT86), .ZN(new_n503));
  NOR4_X1   g302(.A1(new_n503), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n504));
  NOR2_X1   g303(.A1(G29gat), .A2(G36gat), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT14), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT86), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n502), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT87), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g309(.A(KEYINPUT87), .B(new_n502), .C1(new_n504), .C2(new_n507), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n501), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n498), .B1(new_n493), .B2(new_n495), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT84), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n502), .B(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n505), .A2(new_n506), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n514), .B1(new_n518), .B2(new_n500), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n512), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n490), .B1(new_n520), .B2(KEYINPUT17), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT17), .ZN(new_n522));
  OAI211_X1 g321(.A(KEYINPUT88), .B(new_n522), .C1(new_n512), .C2(new_n519), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n521), .A2(new_n523), .B1(KEYINPUT17), .B2(new_n520), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT101), .ZN(new_n525));
  OAI211_X1 g324(.A(G85gat), .B(G92gat), .C1(new_n525), .C2(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g325(.A1(G85gat), .A2(G92gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(KEYINPUT101), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n528), .A2(KEYINPUT101), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT8), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n534), .B1(G99gat), .B2(G106gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT102), .B(G92gat), .ZN(new_n536));
  INV_X1    g335(.A(G85gat), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(G99gat), .A2(G106gat), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT103), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G99gat), .ZN(new_n543));
  INV_X1    g342(.A(G106gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT103), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n545), .A2(new_n546), .A3(new_n539), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n533), .A2(new_n538), .A3(new_n542), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n542), .A2(new_n547), .ZN(new_n549));
  INV_X1    g348(.A(G92gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT102), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT102), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(G92gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n553), .A3(new_n537), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT8), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n531), .B1(new_n526), .B2(new_n529), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n549), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n548), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n524), .A2(KEYINPUT104), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n520), .A2(KEYINPUT17), .ZN(new_n562));
  INV_X1    g361(.A(new_n501), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n517), .A2(new_n503), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n505), .A2(KEYINPUT86), .A3(new_n506), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT87), .B1(new_n566), .B2(new_n502), .ZN(new_n567));
  INV_X1    g366(.A(new_n511), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n563), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n518), .A2(new_n500), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(new_n513), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT88), .B1(new_n572), .B2(new_n522), .ZN(new_n573));
  INV_X1    g372(.A(new_n523), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n562), .B(new_n560), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT104), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT41), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n581), .B1(new_n520), .B2(new_n560), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G190gat), .B(G218gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n585), .B(KEYINPUT105), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n578), .A2(new_n586), .A3(new_n583), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n580), .A2(KEYINPUT41), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT99), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n588), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n586), .B1(new_n578), .B2(new_n583), .ZN(new_n594));
  AOI211_X1 g393(.A(new_n587), .B(new_n582), .C1(new_n561), .C2(new_n577), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n591), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G134gat), .B(G162gat), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT100), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n593), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(new_n593), .B2(new_n596), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G113gat), .B(G141gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT11), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(new_n228), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(new_n289), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT12), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n477), .A2(KEYINPUT90), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT90), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n474), .A2(new_n608), .A3(new_n476), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n562), .B(new_n610), .C1(new_n573), .C2(new_n574), .ZN(new_n611));
  NAND2_X1  g410(.A1(G229gat), .A2(G233gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n572), .A2(new_n477), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT18), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(KEYINPUT91), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n520), .B(new_n477), .ZN(new_n617));
  XOR2_X1   g416(.A(KEYINPUT92), .B(KEYINPUT13), .Z(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(new_n612), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n615), .B1(new_n614), .B2(KEYINPUT91), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n606), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n622), .ZN(new_n624));
  INV_X1    g423(.A(new_n606), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n624), .A2(new_n616), .A3(new_n620), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G120gat), .B(G148gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(G176gat), .B(G204gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT107), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n549), .A2(new_n556), .A3(new_n557), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n533), .A2(new_n538), .B1(new_n542), .B2(new_n547), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n457), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT10), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n548), .A2(new_n483), .A3(new_n558), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT106), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n635), .A2(KEYINPUT106), .A3(new_n636), .A4(new_n637), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n560), .A2(new_n636), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n485), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n632), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n548), .A2(new_n483), .A3(new_n558), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n483), .B1(new_n548), .B2(new_n558), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n648), .A2(new_n631), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n630), .B1(new_n645), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n630), .ZN(new_n651));
  AOI22_X1  g450(.A1(new_n640), .A2(new_n641), .B1(new_n485), .B2(new_n643), .ZN(new_n652));
  INV_X1    g451(.A(new_n631), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n489), .A2(new_n601), .A3(new_n627), .A4(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n434), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n365), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n390), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT16), .B(G8gat), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT42), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(KEYINPUT108), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT108), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n664), .A2(new_n667), .A3(KEYINPUT42), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n669), .B1(new_n662), .B2(G8gat), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n666), .B(new_n668), .C1(new_n664), .C2(new_n670), .ZN(G1325gat));
  INV_X1    g470(.A(new_n658), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n431), .A2(new_n432), .ZN(new_n673));
  OAI21_X1  g472(.A(G15gat), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n429), .A2(G15gat), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n674), .B1(new_n672), .B2(new_n675), .ZN(G1326gat));
  NAND2_X1  g475(.A1(new_n658), .A2(new_n401), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT43), .B(G22gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  INV_X1    g478(.A(new_n601), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(new_n400), .B2(new_n433), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n334), .A2(new_n393), .ZN(new_n684));
  INV_X1    g483(.A(new_n398), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n365), .A2(new_n391), .A3(KEYINPUT82), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n334), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n684), .B1(new_n687), .B2(new_n392), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n402), .A2(new_n428), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n673), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n691), .A2(KEYINPUT44), .A3(new_n680), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n683), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n623), .A2(new_n626), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n489), .A2(new_n694), .A3(new_n655), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(new_n659), .A3(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n693), .A2(KEYINPUT109), .A3(new_n659), .A4(new_n695), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(G29gat), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n681), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n695), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n702), .A2(G29gat), .A3(new_n365), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n703), .A2(KEYINPUT45), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(KEYINPUT45), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n700), .A2(new_n704), .A3(new_n705), .ZN(G1328gat));
  NOR3_X1   g505(.A1(new_n702), .A2(G36gat), .A3(new_n391), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT46), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n390), .A3(new_n695), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G36gat), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(G1329gat));
  INV_X1    g510(.A(new_n673), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n683), .A2(new_n692), .A3(new_n712), .A4(new_n695), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(G43gat), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n701), .A2(new_n491), .A3(new_n395), .A4(new_n695), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT47), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n713), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n713), .A2(new_n719), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n491), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n715), .A2(KEYINPUT47), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n718), .B1(new_n722), .B2(new_n723), .ZN(G1330gat));
  NAND4_X1  g523(.A1(new_n693), .A2(G50gat), .A3(new_n401), .A4(new_n695), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n492), .B1(new_n702), .B2(new_n333), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n725), .A2(KEYINPUT48), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT48), .B1(new_n725), .B2(new_n726), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(G1331gat));
  NAND3_X1  g528(.A1(new_n489), .A2(new_n601), .A3(new_n694), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n656), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n691), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(new_n365), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(new_n440), .ZN(G1332gat));
  AOI211_X1 g533(.A(new_n391), .B(new_n732), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n735));
  NOR2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1333gat));
  INV_X1    g536(.A(new_n732), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n738), .A2(G71gat), .A3(new_n712), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n732), .A2(new_n429), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(G71gat), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g541(.A1(new_n738), .A2(new_n401), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g543(.A1(new_n489), .A2(new_n627), .A3(new_n656), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n693), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(G85gat), .B1(new_n746), .B2(new_n365), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n489), .A2(new_n627), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n701), .A2(KEYINPUT111), .A3(KEYINPUT51), .A4(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n691), .A2(KEYINPUT51), .A3(new_n680), .A4(new_n748), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n680), .B(new_n748), .C1(new_n400), .C2(new_n433), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n749), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n756), .A2(new_n537), .A3(new_n659), .A4(new_n655), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n747), .A2(new_n757), .ZN(G1336gat));
  NOR3_X1   g557(.A1(new_n391), .A2(G92gat), .A3(new_n656), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n683), .A2(new_n692), .A3(new_n390), .A4(new_n745), .ZN(new_n761));
  INV_X1    g560(.A(new_n536), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XOR2_X1   g562(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n755), .A2(new_n750), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n761), .A2(new_n762), .B1(new_n767), .B2(new_n759), .ZN(new_n768));
  OAI22_X1  g567(.A1(new_n760), .A2(new_n765), .B1(new_n766), .B2(new_n768), .ZN(G1337gat));
  OAI21_X1  g568(.A(G99gat), .B1(new_n746), .B2(new_n673), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n756), .A2(new_n543), .A3(new_n395), .A4(new_n655), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(G1338gat));
  NAND3_X1  g571(.A1(new_n401), .A2(new_n544), .A3(new_n655), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n773), .B(KEYINPUT113), .Z(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n756), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n683), .A2(new_n692), .A3(new_n401), .A4(new_n745), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT53), .B1(new_n777), .B2(G106gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n777), .A2(G106gat), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n767), .B2(new_n775), .ZN(new_n782));
  AOI211_X1 g581(.A(KEYINPUT114), .B(new_n774), .C1(new_n755), .C2(new_n750), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n779), .B1(new_n784), .B2(new_n785), .ZN(G1339gat));
  NOR2_X1   g585(.A1(new_n694), .A2(new_n207), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n730), .A2(new_n655), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n630), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n645), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT106), .B1(new_n648), .B2(new_n636), .ZN(new_n793));
  INV_X1    g592(.A(new_n641), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n644), .B(new_n632), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n795), .B(KEYINPUT54), .C1(new_n653), .C2(new_n652), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n792), .A2(new_n796), .A3(KEYINPUT55), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n654), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n797), .A2(KEYINPUT115), .A3(new_n654), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n792), .A2(new_n796), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n800), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n605), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n612), .B1(new_n611), .B2(new_n613), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n617), .A2(new_n619), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n626), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n806), .B(new_n811), .C1(new_n599), .C2(new_n600), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n626), .A2(new_n655), .A3(new_n810), .ZN(new_n813));
  OAI211_X1 g612(.A(KEYINPUT116), .B(new_n813), .C1(new_n805), .C2(new_n694), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n601), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n627), .A2(new_n801), .A3(new_n800), .A4(new_n804), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT116), .B1(new_n816), .B2(new_n813), .ZN(new_n817));
  OAI211_X1 g616(.A(KEYINPUT117), .B(new_n812), .C1(new_n815), .C2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n489), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n813), .B1(new_n805), .B2(new_n694), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(new_n601), .A3(new_n814), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT117), .B1(new_n824), .B2(new_n812), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n789), .B1(new_n820), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n659), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n334), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n828), .A2(KEYINPUT118), .A3(new_n391), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT118), .B1(new_n828), .B2(new_n391), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n787), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n828), .A2(new_n391), .ZN(new_n832));
  OAI21_X1  g631(.A(G113gat), .B1(new_n832), .B2(new_n694), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(G1340gat));
  OAI211_X1 g633(.A(new_n205), .B(new_n655), .C1(new_n829), .C2(new_n830), .ZN(new_n835));
  OAI21_X1  g634(.A(G120gat), .B1(new_n832), .B2(new_n656), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(G1341gat));
  NOR2_X1   g636(.A1(new_n832), .A2(new_n819), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(new_n212), .ZN(G1342gat));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840));
  INV_X1    g639(.A(new_n334), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n601), .A2(new_n390), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n826), .A2(new_n659), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n845), .A3(new_n219), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n843), .A2(G134gat), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n845), .B1(new_n844), .B2(new_n219), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n840), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n849), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n851), .A2(new_n846), .A3(KEYINPUT119), .A4(new_n847), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(G1343gat));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n826), .A2(new_n854), .A3(new_n401), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n673), .A2(new_n659), .A3(new_n391), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n804), .A2(new_n654), .A3(new_n797), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n858), .B1(new_n623), .B2(new_n626), .ZN(new_n859));
  INV_X1    g658(.A(new_n813), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI211_X1 g660(.A(KEYINPUT120), .B(new_n813), .C1(new_n694), .C2(new_n858), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n862), .A3(new_n601), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n489), .B1(new_n863), .B2(new_n812), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n401), .B1(new_n864), .B2(new_n788), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n856), .B1(new_n865), .B2(KEYINPUT57), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n855), .A2(new_n627), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n395), .A2(KEYINPUT36), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n283), .A2(KEYINPUT36), .A3(new_n286), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n401), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n673), .A2(KEYINPUT121), .A3(new_n401), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n826), .A2(new_n659), .A3(new_n391), .A4(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n694), .A2(G141gat), .ZN(new_n877));
  AOI22_X1  g676(.A1(new_n867), .A2(G141gat), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n879), .B1(new_n867), .B2(G141gat), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n878), .A2(new_n880), .A3(KEYINPUT58), .ZN(new_n881));
  INV_X1    g680(.A(new_n877), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n875), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884));
  AOI221_X4 g683(.A(new_n883), .B1(new_n879), .B2(new_n884), .C1(G141gat), .C2(new_n867), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n881), .A2(new_n885), .ZN(G1344gat));
  INV_X1    g685(.A(G148gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n876), .A2(new_n887), .A3(new_n655), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n865), .A2(KEYINPUT57), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n826), .A2(new_n401), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(KEYINPUT57), .ZN(new_n892));
  INV_X1    g691(.A(new_n856), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n655), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n889), .B1(new_n894), .B2(G148gat), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n855), .A2(new_n866), .ZN(new_n896));
  AOI211_X1 g695(.A(KEYINPUT59), .B(new_n887), .C1(new_n896), .C2(new_n655), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n888), .B1(new_n895), .B2(new_n897), .ZN(G1345gat));
  INV_X1    g697(.A(G155gat), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n876), .A2(new_n899), .A3(new_n489), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n896), .A2(new_n489), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(new_n899), .ZN(G1346gat));
  NAND2_X1  g701(.A1(new_n896), .A2(new_n680), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(G162gat), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n601), .A2(G162gat), .A3(new_n390), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n826), .A2(new_n659), .A3(new_n874), .A4(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1347gat));
  NOR2_X1   g706(.A1(new_n659), .A2(new_n391), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n826), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n841), .ZN(new_n910));
  OR4_X1    g709(.A1(KEYINPUT123), .A2(new_n910), .A3(G169gat), .A4(new_n694), .ZN(new_n911));
  INV_X1    g710(.A(new_n910), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n627), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT123), .B1(new_n913), .B2(G169gat), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n913), .A2(G169gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n911), .B1(new_n914), .B2(new_n915), .ZN(G1348gat));
  NAND3_X1  g715(.A1(new_n909), .A2(new_n841), .A3(new_n655), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n917), .A2(new_n918), .A3(new_n236), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n917), .B2(new_n236), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n917), .A2(new_n227), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(G1349gat));
  AOI21_X1  g721(.A(new_n231), .B1(new_n912), .B2(new_n489), .ZN(new_n923));
  INV_X1    g722(.A(new_n249), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n910), .A2(new_n924), .A3(new_n819), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT60), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n912), .A2(new_n249), .A3(new_n489), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT60), .ZN(new_n928));
  OAI21_X1  g727(.A(G183gat), .B1(new_n910), .B2(new_n819), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n926), .A2(new_n930), .ZN(G1350gat));
  NAND3_X1  g730(.A1(new_n909), .A2(new_n841), .A3(new_n680), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n932), .A2(new_n933), .A3(G190gat), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n932), .B2(G190gat), .ZN(new_n935));
  OAI22_X1  g734(.A1(new_n934), .A2(new_n935), .B1(G190gat), .B2(new_n932), .ZN(G1351gat));
  INV_X1    g735(.A(new_n870), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n909), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g737(.A(KEYINPUT125), .B(G197gat), .Z(new_n939));
  OR3_X1    g738(.A1(new_n938), .A2(new_n694), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n673), .A2(new_n908), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n892), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT126), .B1(new_n943), .B2(new_n627), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n892), .A2(KEYINPUT126), .A3(new_n627), .A4(new_n942), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n939), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n940), .B1(new_n944), .B2(new_n946), .ZN(G1352gat));
  NAND3_X1  g746(.A1(new_n892), .A2(new_n655), .A3(new_n942), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G204gat), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n909), .A2(new_n287), .A3(new_n655), .A4(new_n937), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n950), .A2(KEYINPUT62), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(KEYINPUT62), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n952), .A2(KEYINPUT127), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n954), .B1(new_n950), .B2(KEYINPUT62), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n949), .B(new_n951), .C1(new_n953), .C2(new_n955), .ZN(G1353gat));
  INV_X1    g755(.A(new_n938), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n957), .A2(new_n291), .A3(new_n489), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n892), .A2(new_n489), .A3(new_n942), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n959), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT63), .B1(new_n959), .B2(G211gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(G1354gat));
  NAND3_X1  g762(.A1(new_n957), .A2(new_n292), .A3(new_n680), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n943), .A2(new_n680), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(new_n292), .ZN(G1355gat));
endmodule


