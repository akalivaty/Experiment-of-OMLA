//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1176, new_n1177,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT65), .Z(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(new_n202), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G50), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT0), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT66), .B(G77), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  AND2_X1   g0021(.A1(new_n221), .A2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G58), .A2(G232), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n216), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n215), .B(new_n219), .C1(new_n228), .C2(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n235), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(new_n243), .B(KEYINPUT68), .Z(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n212), .B1(new_n216), .B2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n204), .A2(G20), .ZN(new_n252));
  INV_X1    g0052(.A(G58), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT8), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT8), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G58), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n249), .A2(G20), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n257), .A2(new_n258), .B1(G150), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n251), .B1(new_n252), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT72), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n262), .A2(KEYINPUT72), .A3(G13), .A4(G20), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G50), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n250), .B1(new_n265), .B2(new_n266), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n269), .B1(new_n262), .B2(G20), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n268), .A2(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n261), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT69), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT69), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G45), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT70), .ZN(new_n281));
  AND3_X1   g0081(.A1(new_n280), .A2(new_n281), .A3(new_n262), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n281), .B1(new_n280), .B2(new_n262), .ZN(new_n283));
  AND2_X1   g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  OAI21_X1  g0084(.A(KEYINPUT71), .B1(new_n284), .B2(new_n212), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT71), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n286), .A2(new_n287), .A3(G1), .A4(G13), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n285), .A2(G274), .A3(new_n288), .ZN(new_n289));
  NOR3_X1   g0089(.A1(new_n282), .A2(new_n283), .A3(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n291));
  AND3_X1   g0091(.A1(new_n285), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n290), .B1(G226), .B2(new_n292), .ZN(new_n293));
  AND2_X1   g0093(.A1(KEYINPUT3), .A2(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(KEYINPUT3), .A2(G33), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G1698), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G223), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT3), .B(G33), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n299), .B1(new_n220), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n296), .A2(G1698), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(G222), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n284), .A2(new_n212), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n293), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n274), .A2(KEYINPUT9), .B1(G200), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  OAI221_X1 g0108(.A(new_n307), .B1(KEYINPUT9), .B2(new_n274), .C1(new_n308), .C2(new_n306), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT10), .ZN(new_n310));
  INV_X1    g0110(.A(new_n257), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n262), .A2(G20), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n257), .A2(new_n312), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n268), .A2(new_n311), .B1(new_n270), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT7), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n300), .B2(G20), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n296), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT76), .ZN(new_n318));
  NOR4_X1   g0118(.A1(new_n294), .A2(new_n295), .A3(new_n315), .A4(G20), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT76), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n318), .A2(G68), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G68), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n253), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(G20), .B1(new_n324), .B2(new_n202), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n259), .A2(G159), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT16), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT7), .B1(new_n296), .B2(new_n213), .ZN(new_n330));
  OAI21_X1  g0130(.A(G68), .B1(new_n330), .B2(new_n319), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(KEYINPUT16), .A3(new_n328), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n250), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n314), .B1(new_n329), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G200), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n285), .A2(G232), .A3(new_n288), .A4(new_n291), .ZN(new_n336));
  NOR2_X1   g0136(.A1(G223), .A2(G1698), .ZN(new_n337));
  INV_X1    g0137(.A(G226), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(G1698), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(new_n300), .B1(G33), .B2(G87), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n336), .B1(new_n340), .B2(new_n305), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n335), .B1(new_n290), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n338), .A2(G1698), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(G223), .B2(G1698), .ZN(new_n344));
  INV_X1    g0144(.A(G87), .ZN(new_n345));
  OAI22_X1  g0145(.A1(new_n344), .A2(new_n296), .B1(new_n249), .B2(new_n345), .ZN(new_n346));
  AOI22_X1  g0146(.A1(G232), .A2(new_n292), .B1(new_n346), .B2(new_n304), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n280), .A2(new_n262), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT70), .ZN(new_n349));
  AND3_X1   g0149(.A1(new_n285), .A2(G274), .A3(new_n288), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n280), .A2(new_n281), .A3(new_n262), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n347), .A2(new_n352), .A3(new_n308), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n342), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(KEYINPUT77), .A2(KEYINPUT17), .ZN(new_n355));
  NAND2_X1  g0155(.A1(KEYINPUT77), .A2(KEYINPUT17), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n334), .A2(new_n354), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n329), .A2(new_n333), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n342), .A2(new_n353), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n359), .A2(new_n314), .A3(new_n360), .A4(new_n356), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(G169), .B1(new_n290), .B2(new_n341), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n347), .A2(new_n352), .A3(G179), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n334), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT18), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT18), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n334), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n362), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G169), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n274), .B1(new_n372), .B2(new_n306), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(G179), .B2(new_n306), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n298), .A2(G238), .B1(G107), .B2(new_n296), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n300), .A2(new_n297), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n232), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n304), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n292), .A2(G244), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n352), .A3(new_n379), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n380), .A2(G179), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n257), .A2(new_n259), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n213), .A2(G33), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT15), .B(G87), .ZN(new_n384));
  OAI221_X1 g0184(.A(new_n382), .B1(new_n213), .B2(new_n220), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n385), .A2(new_n250), .B1(new_n220), .B2(new_n268), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n270), .A2(G77), .A3(new_n312), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT73), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT73), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n386), .A2(new_n390), .A3(new_n387), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n380), .A2(new_n372), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n381), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n380), .A2(G200), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n378), .A2(new_n379), .A3(G190), .A4(new_n352), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n395), .A2(new_n391), .A3(new_n389), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  XOR2_X1   g0198(.A(new_n398), .B(KEYINPUT74), .Z(new_n399));
  NAND4_X1  g0199(.A1(new_n310), .A2(new_n371), .A3(new_n374), .A4(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n268), .A2(new_n323), .ZN(new_n401));
  XNOR2_X1  g0201(.A(new_n401), .B(KEYINPUT12), .ZN(new_n402));
  INV_X1    g0202(.A(new_n259), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(new_n269), .ZN(new_n404));
  INV_X1    g0204(.A(G77), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n383), .A2(new_n405), .B1(new_n213), .B2(G68), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n250), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT11), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n270), .A2(G68), .A3(new_n312), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n402), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n285), .A2(G238), .A3(new_n288), .A4(new_n291), .ZN(new_n411));
  NOR2_X1   g0211(.A1(G226), .A2(G1698), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n232), .B2(G1698), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n300), .B1(G33), .B2(G97), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n411), .B1(new_n414), .B2(new_n305), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT13), .B1(new_n290), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G97), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n232), .A2(G1698), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(G226), .B2(G1698), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n417), .B1(new_n419), .B2(new_n296), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n292), .A2(G238), .B1(new_n420), .B2(new_n304), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT13), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n352), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT75), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n416), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n421), .A2(new_n352), .A3(KEYINPUT75), .A4(new_n422), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(G169), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT14), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n425), .A2(KEYINPUT14), .A3(G169), .A4(new_n426), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n416), .A2(G179), .A3(new_n423), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n410), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n425), .A2(G200), .A3(new_n426), .ZN(new_n434));
  INV_X1    g0234(.A(new_n410), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n416), .A2(G190), .A3(new_n423), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n400), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(G257), .B(new_n297), .C1(new_n294), .C2(new_n295), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT80), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n440), .B(new_n441), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n298), .A2(G264), .B1(G303), .B2(new_n296), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n305), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT5), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n262), .B(G45), .C1(new_n445), .C2(G41), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n276), .A2(new_n278), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n446), .B1(new_n447), .B2(new_n445), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n350), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(G270), .ZN(new_n450));
  AOI21_X1  g0250(.A(KEYINPUT5), .B1(new_n276), .B2(new_n278), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n285), .B(new_n288), .C1(new_n451), .C2(new_n446), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n449), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n444), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(new_n372), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT81), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G283), .ZN(new_n457));
  INV_X1    g0257(.A(G97), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n457), .B(new_n213), .C1(G33), .C2(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n459), .B(new_n250), .C1(new_n213), .C2(G116), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n460), .B(KEYINPUT20), .ZN(new_n461));
  INV_X1    g0261(.A(G116), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n268), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n262), .A2(G33), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n270), .A2(G116), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n456), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT20), .ZN(new_n468));
  XNOR2_X1  g0268(.A(new_n460), .B(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n469), .A2(KEYINPUT81), .A3(new_n465), .A4(new_n463), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT21), .B1(new_n455), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT82), .ZN(new_n473));
  OAI211_X1 g0273(.A(KEYINPUT21), .B(G169), .C1(new_n444), .C2(new_n453), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n442), .A2(new_n443), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n304), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n285), .A2(new_n288), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n448), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(G270), .B1(new_n350), .B2(new_n448), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n476), .A2(G179), .A3(new_n479), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n471), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n473), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n474), .A2(new_n480), .B1(new_n467), .B2(new_n470), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT82), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n472), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n454), .A2(G190), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n482), .B(new_n487), .C1(new_n335), .C2(new_n454), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n318), .A2(G107), .A3(new_n321), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n259), .A2(G77), .ZN(new_n492));
  XNOR2_X1  g0292(.A(new_n492), .B(KEYINPUT78), .ZN(new_n493));
  INV_X1    g0293(.A(G107), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(KEYINPUT6), .A3(G97), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n458), .A2(new_n494), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(new_n206), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n495), .B1(new_n497), .B2(KEYINPUT6), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n493), .B1(G20), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n251), .B1(new_n491), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n270), .A2(G97), .A3(new_n464), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n501), .B1(G97), .B2(new_n267), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n300), .A2(G250), .A3(G1698), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n300), .A2(G244), .A3(new_n297), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT4), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n457), .B(new_n504), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT4), .B1(new_n302), .B2(G244), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n304), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n478), .A2(G257), .B1(new_n350), .B2(new_n448), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G200), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n503), .B(new_n512), .C1(new_n308), .C2(new_n511), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n372), .ZN(new_n514));
  INV_X1    g0314(.A(G179), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n509), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n514), .B(new_n516), .C1(new_n500), .C2(new_n502), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT23), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n213), .B2(G107), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n494), .A2(KEYINPUT23), .A3(G20), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n520), .A2(new_n521), .B1(new_n258), .B2(G116), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT22), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n296), .A2(G20), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(G87), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n300), .A2(new_n213), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n526), .A2(KEYINPUT22), .A3(new_n345), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n522), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT24), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n251), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(KEYINPUT24), .B(new_n522), .C1(new_n525), .C2(new_n527), .ZN(new_n531));
  OR3_X1    g0331(.A1(new_n267), .A2(KEYINPUT25), .A3(G107), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n270), .A2(G107), .A3(new_n464), .ZN(new_n533));
  OAI21_X1  g0333(.A(KEYINPUT25), .B1(new_n267), .B2(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT83), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT83), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n532), .A2(new_n533), .A3(new_n534), .A4(new_n537), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n530), .A2(new_n531), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n300), .A2(G257), .A3(G1698), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G294), .ZN(new_n541));
  INV_X1    g0341(.A(G250), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n540), .B(new_n541), .C1(new_n376), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n304), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n478), .A2(G264), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(new_n545), .A3(new_n449), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n335), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n544), .A2(new_n545), .A3(new_n308), .A4(new_n449), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(KEYINPUT84), .A3(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT84), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n546), .A2(new_n550), .A3(new_n335), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n539), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n518), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n546), .A2(new_n372), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(G179), .B2(new_n546), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n539), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n300), .A2(G238), .A3(new_n297), .ZN(new_n557));
  OAI211_X1 g0357(.A(G244), .B(G1698), .C1(new_n294), .C2(new_n295), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G33), .A2(G116), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n304), .ZN(new_n561));
  OR3_X1    g0361(.A1(new_n279), .A2(G1), .A3(G274), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n542), .B1(new_n279), .B2(G1), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n285), .A2(new_n562), .A3(new_n288), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G200), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT19), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n213), .B1(new_n417), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(G87), .B2(new_n207), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n567), .B1(new_n383), .B2(new_n458), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n569), .B(new_n570), .C1(new_n526), .C2(new_n323), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n571), .A2(new_n250), .B1(new_n268), .B2(new_n384), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n561), .A2(G190), .A3(new_n564), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n270), .A2(G87), .A3(new_n464), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n566), .A2(new_n572), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  XOR2_X1   g0375(.A(new_n384), .B(KEYINPUT79), .Z(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(new_n270), .A3(new_n464), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(G179), .B2(new_n565), .ZN(new_n579));
  INV_X1    g0379(.A(new_n565), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n580), .A2(G169), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n575), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n553), .A2(new_n556), .A3(new_n582), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n439), .A2(new_n490), .A3(new_n583), .ZN(G372));
  INV_X1    g0384(.A(KEYINPUT86), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n564), .A2(new_n585), .ZN(new_n586));
  OR2_X1    g0386(.A1(new_n564), .A2(new_n585), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT85), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n560), .A2(new_n588), .A3(new_n304), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n588), .B1(new_n560), .B2(new_n304), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n586), .B(new_n587), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n372), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n580), .A2(new_n515), .B1(new_n572), .B2(new_n577), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n591), .A2(G200), .B1(G190), .B2(new_n580), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n572), .A2(new_n574), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT87), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT87), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n572), .A2(new_n598), .A3(new_n574), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n595), .A2(new_n600), .B1(new_n592), .B2(new_n593), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n601), .A2(new_n552), .A3(new_n517), .A4(new_n513), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n556), .A2(new_n472), .A3(new_n484), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n594), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n514), .A2(new_n516), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n605), .A2(new_n503), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT26), .B1(new_n601), .B2(new_n606), .ZN(new_n607));
  XOR2_X1   g0407(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n608));
  NOR3_X1   g0408(.A1(new_n582), .A2(new_n517), .A3(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  OR2_X1    g0410(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n439), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n437), .A2(new_n381), .A3(new_n392), .A4(new_n393), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n362), .B1(new_n433), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n310), .B1(new_n370), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n374), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n612), .A2(new_n617), .ZN(G369));
  NAND3_X1  g0418(.A1(new_n262), .A2(new_n213), .A3(G13), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n619), .A2(KEYINPUT27), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n620), .B(KEYINPUT89), .ZN(new_n621));
  INV_X1    g0421(.A(G213), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n619), .B2(KEYINPUT27), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(G343), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n482), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n472), .B2(new_n484), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n489), .B2(new_n627), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(G330), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n556), .A2(new_n626), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n539), .A2(new_n626), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n632), .A2(new_n552), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n631), .B1(new_n633), .B2(new_n556), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n634), .ZN(new_n636));
  INV_X1    g0436(.A(new_n626), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n486), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n631), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n635), .A2(new_n640), .ZN(G399));
  INV_X1    g0441(.A(new_n217), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(new_n447), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(G1), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n210), .B2(new_n644), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n647), .B(KEYINPUT28), .ZN(new_n648));
  INV_X1    g0448(.A(new_n556), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n602), .B1(new_n486), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n595), .A2(new_n600), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n606), .A2(new_n651), .A3(KEYINPUT26), .A4(new_n594), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n608), .B1(new_n582), .B2(new_n517), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n594), .ZN(new_n655));
  OAI211_X1 g0455(.A(KEYINPUT29), .B(new_n626), .C1(new_n650), .C2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(KEYINPUT93), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT93), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n611), .A2(new_n626), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT29), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n657), .B1(new_n661), .B2(new_n656), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT92), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT90), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n480), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n476), .A2(KEYINPUT90), .A3(G179), .A4(new_n479), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n544), .A2(new_n545), .A3(new_n561), .A4(new_n564), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n511), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT30), .ZN(new_n670));
  INV_X1    g0470(.A(new_n511), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n546), .A2(new_n515), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n671), .A2(new_n672), .A3(new_n454), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n669), .A2(new_n670), .B1(new_n673), .B2(new_n591), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n665), .A2(KEYINPUT30), .A3(new_n666), .A4(new_n668), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n675), .A2(KEYINPUT91), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(KEYINPUT91), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n678), .A2(KEYINPUT31), .A3(new_n637), .ZN(new_n679));
  AOI21_X1  g0479(.A(KEYINPUT31), .B1(new_n678), .B2(new_n637), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n663), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n678), .A2(new_n637), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT31), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n678), .A2(KEYINPUT31), .A3(new_n637), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(KEYINPUT92), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n490), .A2(new_n583), .A3(new_n626), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n681), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G330), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n662), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n648), .B1(new_n691), .B2(G1), .ZN(G364));
  AND2_X1   g0492(.A1(new_n213), .A2(G13), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n262), .B1(new_n693), .B2(G45), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OR3_X1    g0495(.A1(new_n695), .A2(new_n643), .A3(KEYINPUT94), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT94), .B1(new_n695), .B2(new_n643), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n699), .B1(new_n629), .B2(G330), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(G330), .B2(new_n629), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n642), .A2(new_n300), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n279), .B2(new_n211), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n247), .B2(new_n279), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n642), .A2(new_n296), .ZN(new_n706));
  AOI22_X1  g0506(.A1(new_n706), .A2(G355), .B1(new_n462), .B2(new_n642), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n705), .A2(KEYINPUT95), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(G13), .A2(G33), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G20), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n212), .B1(G20), .B2(new_n372), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT95), .B1(new_n705), .B2(new_n707), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n699), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n213), .A2(new_n515), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(new_n308), .A3(new_n335), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n300), .B1(new_n718), .B2(new_n220), .ZN(new_n719));
  NOR4_X1   g0519(.A1(new_n213), .A2(new_n335), .A3(G179), .A4(G190), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n494), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n717), .A2(G190), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n335), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n722), .B1(G50), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n723), .A2(G200), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR4_X1   g0527(.A1(new_n213), .A2(new_n308), .A3(new_n335), .A4(G179), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI221_X1 g0529(.A(new_n725), .B1(new_n253), .B2(new_n727), .C1(new_n345), .C2(new_n729), .ZN(new_n730));
  NOR4_X1   g0530(.A1(new_n213), .A2(new_n515), .A3(new_n335), .A4(G190), .ZN(new_n731));
  AOI211_X1 g0531(.A(new_n719), .B(new_n730), .C1(G68), .C2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G179), .A2(G200), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT96), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n734), .A2(new_n213), .A3(G190), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G159), .ZN(new_n737));
  OR3_X1    g0537(.A1(new_n736), .A2(KEYINPUT32), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(G20), .B1(new_n734), .B2(new_n308), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G97), .ZN(new_n740));
  OAI21_X1  g0540(.A(KEYINPUT32), .B1(new_n736), .B2(new_n737), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n732), .A2(new_n738), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n739), .ZN(new_n743));
  INV_X1    g0543(.A(G294), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G322), .ZN(new_n746));
  INV_X1    g0546(.A(new_n724), .ZN(new_n747));
  INV_X1    g0547(.A(G326), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n746), .A2(new_n727), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G303), .ZN(new_n750));
  INV_X1    g0550(.A(G283), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n729), .A2(new_n750), .B1(new_n721), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(KEYINPUT33), .B(G317), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n731), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n718), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n300), .B(new_n755), .C1(G311), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n735), .A2(G329), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n753), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n742), .B1(new_n745), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n716), .B1(new_n760), .B2(new_n712), .ZN(new_n761));
  INV_X1    g0561(.A(new_n711), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n761), .B1(new_n629), .B2(new_n762), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n701), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(G396));
  NOR2_X1   g0565(.A1(new_n394), .A2(new_n637), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n392), .A2(new_n637), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT100), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n392), .A2(KEYINPUT100), .A3(new_n637), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n769), .A2(new_n397), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n766), .B1(new_n771), .B2(new_n394), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n659), .B(new_n772), .Z(new_n773));
  AOI21_X1  g0573(.A(new_n699), .B1(new_n773), .B2(new_n689), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(new_n689), .B2(new_n773), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n712), .A2(new_n709), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n698), .B1(new_n405), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n712), .ZN(new_n778));
  INV_X1    g0578(.A(new_n731), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n296), .B1(new_n462), .B2(new_n718), .C1(new_n779), .C2(new_n751), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(G311), .B2(new_n735), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n726), .A2(G294), .B1(G87), .B2(new_n720), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n724), .A2(G303), .B1(G107), .B2(new_n728), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n781), .A2(new_n740), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT97), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n296), .B1(new_n735), .B2(G132), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT99), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n721), .A2(new_n323), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(G50), .B2(new_n728), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n787), .B(new_n789), .C1(new_n253), .C2(new_n743), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n756), .A2(G159), .B1(new_n731), .B2(G150), .ZN(new_n791));
  INV_X1    g0591(.A(G143), .ZN(new_n792));
  INV_X1    g0592(.A(G137), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n791), .B1(new_n727), .B2(new_n792), .C1(new_n793), .C2(new_n747), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT98), .Z(new_n795));
  AOI21_X1  g0595(.A(new_n790), .B1(KEYINPUT34), .B2(new_n795), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n795), .A2(KEYINPUT34), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n785), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n777), .B1(new_n778), .B2(new_n798), .C1(new_n772), .C2(new_n710), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n775), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(G384));
  NOR2_X1   g0601(.A1(new_n693), .A2(new_n262), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT38), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT37), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n316), .A2(new_n317), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n327), .B1(new_n805), .B2(G68), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(KEYINPUT16), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n314), .B1(new_n807), .B2(new_n333), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n365), .B2(new_n625), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n360), .B(new_n314), .C1(new_n329), .C2(new_n333), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n804), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n366), .A2(new_n810), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT104), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n334), .A2(new_n625), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n812), .A2(new_n813), .A3(new_n804), .A4(new_n814), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n366), .A2(new_n814), .A3(new_n810), .A4(new_n804), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(KEYINPUT104), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n811), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n808), .A2(new_n625), .ZN(new_n819));
  INV_X1    g0619(.A(new_n370), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n358), .A2(new_n361), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n803), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n811), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n816), .A2(KEYINPUT104), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n816), .A2(KEYINPUT104), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n625), .B(new_n808), .C1(new_n362), .C2(new_n370), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n827), .A2(KEYINPUT38), .A3(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT105), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n823), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  OAI211_X1 g0631(.A(KEYINPUT105), .B(new_n803), .C1(new_n818), .C2(new_n822), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT39), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT107), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n370), .B1(new_n362), .B2(KEYINPUT106), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT106), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n821), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n814), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n804), .B1(new_n812), .B2(new_n814), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(new_n815), .B2(new_n817), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n803), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(KEYINPUT39), .B1(new_n842), .B2(new_n829), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n834), .A2(new_n835), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n433), .A2(new_n637), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT39), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n831), .B2(new_n832), .ZN(new_n848));
  OAI21_X1  g0648(.A(KEYINPUT107), .B1(new_n848), .B2(new_n843), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n845), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n833), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n432), .B1(new_n429), .B2(new_n430), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n437), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n853), .A2(new_n410), .A3(new_n637), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n410), .A2(new_n637), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT102), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n433), .A2(KEYINPUT103), .A3(new_n437), .A4(new_n856), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n856), .B(new_n437), .C1(new_n852), .C2(new_n435), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT103), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n772), .B(new_n626), .C1(new_n604), .C2(new_n610), .ZN(new_n862));
  INV_X1    g0662(.A(new_n766), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n854), .A2(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n851), .A2(new_n864), .B1(new_n370), .B2(new_n624), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n850), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n439), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n867), .A2(new_n662), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n868), .A2(new_n616), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n866), .B(new_n869), .Z(new_n870));
  INV_X1    g0670(.A(G330), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT40), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n861), .A2(new_n854), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n687), .A2(new_n684), .A3(new_n685), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n873), .A2(new_n874), .A3(new_n772), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n872), .B1(new_n875), .B2(new_n833), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n872), .B1(new_n842), .B2(new_n829), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n877), .A2(new_n772), .A3(new_n873), .A4(new_n874), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n439), .A2(new_n874), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n871), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n881), .B2(new_n880), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n802), .B1(new_n870), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n870), .B2(new_n883), .ZN(new_n885));
  OR2_X1    g0685(.A1(new_n498), .A2(KEYINPUT35), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n498), .A2(KEYINPUT35), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n886), .A2(G116), .A3(new_n214), .A4(new_n887), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n888), .B(KEYINPUT36), .Z(new_n889));
  NOR3_X1   g0689(.A1(new_n210), .A2(new_n220), .A3(new_n324), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n890), .A2(KEYINPUT101), .B1(G68), .B2(new_n201), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(KEYINPUT101), .B2(new_n890), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n262), .A2(G13), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n885), .A2(new_n894), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n895), .B(KEYINPUT108), .Z(G367));
  OAI21_X1  g0696(.A(new_n518), .B1(new_n503), .B2(new_n626), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n606), .A2(new_n637), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n640), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT45), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT44), .B1(new_n640), .B2(new_n900), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n640), .A2(KEYINPUT44), .A3(new_n900), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(new_n635), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n634), .B(new_n638), .Z(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(new_n630), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n691), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n643), .B(KEYINPUT41), .Z(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n695), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n636), .A2(new_n638), .A3(new_n899), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n916), .A2(KEYINPUT42), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n517), .B1(new_n897), .B2(new_n649), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n916), .A2(KEYINPUT42), .B1(new_n626), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n601), .B1(new_n600), .B2(new_n626), .ZN(new_n920));
  OR3_X1    g0720(.A1(new_n594), .A2(new_n600), .A3(new_n626), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n917), .A2(new_n919), .B1(KEYINPUT43), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n923), .B(new_n924), .Z(new_n925));
  NOR3_X1   g0725(.A1(new_n630), .A2(new_n634), .A3(new_n900), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n925), .B(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n920), .A2(new_n711), .A3(new_n921), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n239), .A2(new_n702), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n713), .B1(new_n217), .B2(new_n384), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n699), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n739), .A2(G68), .ZN(new_n932));
  INV_X1    g0732(.A(G150), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n932), .B1(new_n792), .B2(new_n747), .C1(new_n933), .C2(new_n727), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT110), .Z(new_n935));
  OAI22_X1  g0735(.A1(new_n729), .A2(new_n253), .B1(new_n721), .B2(new_n220), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n300), .B1(new_n201), .B2(new_n718), .C1(new_n779), .C2(new_n737), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n936), .B(new_n937), .C1(G137), .C2(new_n735), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n296), .B1(new_n751), .B2(new_n718), .C1(new_n779), .C2(new_n744), .ZN(new_n939));
  INV_X1    g0739(.A(G317), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT46), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n728), .A2(G116), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n736), .A2(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n939), .B(new_n943), .C1(new_n941), .C2(new_n942), .ZN(new_n944));
  XOR2_X1   g0744(.A(KEYINPUT109), .B(G311), .Z(new_n945));
  AOI22_X1  g0745(.A1(new_n724), .A2(new_n945), .B1(G97), .B2(new_n720), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n750), .B2(new_n727), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(G107), .B2(new_n739), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n935), .A2(new_n938), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT47), .Z(new_n950));
  AOI21_X1  g0750(.A(new_n931), .B1(new_n950), .B2(new_n712), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n915), .A2(new_n927), .B1(new_n928), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(G387));
  INV_X1    g0753(.A(new_n645), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n954), .A2(new_n706), .B1(new_n494), .B2(new_n642), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n235), .A2(new_n279), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n257), .A2(new_n269), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT50), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n645), .B(new_n279), .C1(new_n323), .C2(new_n405), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n702), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n955), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n698), .B1(new_n961), .B2(new_n713), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n576), .A2(new_n739), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n300), .B1(new_n323), .B2(new_n718), .C1(new_n779), .C2(new_n311), .ZN(new_n964));
  XNOR2_X1  g0764(.A(KEYINPUT111), .B(G150), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n964), .B1(new_n735), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n729), .A2(new_n220), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(G97), .B2(new_n720), .ZN(new_n968));
  AOI22_X1  g0768(.A1(G50), .A2(new_n726), .B1(new_n724), .B2(G159), .ZN(new_n969));
  AND4_X1   g0769(.A1(new_n963), .A2(new_n966), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n736), .A2(new_n748), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n296), .B1(new_n721), .B2(new_n462), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n756), .A2(G303), .B1(new_n731), .B2(new_n945), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n973), .B1(new_n727), .B2(new_n940), .C1(new_n746), .C2(new_n747), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT48), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n975), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n739), .A2(G283), .B1(G294), .B2(new_n728), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n971), .B(new_n972), .C1(new_n980), .C2(KEYINPUT49), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n980), .A2(KEYINPUT49), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n970), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n962), .B1(new_n983), .B2(new_n778), .C1(new_n636), .C2(new_n762), .ZN(new_n984));
  INV_X1    g0784(.A(new_n910), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n691), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n643), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n691), .A2(new_n985), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n984), .B1(new_n694), .B2(new_n910), .C1(new_n987), .C2(new_n988), .ZN(G393));
  OAI221_X1 g0789(.A(new_n713), .B1(new_n458), .B2(new_n217), .C1(new_n243), .C2(new_n703), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n699), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT112), .Z(new_n992));
  OAI221_X1 g0792(.A(new_n296), .B1(new_n744), .B2(new_n718), .C1(new_n779), .C2(new_n750), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n722), .B(new_n993), .C1(G283), .C2(new_n728), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G311), .A2(new_n726), .B1(new_n724), .B2(G317), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT52), .Z(new_n996));
  NAND2_X1  g0796(.A1(new_n739), .A2(G116), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n735), .A2(G322), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n994), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G150), .A2(new_n724), .B1(new_n726), .B2(G159), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT114), .ZN(new_n1001));
  XOR2_X1   g0801(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n739), .A2(G77), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n735), .A2(G143), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n300), .B1(new_n311), .B2(new_n718), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n729), .A2(new_n323), .B1(new_n721), .B2(new_n345), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n201), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1006), .B(new_n1007), .C1(new_n1008), .C2(new_n731), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .A4(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n999), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n992), .B1(new_n1012), .B2(new_n712), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n899), .B2(new_n762), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n908), .B2(new_n694), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n908), .A2(new_n986), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1016), .A2(new_n644), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n908), .A2(new_n986), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(G390));
  NAND2_X1  g0820(.A1(new_n771), .A2(new_n394), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n626), .B(new_n1021), .C1(new_n650), .C2(new_n655), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n863), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n873), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n846), .B1(new_n842), .B2(new_n829), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT115), .ZN(new_n1026));
  AND3_X1   g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1026), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n845), .A2(new_n849), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT116), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n864), .B2(new_n846), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n862), .A2(new_n863), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n873), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n846), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1034), .A2(KEYINPUT116), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1029), .B1(new_n1030), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n875), .A2(new_n871), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(KEYINPUT117), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n688), .A2(G330), .A3(new_n772), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n873), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1039), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT117), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1037), .B1(new_n849), .B2(new_n845), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1047), .B(new_n1040), .C1(new_n1048), .C2(new_n1029), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1042), .A2(new_n1046), .A3(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1050), .A2(new_n694), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1030), .A2(new_n709), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n776), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n699), .B1(new_n257), .B2(new_n1053), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n462), .A2(new_n727), .B1(new_n747), .B2(new_n751), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n788), .B(new_n1055), .C1(G87), .C2(new_n728), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n735), .A2(G294), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n296), .B1(new_n779), .B2(new_n494), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G97), .B2(new_n756), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1056), .A2(new_n1004), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n300), .B1(new_n721), .B2(new_n201), .ZN(new_n1061));
  INV_X1    g0861(.A(G132), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n727), .A2(new_n1062), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1061), .B(new_n1063), .C1(G128), .C2(new_n724), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n739), .A2(G159), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n728), .A2(new_n965), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(KEYINPUT53), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(KEYINPUT54), .B(G143), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n756), .A2(new_n1069), .B1(new_n731), .B2(G137), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(KEYINPUT118), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .A4(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n735), .A2(G125), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(KEYINPUT53), .B2(new_n1066), .C1(KEYINPUT118), .C2(new_n1070), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1060), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1054), .B1(new_n1075), .B2(new_n712), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1051), .B1(new_n1052), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n439), .A2(G330), .A3(new_n874), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1078), .B(new_n617), .C1(new_n662), .C2(new_n867), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n1041), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n1033), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n874), .A2(G330), .A3(new_n772), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1023), .B1(new_n1083), .B2(new_n1044), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1045), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1079), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1050), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1042), .A2(new_n1046), .A3(new_n1049), .A4(new_n1086), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1088), .A2(new_n643), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1077), .A2(new_n1090), .ZN(G378));
  NAND2_X1  g0891(.A1(new_n310), .A2(new_n374), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n274), .A2(new_n624), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT55), .Z(new_n1094));
  XNOR2_X1  g0894(.A(new_n1092), .B(new_n1094), .ZN(new_n1095));
  XOR2_X1   g0895(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1096));
  XOR2_X1   g0896(.A(new_n1095), .B(new_n1096), .Z(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n876), .A2(G330), .A3(new_n878), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n850), .A2(new_n865), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1099), .B1(new_n850), .B2(new_n865), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1098), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1102), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1104), .A2(new_n1100), .A3(new_n1097), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1098), .A2(new_n709), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n699), .B1(new_n1008), .B2(new_n1053), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n249), .B(new_n275), .C1(new_n721), .C2(new_n737), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n779), .A2(new_n1062), .B1(new_n793), .B2(new_n718), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n728), .B2(new_n1069), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(G125), .A2(new_n724), .B1(new_n726), .B2(G128), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1111), .B(new_n1112), .C1(new_n933), .C2(new_n743), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1113), .A2(KEYINPUT59), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1109), .B(new_n1114), .C1(G124), .C2(new_n735), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(KEYINPUT59), .B2(new_n1113), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n721), .A2(new_n253), .ZN(new_n1117));
  NOR4_X1   g0917(.A1(new_n967), .A2(new_n1117), .A3(new_n447), .A4(new_n300), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n751), .B2(new_n736), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n726), .A2(G107), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT120), .Z(new_n1122));
  NAND2_X1  g0922(.A1(new_n576), .A2(new_n756), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n724), .A2(G116), .B1(G97), .B2(new_n731), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1123), .A2(new_n932), .A3(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1120), .A2(new_n1122), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT58), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  OR2_X1    g0928(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n269), .B1(G33), .B2(G41), .C1(new_n447), .C2(new_n300), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1116), .A2(new_n1128), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1108), .B1(new_n1131), .B2(new_n712), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1106), .A2(new_n695), .B1(new_n1107), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1079), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1089), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT122), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1089), .A2(KEYINPUT122), .A3(new_n1134), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(KEYINPUT57), .B1(new_n1139), .B2(new_n1106), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1103), .A2(new_n1105), .A3(KEYINPUT57), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1089), .A2(KEYINPUT122), .A3(new_n1134), .ZN(new_n1142));
  AOI21_X1  g0942(.A(KEYINPUT122), .B1(new_n1089), .B2(new_n1134), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n643), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1133), .B1(new_n1140), .B2(new_n1145), .ZN(G375));
  NAND3_X1  g0946(.A1(new_n1082), .A2(new_n1079), .A3(new_n1085), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1087), .A2(new_n913), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n694), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n873), .A2(new_n710), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1150), .A2(KEYINPUT123), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(KEYINPUT123), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n1062), .A2(new_n747), .B1(new_n727), .B2(new_n793), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1117), .B(new_n1153), .C1(G159), .C2(new_n728), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n300), .B1(new_n718), .B2(new_n933), .C1(new_n779), .C2(new_n1068), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G128), .B2(new_n735), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1154), .B(new_n1156), .C1(new_n269), .C2(new_n743), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n747), .A2(new_n744), .B1(new_n458), .B2(new_n729), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n727), .A2(new_n751), .B1(new_n405), .B2(new_n721), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n735), .A2(G303), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n296), .B1(new_n718), .B2(new_n494), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G116), .B2(new_n731), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1160), .A2(new_n963), .A3(new_n1161), .A4(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n778), .B1(new_n1157), .B2(new_n1164), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n698), .B(new_n1165), .C1(new_n323), .C2(new_n776), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT124), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n1151), .A2(new_n1152), .A3(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1149), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1148), .A2(new_n1169), .ZN(G381));
  OR4_X1    g0970(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1171), .A2(G387), .A3(G381), .ZN(new_n1172));
  INV_X1    g0972(.A(G378), .ZN(new_n1173));
  INV_X1    g0973(.A(G375), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(G407));
  NOR2_X1   g0975(.A1(new_n622), .A2(G343), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1173), .A3(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(G407), .A2(G213), .A3(new_n1177), .ZN(G409));
  OAI211_X1 g0978(.A(G378), .B(new_n1133), .C1(new_n1140), .C2(new_n1145), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n913), .B(new_n1106), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n1133), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n1173), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1176), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1147), .A2(KEYINPUT125), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT60), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1147), .A2(KEYINPUT125), .A3(KEYINPUT60), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n644), .B(new_n1086), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1169), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n800), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1193), .A2(new_n643), .A3(new_n1087), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1194), .A2(G384), .A3(new_n1169), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1192), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1176), .A2(G2897), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1196), .A2(G2897), .A3(new_n1176), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT61), .B1(new_n1185), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT63), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n1185), .B2(new_n1196), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(G393), .B(new_n764), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G387), .B2(KEYINPUT126), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1206), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n952), .A2(new_n1208), .ZN(new_n1209));
  OR3_X1    g1009(.A1(new_n1207), .A2(new_n1019), .A3(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1019), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1176), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1213), .A2(KEYINPUT63), .A3(new_n1197), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1203), .A2(new_n1205), .A3(new_n1212), .A4(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT62), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1213), .A2(new_n1216), .A3(new_n1197), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT61), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n1213), .B2(new_n1201), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1216), .B1(new_n1213), .B2(new_n1197), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(new_n1217), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1215), .B1(new_n1221), .B2(new_n1212), .ZN(G405));
  NAND3_X1  g1022(.A1(G375), .A2(new_n1197), .A3(new_n1173), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1197), .B1(G375), .B2(new_n1173), .ZN(new_n1225));
  OAI211_X1 g1025(.A(KEYINPUT127), .B(new_n1179), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1225), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1179), .A2(KEYINPUT127), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n1229), .A3(new_n1223), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1226), .A2(new_n1227), .A3(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1227), .B1(new_n1226), .B2(new_n1230), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(G402));
endmodule


