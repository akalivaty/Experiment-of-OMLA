//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT25), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  INV_X1    g003(.A(G176gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AND2_X1   g005(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n207));
  NOR2_X1   g006(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT66), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n206), .B(new_n211), .C1(new_n207), .C2(new_n208), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n204), .A2(new_n205), .A3(KEYINPUT23), .ZN(new_n213));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT67), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n213), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  AOI22_X1  g017(.A1(new_n210), .A2(new_n212), .B1(new_n218), .B2(KEYINPUT68), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n213), .A2(new_n216), .A3(new_n217), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT68), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n222));
  INV_X1    g021(.A(G183gat), .ZN(new_n223));
  INV_X1    g022(.A(G190gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n220), .A2(new_n221), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n203), .B1(new_n219), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n210), .A2(new_n212), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n203), .A3(new_n214), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n230), .B1(new_n226), .B2(new_n225), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n223), .A2(KEYINPUT27), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT27), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G183gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n235), .A3(new_n224), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT28), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT27), .B(G183gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(KEYINPUT28), .A3(new_n224), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n204), .A2(new_n205), .A3(KEYINPUT26), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT26), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n243), .B1(G169gat), .B2(G176gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n245), .A2(new_n214), .B1(G183gat), .B2(G190gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n228), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n250));
  INV_X1    g049(.A(G134gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G127gat), .ZN(new_n252));
  INV_X1    g051(.A(G127gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G134gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G113gat), .B(G120gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n255), .B1(new_n256), .B2(KEYINPUT1), .ZN(new_n257));
  INV_X1    g056(.A(G120gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G113gat), .ZN(new_n259));
  INV_X1    g058(.A(G113gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G120gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G127gat), .B(G134gat), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT1), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n257), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n249), .A2(new_n250), .A3(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n213), .A2(new_n216), .A3(KEYINPUT68), .A4(new_n217), .ZN(new_n268));
  INV_X1    g067(.A(new_n212), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT65), .B(KEYINPUT23), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n211), .B1(new_n270), .B2(new_n206), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n268), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n225), .A2(new_n226), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(new_n218), .B2(KEYINPUT68), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT25), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n229), .A2(new_n231), .B1(new_n241), .B2(new_n246), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n257), .A2(new_n265), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT69), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT70), .B1(new_n277), .B2(new_n278), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n281));
  AOI211_X1 g080(.A(new_n281), .B(new_n266), .C1(new_n275), .C2(new_n276), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n267), .B(new_n279), .C1(new_n280), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G227gat), .A2(G233gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT34), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT71), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n288), .B(KEYINPUT34), .C1(new_n283), .C2(new_n285), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n284), .B(KEYINPUT64), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n290), .A2(KEYINPUT34), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n283), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n287), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT33), .B1(new_n283), .B2(new_n290), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT32), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n296), .B1(new_n283), .B2(new_n290), .ZN(new_n297));
  XOR2_X1   g096(.A(G15gat), .B(G43gat), .Z(new_n298));
  XNOR2_X1  g097(.A(G71gat), .B(G99gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NOR3_X1   g100(.A1(new_n295), .A2(new_n297), .A3(new_n301), .ZN(new_n302));
  AOI221_X4 g101(.A(new_n296), .B1(KEYINPUT33), .B2(new_n300), .C1(new_n283), .C2(new_n290), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n294), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n283), .A2(new_n290), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT33), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(KEYINPUT32), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n308), .A3(new_n300), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n297), .B1(new_n295), .B2(new_n301), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n292), .B1(new_n286), .B2(KEYINPUT71), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n309), .A2(new_n310), .B1(new_n311), .B2(new_n289), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n202), .B1(new_n304), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(G155gat), .A2(G162gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G148gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G141gat), .ZN(new_n318));
  INV_X1    g117(.A(G141gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G148gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT2), .ZN(new_n322));
  AOI211_X1 g121(.A(new_n314), .B(new_n316), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n317), .A2(KEYINPUT73), .A3(G141gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT73), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n326), .B1(new_n319), .B2(G148gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n319), .A2(G148gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n325), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n314), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n315), .B1(new_n330), .B2(KEYINPUT2), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n329), .A2(KEYINPUT74), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT74), .B1(new_n329), .B2(new_n331), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n324), .B(new_n266), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT78), .B1(new_n334), .B2(KEYINPUT4), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(KEYINPUT4), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n334), .A2(KEYINPUT78), .A3(KEYINPUT4), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n278), .A2(KEYINPUT75), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n341), .B1(new_n257), .B2(new_n265), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n317), .A2(KEYINPUT73), .A3(G141gat), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT73), .B1(new_n317), .B2(G141gat), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n346), .B1(new_n318), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n316), .B1(new_n322), .B2(new_n314), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n329), .A2(KEYINPUT74), .A3(new_n331), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n323), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT3), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n324), .B1(new_n332), .B2(new_n333), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT3), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n344), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G225gat), .A2(G233gat), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n359), .A2(KEYINPUT5), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n339), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n352), .A2(new_n362), .A3(new_n266), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n336), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n357), .A2(new_n364), .A3(new_n358), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT5), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n334), .B1(new_n343), .B2(new_n352), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n366), .B1(new_n367), .B2(new_n359), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n361), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G57gat), .B(G85gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n371), .B(KEYINPUT77), .ZN(new_n372));
  XOR2_X1   g171(.A(G1gat), .B(G29gat), .Z(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n370), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT6), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G8gat), .B(G36gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(G64gat), .B(G92gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  XOR2_X1   g184(.A(G211gat), .B(G218gat), .Z(new_n386));
  INV_X1    g185(.A(G218gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT72), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT72), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(G218gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT22), .B1(new_n391), .B2(G211gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(G197gat), .B(G204gat), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n386), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n386), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT72), .B(G218gat), .ZN(new_n397));
  INV_X1    g196(.A(G211gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n393), .B(new_n396), .C1(new_n399), .C2(KEYINPUT22), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G226gat), .A2(G233gat), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(new_n249), .B2(KEYINPUT29), .ZN(new_n404));
  INV_X1    g203(.A(new_n403), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n405), .B1(new_n228), .B2(new_n248), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n402), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT29), .B1(new_n275), .B2(new_n276), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n406), .B(new_n402), .C1(new_n408), .C2(new_n405), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n385), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n406), .B1(new_n408), .B2(new_n405), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n401), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n413), .A2(new_n384), .A3(new_n409), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(KEYINPUT30), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n384), .B1(new_n413), .B2(new_n409), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT30), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n361), .A2(new_n369), .A3(new_n376), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT79), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT79), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n361), .A2(new_n369), .A3(new_n422), .A4(new_n376), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT6), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n381), .B(new_n419), .C1(new_n424), .C2(new_n379), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n294), .B1(new_n302), .B2(new_n303), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n309), .A2(new_n289), .A3(new_n311), .A4(new_n310), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n428), .A3(KEYINPUT84), .ZN(new_n429));
  NAND2_X1  g228(.A1(G228gat), .A2(G233gat), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT29), .B1(new_n395), .B2(new_n400), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n355), .B1(new_n431), .B2(KEYINPUT3), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT80), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n430), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT29), .B1(new_n352), .B2(new_n353), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n432), .B1(new_n435), .B2(new_n401), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  OAI221_X1 g236(.A(new_n432), .B1(new_n433), .B2(new_n430), .C1(new_n435), .C2(new_n401), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(G22gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT81), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n437), .A2(G22gat), .A3(new_n438), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G78gat), .B(G106gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT31), .B(G50gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n443), .A2(new_n445), .A3(new_n449), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n441), .B(new_n444), .C1(new_n442), .C2(new_n448), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT35), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n313), .A2(new_n426), .A3(new_n429), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n451), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n427), .A2(new_n454), .A3(new_n428), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n426), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n453), .A2(KEYINPUT85), .B1(KEYINPUT35), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n429), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT84), .B1(new_n427), .B2(new_n428), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT85), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n460), .A2(new_n461), .A3(new_n426), .A4(new_n452), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n378), .A2(KEYINPUT6), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n343), .B1(KEYINPUT3), .B2(new_n355), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n337), .A2(new_n338), .B1(new_n464), .B2(new_n354), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n465), .A2(new_n360), .B1(new_n365), .B2(new_n368), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n422), .B1(new_n466), .B2(new_n376), .ZN(new_n467));
  INV_X1    g266(.A(new_n423), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n380), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n463), .B1(new_n469), .B2(new_n378), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT37), .B1(new_n407), .B2(new_n410), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT37), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n413), .A2(new_n473), .A3(new_n409), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n385), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT38), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n471), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n416), .B1(new_n475), .B2(new_n476), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n413), .A2(new_n473), .A3(new_n409), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n473), .B1(new_n413), .B2(new_n409), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n384), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(KEYINPUT83), .A3(KEYINPUT38), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n477), .A2(new_n478), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n470), .A2(new_n483), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n415), .A2(new_n418), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n378), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n367), .A2(new_n359), .ZN(new_n487));
  OAI211_X1 g286(.A(KEYINPUT39), .B(new_n487), .C1(new_n465), .C2(new_n358), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT39), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n334), .A2(KEYINPUT78), .A3(KEYINPUT4), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n490), .B1(new_n336), .B2(new_n335), .ZN(new_n491));
  INV_X1    g290(.A(new_n357), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n489), .B(new_n359), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT82), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n493), .A2(new_n494), .A3(new_n376), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n494), .B1(new_n493), .B2(new_n376), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n488), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT40), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT40), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n499), .B(new_n488), .C1(new_n495), .C2(new_n496), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n486), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n454), .B1(new_n484), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n454), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n426), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n427), .A2(new_n428), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT36), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n457), .A2(new_n462), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT89), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT16), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(G1gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(G15gat), .B(G22gat), .ZN(new_n513));
  MUX2_X1   g312(.A(G1gat), .B(new_n512), .S(new_n513), .Z(new_n514));
  XOR2_X1   g313(.A(new_n514), .B(G8gat), .Z(new_n515));
  NOR3_X1   g314(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT86), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g318(.A(KEYINPUT86), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n521), .A2(KEYINPUT88), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(KEYINPUT88), .ZN(new_n523));
  INV_X1    g322(.A(G50gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(G43gat), .ZN(new_n525));
  INV_X1    g324(.A(G43gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(G50gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT87), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT15), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n525), .B(new_n527), .C1(new_n529), .C2(KEYINPUT15), .ZN(new_n533));
  INV_X1    g332(.A(G29gat), .ZN(new_n534));
  INV_X1    g333(.A(G36gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n532), .A2(new_n533), .A3(new_n537), .ZN(new_n538));
  OR3_X1    g337(.A1(new_n522), .A2(new_n523), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n521), .A2(new_n536), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n540), .A2(new_n531), .A3(new_n528), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT17), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n539), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n522), .A2(new_n523), .A3(new_n538), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT17), .B1(new_n545), .B2(new_n541), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n515), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n545), .A2(new_n541), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n514), .B(G8gat), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G229gat), .A2(G233gat), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NOR3_X1   g351(.A1(new_n547), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n510), .B1(new_n553), .B2(KEYINPUT18), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n544), .A2(new_n546), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n549), .ZN(new_n556));
  INV_X1    g355(.A(new_n550), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT18), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(KEYINPUT89), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n556), .A2(KEYINPUT18), .A3(new_n551), .A4(new_n557), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n548), .B(new_n549), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n551), .B(KEYINPUT13), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G113gat), .B(G141gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT11), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(new_n204), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(G197gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT12), .ZN(new_n571));
  INV_X1    g370(.A(G197gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n569), .B(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT12), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n561), .A2(new_n566), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n558), .A2(new_n559), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n566), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n576), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n509), .A2(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(G183gat), .B(G211gat), .Z(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  OR2_X1    g385(.A1(G57gat), .A2(G64gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(G57gat), .A2(G64gat), .ZN(new_n588));
  AND2_X1   g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n587), .B(new_n588), .C1(new_n589), .C2(KEYINPUT9), .ZN(new_n590));
  XOR2_X1   g389(.A(G71gat), .B(G78gat), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT21), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G127gat), .B(G155gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n592), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n515), .B1(KEYINPUT21), .B2(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n602), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n586), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n603), .A2(new_n604), .A3(new_n586), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G134gat), .B(G162gat), .Z(new_n609));
  NAND2_X1  g408(.A1(G85gat), .A2(G92gat), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT90), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT7), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n610), .B(KEYINPUT90), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT7), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G99gat), .A2(G106gat), .ZN(new_n617));
  INV_X1    g416(.A(G85gat), .ZN(new_n618));
  INV_X1    g417(.A(G92gat), .ZN(new_n619));
  AOI22_X1  g418(.A1(KEYINPUT8), .A2(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n613), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G99gat), .B(G106gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n613), .A2(new_n616), .A3(new_n622), .A4(new_n620), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n627), .B1(new_n544), .B2(new_n546), .ZN(new_n628));
  AND2_X1   g427(.A1(G232gat), .A2(G233gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT41), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n630), .B1(new_n548), .B2(new_n626), .ZN(new_n631));
  XNOR2_X1  g430(.A(G190gat), .B(G218gat), .ZN(new_n632));
  OR3_X1    g431(.A1(new_n628), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n629), .A2(KEYINPUT41), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n632), .B1(new_n628), .B2(new_n631), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n635), .B1(new_n633), .B2(new_n636), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n609), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n639), .ZN(new_n641));
  INV_X1    g440(.A(new_n609), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n641), .A2(new_n637), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n608), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT10), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n625), .A2(KEYINPUT91), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n624), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n621), .A2(KEYINPUT91), .A3(new_n623), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n592), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n626), .A2(new_n601), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n647), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n624), .A2(new_n601), .A3(KEYINPUT10), .A4(new_n625), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT92), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(G230gat), .A2(G233gat), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OR3_X1    g457(.A1(new_n651), .A2(new_n652), .A3(new_n657), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G120gat), .B(G148gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(G176gat), .B(G204gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n663), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n658), .A2(new_n659), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n646), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n584), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n470), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT93), .B(G1gat), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1324gat));
  INV_X1    g472(.A(KEYINPUT94), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT16), .B(G8gat), .Z(new_n675));
  NAND3_X1  g474(.A1(new_n669), .A2(new_n485), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n584), .A2(new_n485), .A3(new_n668), .ZN(new_n679));
  INV_X1    g478(.A(new_n675), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n681), .A2(KEYINPUT94), .A3(KEYINPUT42), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n679), .A2(G8gat), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n684), .A2(KEYINPUT95), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(KEYINPUT95), .ZN(new_n686));
  OAI22_X1  g485(.A1(new_n685), .A2(new_n686), .B1(new_n677), .B2(new_n676), .ZN(new_n687));
  OR3_X1    g486(.A1(new_n683), .A2(new_n687), .A3(KEYINPUT96), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT96), .B1(new_n683), .B2(new_n687), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(G1325gat));
  INV_X1    g489(.A(new_n669), .ZN(new_n691));
  OAI21_X1  g490(.A(G15gat), .B1(new_n691), .B2(new_n508), .ZN(new_n692));
  INV_X1    g491(.A(new_n460), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(G15gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n691), .B2(new_n694), .ZN(G1326gat));
  NAND2_X1  g494(.A1(new_n669), .A2(new_n503), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT97), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT43), .B(G22gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  OAI21_X1  g498(.A(KEYINPUT44), .B1(new_n509), .B2(new_n645), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n457), .A2(new_n462), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n505), .A2(new_n508), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n645), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT99), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT99), .ZN(new_n706));
  NOR4_X1   g505(.A1(new_n509), .A2(new_n706), .A3(KEYINPUT44), .A4(new_n645), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n700), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n608), .A2(KEYINPUT98), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT98), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n606), .A2(new_n710), .A3(new_n607), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n712), .A2(new_n583), .A3(new_n667), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n708), .A2(new_n670), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT100), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n708), .A2(KEYINPUT100), .A3(new_n670), .A4(new_n713), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n716), .A2(G29gat), .A3(new_n717), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n608), .A2(new_n645), .A3(new_n667), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n584), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n721), .A2(new_n534), .A3(new_n670), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT45), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT101), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n718), .A2(KEYINPUT101), .A3(new_n723), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1328gat));
  NOR3_X1   g527(.A1(new_n720), .A2(G36gat), .A3(new_n419), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT46), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n708), .A2(new_n485), .A3(new_n713), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n731), .B2(new_n535), .ZN(G1329gat));
  NAND4_X1  g531(.A1(new_n708), .A2(G43gat), .A3(new_n507), .A4(new_n713), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n720), .A2(new_n693), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(G43gat), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g535(.A1(new_n708), .A2(G50gat), .A3(new_n503), .A4(new_n713), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n524), .B1(new_n720), .B2(new_n454), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g539(.A1(new_n701), .A2(new_n702), .ZN(new_n741));
  INV_X1    g540(.A(new_n667), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n646), .A2(new_n582), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n470), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT102), .B(G57gat), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1332gat));
  INV_X1    g546(.A(new_n744), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT49), .ZN(new_n749));
  INV_X1    g548(.A(G64gat), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n485), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT103), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n749), .A2(new_n750), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1333gat));
  NAND3_X1  g554(.A1(new_n748), .A2(G71gat), .A3(new_n507), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n744), .A2(new_n693), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(G71gat), .B2(new_n757), .ZN(new_n758));
  XOR2_X1   g557(.A(KEYINPUT104), .B(KEYINPUT50), .Z(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1334gat));
  NAND2_X1  g559(.A1(new_n748), .A2(new_n503), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g561(.A1(new_n608), .A2(new_n582), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n703), .B(new_n763), .C1(KEYINPUT106), .C2(KEYINPUT51), .ZN(new_n764));
  NAND2_X1  g563(.A1(KEYINPUT106), .A2(KEYINPUT51), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(KEYINPUT107), .Z(new_n767));
  NAND3_X1  g566(.A1(new_n670), .A2(new_n618), .A3(new_n667), .ZN(new_n768));
  INV_X1    g567(.A(new_n708), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n763), .A2(new_n667), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT105), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n769), .A2(new_n470), .A3(new_n771), .ZN(new_n772));
  OAI22_X1  g571(.A1(new_n767), .A2(new_n768), .B1(new_n618), .B2(new_n772), .ZN(G1336gat));
  NAND4_X1  g572(.A1(new_n766), .A2(new_n619), .A3(new_n485), .A4(new_n667), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n769), .A2(new_n419), .A3(new_n771), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n775), .B2(new_n619), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT52), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n774), .B(new_n778), .C1(new_n775), .C2(new_n619), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1337gat));
  INV_X1    g579(.A(G99gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n460), .A2(new_n781), .A3(new_n667), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n769), .A2(new_n508), .A3(new_n771), .ZN(new_n783));
  OAI22_X1  g582(.A1(new_n767), .A2(new_n782), .B1(new_n781), .B2(new_n783), .ZN(G1338gat));
  INV_X1    g583(.A(G106gat), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n766), .A2(new_n785), .A3(new_n503), .A4(new_n667), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n769), .A2(new_n454), .A3(new_n771), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n787), .B2(new_n785), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT53), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n786), .B(new_n790), .C1(new_n787), .C2(new_n785), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(G1339gat));
  INV_X1    g591(.A(new_n712), .ZN(new_n793));
  INV_X1    g592(.A(new_n657), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n653), .A2(new_n655), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT108), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT108), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n653), .A2(new_n655), .A3(new_n797), .A4(new_n794), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n794), .B1(new_n653), .B2(new_n655), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n665), .B1(new_n800), .B2(new_n801), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n803), .A2(KEYINPUT55), .A3(new_n804), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n807), .A2(new_n582), .A3(new_n666), .A4(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n562), .A2(new_n576), .A3(new_n565), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n554), .B2(new_n560), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n563), .A2(new_n564), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n552), .B1(new_n547), .B2(new_n550), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n573), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n667), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n644), .B1(new_n809), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n644), .A2(new_n807), .A3(new_n815), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n808), .A2(new_n666), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT109), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n817), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n663), .B1(new_n658), .B2(KEYINPUT54), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n799), .B2(new_n802), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n576), .B1(new_n566), .B2(new_n578), .ZN(new_n825));
  OAI22_X1  g624(.A1(new_n824), .A2(KEYINPUT55), .B1(new_n825), .B2(new_n811), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n816), .B1(new_n826), .B2(new_n819), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n645), .ZN(new_n828));
  INV_X1    g627(.A(new_n819), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n829), .A2(new_n644), .A3(new_n815), .A4(new_n807), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT109), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n793), .B1(new_n822), .B2(new_n831), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n646), .A2(new_n582), .A3(new_n667), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(KEYINPUT110), .A3(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT110), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n821), .B1(new_n817), .B2(new_n820), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n828), .A2(KEYINPUT109), .A3(new_n830), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n712), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n836), .B1(new_n839), .B2(new_n833), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n835), .A2(new_n840), .A3(new_n670), .A4(new_n455), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n485), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT112), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n841), .A2(KEYINPUT112), .A3(new_n485), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n260), .B(new_n582), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n835), .A2(new_n840), .A3(new_n454), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT111), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n835), .A2(new_n840), .A3(KEYINPUT111), .A4(new_n454), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n670), .A2(new_n419), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n693), .A2(new_n852), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n851), .A2(new_n582), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n846), .B1(new_n260), .B2(new_n854), .ZN(G1340gat));
  NAND2_X1  g654(.A1(new_n667), .A2(new_n258), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT113), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n857), .B1(new_n844), .B2(new_n845), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n851), .A2(new_n667), .A3(new_n853), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n258), .B2(new_n859), .ZN(G1341gat));
  NAND4_X1  g659(.A1(new_n851), .A2(G127gat), .A3(new_n712), .A4(new_n853), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n842), .A2(KEYINPUT114), .A3(new_n608), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n253), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT114), .B1(new_n842), .B2(new_n608), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT115), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n867), .B(new_n861), .C1(new_n863), .C2(new_n864), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n868), .ZN(G1342gat));
  NOR2_X1   g668(.A1(new_n645), .A2(new_n485), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n841), .A2(G134gat), .A3(new_n871), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT56), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n851), .A2(new_n644), .A3(new_n853), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(new_n251), .ZN(G1343gat));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n835), .A2(new_n840), .A3(new_n876), .A4(new_n503), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n608), .B1(new_n828), .B2(new_n830), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n503), .B1(new_n833), .B2(new_n878), .ZN(new_n879));
  AOI211_X1 g678(.A(new_n507), .B(new_n852), .C1(new_n879), .C2(KEYINPUT57), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(G141gat), .B1(new_n881), .B2(new_n583), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT58), .B1(new_n882), .B2(KEYINPUT118), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n835), .A2(new_n840), .A3(new_n670), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n835), .A2(new_n840), .A3(KEYINPUT116), .A4(new_n670), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n507), .A2(new_n454), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n886), .A2(new_n419), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n582), .A2(new_n319), .ZN(new_n890));
  XOR2_X1   g689(.A(new_n890), .B(KEYINPUT117), .Z(new_n891));
  OAI21_X1  g690(.A(new_n882), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  XOR2_X1   g691(.A(new_n883), .B(new_n892), .Z(G1344gat));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n894), .B(G148gat), .C1(new_n881), .C2(new_n742), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n835), .A2(new_n840), .A3(KEYINPUT57), .A4(new_n503), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n828), .A2(new_n830), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n897), .A2(KEYINPUT119), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n608), .B1(new_n897), .B2(KEYINPUT119), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n833), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n876), .B1(new_n900), .B2(new_n454), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  OR3_X1    g701(.A1(new_n507), .A2(new_n742), .A3(new_n852), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n317), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n895), .B1(new_n905), .B2(new_n894), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n667), .A2(new_n317), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n889), .B2(new_n907), .ZN(G1345gat));
  OAI21_X1  g707(.A(G155gat), .B1(new_n881), .B2(new_n793), .ZN(new_n909));
  INV_X1    g708(.A(new_n608), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n910), .A2(G155gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n909), .B1(new_n889), .B2(new_n911), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(KEYINPUT120), .Z(G1346gat));
  OAI21_X1  g712(.A(G162gat), .B1(new_n881), .B2(new_n645), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n871), .A2(G162gat), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n886), .A2(new_n887), .A3(new_n888), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1347gat));
  AND4_X1   g716(.A1(new_n470), .A2(new_n835), .A3(new_n840), .A4(new_n485), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n455), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n918), .A2(KEYINPUT121), .A3(new_n455), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n921), .A2(new_n582), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n470), .A2(new_n485), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT122), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n925), .A2(new_n693), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n927), .B1(new_n849), .B2(new_n850), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n583), .A2(new_n204), .ZN(new_n929));
  AOI22_X1  g728(.A1(new_n923), .A2(new_n204), .B1(new_n928), .B2(new_n929), .ZN(G1348gat));
  NAND4_X1  g729(.A1(new_n921), .A2(new_n205), .A3(new_n667), .A4(new_n922), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n928), .A2(new_n667), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n932), .B2(new_n205), .ZN(G1349gat));
  NAND3_X1  g732(.A1(new_n851), .A2(new_n712), .A3(new_n926), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G183gat), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n918), .A2(new_n239), .A3(new_n455), .A4(new_n608), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n935), .A2(new_n936), .A3(KEYINPUT60), .A4(new_n937), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n936), .A2(KEYINPUT60), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n936), .A2(KEYINPUT60), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n223), .B1(new_n928), .B2(new_n712), .ZN(new_n941));
  INV_X1    g740(.A(new_n937), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n939), .B(new_n940), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n938), .A2(new_n943), .ZN(G1350gat));
  NAND4_X1  g743(.A1(new_n921), .A2(new_n224), .A3(new_n644), .A4(new_n922), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n928), .A2(new_n644), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n946), .B1(new_n947), .B2(G190gat), .ZN(new_n948));
  AOI211_X1 g747(.A(KEYINPUT61), .B(new_n224), .C1(new_n928), .C2(new_n644), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G1351gat));
  AND2_X1   g749(.A1(new_n918), .A2(new_n888), .ZN(new_n951));
  XOR2_X1   g750(.A(KEYINPUT124), .B(G197gat), .Z(new_n952));
  NOR2_X1   g751(.A1(new_n583), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n925), .A2(new_n507), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n955), .B1(new_n902), .B2(KEYINPUT125), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n896), .A2(new_n957), .A3(new_n901), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT126), .B1(new_n959), .B2(new_n582), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n956), .A2(KEYINPUT126), .A3(new_n582), .A4(new_n958), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(new_n952), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n954), .B1(new_n960), .B2(new_n962), .ZN(G1352gat));
  NAND2_X1  g762(.A1(new_n959), .A2(new_n667), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G204gat), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n742), .A2(G204gat), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n966), .B1(new_n951), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n951), .A2(new_n966), .A3(new_n967), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n951), .A2(KEYINPUT127), .A3(new_n966), .A4(new_n967), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n965), .A2(new_n973), .ZN(G1353gat));
  NOR2_X1   g773(.A1(new_n955), .A2(new_n910), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n398), .B1(new_n902), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT63), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n951), .A2(new_n398), .A3(new_n608), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(G1354gat));
  AOI21_X1  g778(.A(G218gat), .B1(new_n951), .B2(new_n644), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n645), .A2(new_n397), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n980), .B1(new_n959), .B2(new_n981), .ZN(G1355gat));
endmodule


