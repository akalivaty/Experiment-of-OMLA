//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT65), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  INV_X1    g0013(.A(new_n206), .ZN(new_n214));
  INV_X1    g0014(.A(G50), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT66), .Z(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G20), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n213), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  AND2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n225), .A2(KEYINPUT67), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(KEYINPUT67), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n229));
  NAND4_X1  g0029(.A1(new_n226), .A2(new_n227), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(new_n210), .ZN(new_n231));
  AND2_X1   g0031(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n233));
  NOR3_X1   g0033(.A1(new_n222), .A2(new_n232), .A3(new_n233), .ZN(G361));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT2), .B(G226), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n238), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n201), .ZN(new_n246));
  XOR2_X1   g0046(.A(KEYINPUT69), .B(G50), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n219), .ZN(new_n254));
  INV_X1    g0054(.A(G20), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n255), .B1(new_n214), .B2(new_n215), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G150), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI22_X1  g0061(.A1(new_n257), .A2(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n254), .B1(new_n256), .B2(new_n262), .ZN(new_n263));
  OR2_X1    g0063(.A1(KEYINPUT71), .A2(G1), .ZN(new_n264));
  NAND2_X1  g0064(.A1(KEYINPUT71), .A2(G1), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n264), .A2(G13), .A3(G20), .A4(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(G50), .ZN(new_n267));
  INV_X1    g0067(.A(new_n265), .ZN(new_n268));
  NOR2_X1   g0068(.A1(KEYINPUT71), .A2(G1), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n254), .B1(new_n270), .B2(G20), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n267), .B1(G50), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(KEYINPUT9), .B1(new_n263), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  INV_X1    g0075(.A(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(G222), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G77), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(G1698), .ZN(new_n283));
  INV_X1    g0083(.A(G223), .ZN(new_n284));
  OAI221_X1 g0084(.A(new_n281), .B1(new_n282), .B2(new_n279), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT73), .B1(new_n287), .B2(new_n219), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT73), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n220), .A2(new_n289), .A3(new_n286), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n264), .A2(new_n265), .ZN(new_n293));
  INV_X1    g0093(.A(G41), .ZN(new_n294));
  INV_X1    g0094(.A(G45), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT72), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT72), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n270), .A2(new_n299), .A3(new_n296), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT70), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(G33), .A3(G41), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n219), .B1(KEYINPUT70), .B2(new_n286), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n298), .A2(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G226), .ZN(new_n305));
  INV_X1    g0105(.A(G274), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(new_n303), .B2(new_n302), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n297), .A2(G1), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n292), .A2(new_n305), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G200), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n292), .A2(new_n305), .A3(G190), .A4(new_n309), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n263), .A2(KEYINPUT9), .A3(new_n272), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n274), .A2(new_n311), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT10), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n310), .A2(G179), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT74), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n263), .A2(new_n272), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n310), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n317), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n315), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n266), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n282), .ZN(new_n324));
  INV_X1    g0124(.A(new_n271), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n324), .B1(new_n325), .B2(new_n282), .ZN(new_n326));
  INV_X1    g0126(.A(new_n254), .ZN(new_n327));
  INV_X1    g0127(.A(new_n257), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n328), .A2(new_n260), .B1(G20), .B2(G77), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT15), .B(G87), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n330), .A2(new_n258), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n327), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n279), .A2(G232), .A3(new_n280), .ZN(new_n334));
  INV_X1    g0134(.A(G107), .ZN(new_n335));
  INV_X1    g0135(.A(G238), .ZN(new_n336));
  OAI221_X1 g0136(.A(new_n334), .B1(new_n335), .B2(new_n279), .C1(new_n283), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n291), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n304), .A2(G244), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(new_n309), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n333), .B1(new_n340), .B2(new_n319), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(G179), .B2(new_n340), .ZN(new_n342));
  INV_X1    g0142(.A(G190), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT75), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n333), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n340), .A2(G200), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n344), .B1(KEYINPUT75), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n342), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n322), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n351), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n352));
  AND2_X1   g0152(.A1(KEYINPUT3), .A2(G33), .ZN(new_n353));
  NOR2_X1   g0153(.A1(KEYINPUT3), .A2(G33), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT77), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT77), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n277), .A2(new_n356), .A3(new_n278), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(new_n357), .A3(new_n255), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT7), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n279), .A2(G20), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT78), .B(KEYINPUT7), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n358), .A2(new_n359), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  OAI211_X1 g0163(.A(KEYINPUT16), .B(new_n352), .C1(new_n363), .C2(new_n202), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT16), .ZN(new_n365));
  INV_X1    g0165(.A(new_n352), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n361), .B1(new_n279), .B2(G20), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n353), .A2(new_n354), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(KEYINPUT7), .A3(new_n255), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n202), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n365), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n364), .A2(new_n371), .A3(new_n254), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n266), .A2(new_n257), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n271), .B2(new_n257), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G33), .A2(G87), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n376), .B(KEYINPUT79), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n284), .A2(new_n280), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(G226), .B2(new_n280), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n377), .B1(new_n368), .B2(new_n379), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n380), .A2(new_n291), .B1(new_n307), .B2(new_n308), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n286), .A2(KEYINPUT70), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n382), .A2(new_n302), .A3(new_n220), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n299), .B1(new_n270), .B2(new_n296), .ZN(new_n384));
  AND4_X1   g0184(.A1(new_n299), .A2(new_n264), .A3(new_n296), .A4(new_n265), .ZN(new_n385));
  OAI211_X1 g0185(.A(G232), .B(new_n383), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G169), .ZN(new_n388));
  INV_X1    g0188(.A(G179), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n388), .B1(new_n389), .B2(new_n387), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n375), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT18), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT18), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n375), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n387), .A2(G200), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n381), .A2(G190), .A3(new_n386), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n372), .A2(new_n395), .A3(new_n374), .A4(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n395), .A2(new_n396), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n400), .A2(KEYINPUT17), .A3(new_n372), .A4(new_n374), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n392), .A2(new_n394), .A3(new_n399), .A4(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n276), .A2(G20), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n404), .A2(G77), .B1(G20), .B2(new_n202), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n215), .B2(new_n261), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n254), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT11), .ZN(new_n408));
  XNOR2_X1  g0208(.A(new_n407), .B(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT12), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n323), .A2(new_n410), .A3(new_n202), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT12), .B1(new_n266), .B2(G68), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n202), .B2(new_n325), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n240), .A2(G1698), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(G226), .B2(G1698), .ZN(new_n418));
  INV_X1    g0218(.A(G97), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n418), .A2(new_n368), .B1(new_n276), .B2(new_n419), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(new_n291), .B1(new_n307), .B2(new_n308), .ZN(new_n421));
  OAI211_X1 g0221(.A(G238), .B(new_n383), .C1(new_n384), .C2(new_n385), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT13), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT13), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n421), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(G179), .A3(new_n426), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n421), .A2(new_n422), .A3(new_n425), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n425), .B1(new_n421), .B2(new_n422), .ZN(new_n429));
  OAI21_X1  g0229(.A(G169), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT76), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT14), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n427), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n424), .A2(new_n426), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n432), .B1(new_n435), .B2(G169), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n416), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(G200), .B1(new_n428), .B2(new_n429), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n424), .A2(G190), .A3(new_n426), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n415), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n350), .A2(new_n403), .A3(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(G264), .B(G1698), .C1(new_n353), .C2(new_n354), .ZN(new_n443));
  OAI211_X1 g0243(.A(G257), .B(new_n280), .C1(new_n353), .C2(new_n354), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n277), .A2(G303), .A3(new_n278), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n446), .A2(new_n291), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n268), .A2(new_n269), .A3(new_n295), .ZN(new_n448));
  AND2_X1   g0248(.A1(KEYINPUT5), .A2(G41), .ZN(new_n449));
  NOR2_X1   g0249(.A1(KEYINPUT5), .A2(G41), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n448), .A2(new_n383), .A3(new_n451), .A4(G274), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n264), .A2(G45), .A3(new_n265), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n449), .A2(new_n450), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n383), .B(G270), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n447), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G190), .ZN(new_n458));
  INV_X1    g0258(.A(G116), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n270), .A2(G13), .A3(G20), .A4(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n264), .A2(G33), .A3(new_n265), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n266), .A2(new_n327), .A3(new_n461), .A4(G116), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n253), .A2(new_n219), .B1(G20), .B2(new_n459), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G283), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n464), .B(new_n255), .C1(G33), .C2(new_n419), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n463), .A2(KEYINPUT20), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT20), .B1(new_n463), .B2(new_n465), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n460), .B(new_n462), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G200), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n458), .B(new_n469), .C1(new_n470), .C2(new_n457), .ZN(new_n471));
  OAI211_X1 g0271(.A(KEYINPUT21), .B(G169), .C1(new_n447), .C2(new_n456), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n446), .A2(new_n291), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n473), .A2(G179), .A3(new_n452), .A4(new_n455), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n468), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n468), .B(G169), .C1(new_n447), .C2(new_n456), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT84), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT21), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n478), .B1(new_n477), .B2(new_n479), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n471), .B(new_n476), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT85), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n477), .A2(new_n479), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT84), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n488), .A2(KEYINPUT85), .A3(new_n476), .A4(new_n471), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n383), .B(G257), .C1(new_n453), .C2(new_n454), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT80), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n448), .A2(new_n451), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n494), .A2(KEYINPUT80), .A3(G257), .A4(new_n383), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(G244), .B(new_n280), .C1(new_n353), .C2(new_n354), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n279), .A2(KEYINPUT4), .A3(G244), .A4(new_n280), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n279), .A2(G250), .A3(G1698), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n499), .A2(new_n500), .A3(new_n464), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n291), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n496), .A2(new_n503), .A3(new_n452), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n319), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n496), .A2(new_n503), .A3(new_n389), .A4(new_n452), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT6), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n507), .A2(new_n419), .A3(G107), .ZN(new_n508));
  XNOR2_X1  g0308(.A(G97), .B(G107), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n508), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  OAI22_X1  g0310(.A1(new_n510), .A2(new_n255), .B1(new_n282), .B2(new_n261), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n335), .B1(new_n367), .B2(new_n369), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n254), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n323), .A2(new_n419), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n266), .A2(new_n327), .A3(new_n461), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G97), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n513), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n505), .A2(new_n506), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT81), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT81), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n505), .A2(new_n521), .A3(new_n506), .A4(new_n518), .ZN(new_n522));
  INV_X1    g0322(.A(new_n518), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n504), .A2(G200), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n523), .B(new_n524), .C1(new_n343), .C2(new_n504), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n520), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n255), .B(G87), .C1(new_n353), .C2(new_n354), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT22), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT22), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n279), .A2(new_n529), .A3(new_n255), .A4(G87), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT24), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT23), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n255), .B2(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n335), .A2(KEYINPUT23), .A3(G20), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n534), .A2(new_n535), .B1(new_n404), .B2(G116), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n531), .A2(new_n532), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n532), .B1(new_n531), .B2(new_n536), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n254), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n266), .A2(G107), .ZN(new_n540));
  XOR2_X1   g0340(.A(KEYINPUT86), .B(KEYINPUT25), .Z(new_n541));
  OR2_X1    g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n541), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n542), .A2(new_n543), .B1(G107), .B2(new_n516), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(G257), .B(G1698), .C1(new_n353), .C2(new_n354), .ZN(new_n546));
  OAI211_X1 g0346(.A(G250), .B(new_n280), .C1(new_n353), .C2(new_n354), .ZN(new_n547));
  INV_X1    g0347(.A(G294), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n546), .B(new_n547), .C1(new_n276), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n291), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n494), .A2(G264), .A3(new_n383), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n550), .A2(new_n452), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G169), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT87), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n550), .A2(G179), .A3(new_n551), .A4(new_n452), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  OR2_X1    g0356(.A1(new_n555), .A2(new_n554), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n545), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(G238), .B(new_n280), .C1(new_n353), .C2(new_n354), .ZN(new_n559));
  OAI211_X1 g0359(.A(G244), .B(G1698), .C1(new_n353), .C2(new_n354), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n559), .B(new_n560), .C1(new_n276), .C2(new_n459), .ZN(new_n561));
  INV_X1    g0361(.A(G250), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n453), .A2(new_n562), .B1(new_n303), .B2(new_n302), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n448), .A2(new_n306), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n291), .A2(new_n561), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n565), .A2(KEYINPUT83), .A3(G190), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n561), .A2(new_n291), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n563), .A2(new_n564), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(G190), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT83), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n565), .A2(new_n470), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n566), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR3_X1   g0373(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n574));
  OR2_X1    g0374(.A1(KEYINPUT82), .A2(KEYINPUT19), .ZN(new_n575));
  NAND2_X1  g0375(.A1(KEYINPUT82), .A2(KEYINPUT19), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n276), .A2(new_n419), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n574), .B1(new_n579), .B2(new_n255), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n279), .A2(new_n255), .A3(G68), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n575), .B(new_n576), .C1(new_n258), .C2(new_n419), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n254), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n323), .A2(new_n330), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n516), .A2(G87), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n573), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n584), .B(new_n585), .C1(new_n330), .C2(new_n515), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n567), .A2(new_n568), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n319), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n565), .A2(new_n389), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n590), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n448), .A2(new_n451), .B1(new_n303), .B2(new_n302), .ZN(new_n595));
  AOI22_X1  g0395(.A1(G264), .A2(new_n595), .B1(new_n549), .B2(new_n291), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n596), .A2(G190), .A3(new_n452), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n552), .A2(G200), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n539), .A2(new_n544), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n558), .A2(new_n589), .A3(new_n594), .A4(new_n599), .ZN(new_n600));
  NOR4_X1   g0400(.A1(new_n442), .A2(new_n490), .A3(new_n526), .A4(new_n600), .ZN(G372));
  AND2_X1   g0401(.A1(new_n401), .A2(new_n399), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT89), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n342), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n341), .B(KEYINPUT89), .C1(G179), .C2(new_n340), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n604), .A2(new_n440), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n437), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n602), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n375), .A2(new_n390), .A3(new_n393), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n393), .B1(new_n375), .B2(new_n390), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n315), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT88), .ZN(new_n614));
  XNOR2_X1  g0414(.A(new_n587), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n573), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n476), .B1(new_n480), .B2(new_n481), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n545), .A2(new_n556), .A3(new_n557), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n599), .B(new_n616), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n594), .B1(new_n619), .B2(new_n526), .ZN(new_n620));
  INV_X1    g0420(.A(new_n519), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT26), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n621), .A2(new_n616), .A3(new_n622), .A4(new_n594), .ZN(new_n623));
  AND4_X1   g0423(.A1(KEYINPUT83), .A2(new_n567), .A3(G190), .A4(new_n568), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n591), .A2(G200), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT83), .B1(new_n565), .B2(G190), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n594), .B1(new_n627), .B2(new_n587), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n520), .B2(new_n522), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n623), .B1(new_n629), .B2(new_n622), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n620), .A2(new_n630), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n613), .B(new_n321), .C1(new_n442), .C2(new_n631), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n632), .B(KEYINPUT90), .ZN(G369));
  INV_X1    g0433(.A(G13), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(G20), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n270), .A2(new_n635), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(G213), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(G343), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(new_n469), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n490), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n617), .A2(new_n643), .ZN(new_n645));
  OAI21_X1  g0445(.A(G330), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n558), .A2(new_n599), .ZN(new_n648));
  INV_X1    g0448(.A(new_n545), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n648), .B1(new_n649), .B2(new_n642), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n618), .A2(new_n641), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n641), .B1(new_n488), .B2(new_n476), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n654), .A2(new_n648), .B1(new_n618), .B2(new_n642), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n653), .A2(new_n655), .ZN(G399));
  NAND2_X1  g0456(.A1(new_n574), .A2(new_n459), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n211), .A2(new_n294), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(G1), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n216), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n660), .B1(new_n661), .B2(new_n659), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT28), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n629), .A2(new_n622), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n616), .A2(new_n594), .ZN(new_n665));
  OAI21_X1  g0465(.A(KEYINPUT26), .B1(new_n665), .B2(new_n519), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n642), .B1(new_n667), .B2(new_n620), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT29), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT29), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n670), .B(new_n642), .C1(new_n620), .C2(new_n630), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n526), .A2(new_n600), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n484), .A2(new_n489), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n674), .A3(new_n642), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT30), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n457), .A2(G179), .A3(new_n565), .A4(new_n596), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n676), .B1(new_n677), .B2(new_n504), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n550), .A2(new_n551), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n474), .A2(new_n591), .A3(new_n679), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n496), .A2(new_n503), .A3(new_n452), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(new_n681), .A3(KEYINPUT30), .ZN(new_n682));
  INV_X1    g0482(.A(new_n456), .ZN(new_n683));
  AOI21_X1  g0483(.A(G179), .B1(new_n683), .B2(new_n473), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n684), .A2(new_n504), .A3(new_n591), .A4(new_n552), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n678), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n686), .A2(KEYINPUT31), .A3(new_n641), .ZN(new_n687));
  AOI21_X1  g0487(.A(KEYINPUT31), .B1(new_n686), .B2(new_n641), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT91), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n686), .A2(new_n641), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT31), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT91), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n686), .A2(KEYINPUT31), .A3(new_n641), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n675), .A2(new_n689), .A3(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n672), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n663), .B1(new_n698), .B2(G1), .ZN(G364));
  NOR2_X1   g0499(.A1(new_n319), .A2(KEYINPUT95), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n255), .B1(KEYINPUT95), .B2(new_n319), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n219), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(G20), .A2(G179), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n705), .B(KEYINPUT96), .Z(new_n706));
  NOR2_X1   g0506(.A1(new_n343), .A2(G200), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n343), .A2(new_n470), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  AOI22_X1  g0512(.A1(G322), .A2(new_n709), .B1(new_n712), .B2(G326), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n707), .A2(new_n389), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G20), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G294), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n255), .A2(G179), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(new_n343), .A3(new_n470), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n279), .B1(new_n719), .B2(G329), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n717), .A2(G190), .A3(G200), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n717), .A2(new_n343), .A3(G200), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n722), .A2(G303), .B1(new_n724), .B2(G283), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n713), .A2(new_n716), .A3(new_n720), .A4(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(G311), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n706), .A2(new_n343), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G200), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n728), .A2(new_n470), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  XOR2_X1   g0532(.A(KEYINPUT33), .B(G317), .Z(new_n733));
  OAI22_X1  g0533(.A1(new_n727), .A2(new_n730), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n726), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT97), .Z(new_n736));
  NAND2_X1  g0536(.A1(new_n715), .A2(G97), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n737), .B(new_n279), .C1(new_n708), .C2(new_n201), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n738), .B1(G50), .B2(new_n712), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n731), .A2(G68), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n729), .A2(G77), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT32), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n742), .B1(new_n719), .B2(G159), .ZN(new_n743));
  INV_X1    g0543(.A(G159), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n718), .A2(KEYINPUT32), .A3(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G87), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n721), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n723), .A2(new_n335), .ZN(new_n748));
  NOR4_X1   g0548(.A1(new_n743), .A2(new_n745), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n739), .A2(new_n740), .A3(new_n741), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n736), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n704), .B1(new_n751), .B2(KEYINPUT98), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(KEYINPUT98), .B2(new_n751), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT94), .Z(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n703), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n355), .A2(new_n357), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n211), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n248), .A2(new_n295), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT93), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n762), .B(new_n764), .C1(new_n295), .C2(new_n217), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n279), .A2(new_n211), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(G355), .B2(KEYINPUT92), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(KEYINPUT92), .B2(G355), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G116), .B2(new_n211), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n759), .B1(new_n765), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n635), .A2(G45), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n771), .A2(G1), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n659), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n753), .A2(new_n770), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n644), .A2(new_n645), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n776), .B1(new_n777), .B2(new_n758), .ZN(new_n778));
  INV_X1    g0578(.A(new_n775), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n646), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G330), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n780), .B1(new_n781), .B2(new_n777), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(G396));
  OAI21_X1  g0584(.A(new_n641), .B1(new_n332), .B2(new_n326), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n604), .A2(new_n605), .A3(new_n786), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n342), .B(new_n785), .C1(new_n346), .C2(new_n348), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(new_n631), .B2(new_n641), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n789), .B(new_n642), .C1(new_n620), .C2(new_n630), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(new_n697), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n697), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n794), .A2(new_n779), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(KEYINPUT99), .B(G143), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G137), .A2(new_n712), .B1(new_n709), .B2(new_n798), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n799), .B1(new_n730), .B2(new_n744), .C1(new_n259), .C2(new_n732), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT34), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n724), .A2(G68), .ZN(new_n802));
  INV_X1    g0602(.A(new_n715), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n802), .B1(new_n215), .B2(new_n721), .C1(new_n803), .C2(new_n201), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n761), .B(new_n804), .C1(G132), .C2(new_n719), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G303), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n548), .A2(new_n708), .B1(new_n711), .B2(new_n807), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n737), .B(new_n368), .C1(new_n727), .C2(new_n718), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n746), .A2(new_n723), .B1(new_n721), .B2(new_n335), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G283), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n811), .B1(new_n459), .B2(new_n730), .C1(new_n812), .C2(new_n732), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n704), .B1(new_n806), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n703), .A2(new_n754), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n779), .B(new_n814), .C1(new_n282), .C2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n755), .B2(new_n789), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n796), .A2(new_n817), .ZN(G384));
  NOR2_X1   g0618(.A1(new_n270), .A2(new_n635), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT37), .ZN(new_n820));
  INV_X1    g0620(.A(new_n639), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n375), .A2(new_n821), .ZN(new_n822));
  AND4_X1   g0622(.A1(new_n820), .A2(new_n391), .A3(new_n822), .A4(new_n397), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n364), .A2(new_n254), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n352), .B1(new_n363), .B2(new_n202), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT102), .ZN(new_n826));
  AOI21_X1  g0626(.A(KEYINPUT16), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI211_X1 g0627(.A(KEYINPUT102), .B(new_n352), .C1(new_n363), .C2(new_n202), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n824), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n374), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n821), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n390), .B1(new_n829), .B2(new_n830), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n831), .A2(new_n832), .A3(new_n397), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n823), .B1(KEYINPUT37), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n831), .B1(new_n602), .B2(new_n611), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT38), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n358), .A2(new_n359), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n360), .A2(new_n362), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n202), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n826), .B1(new_n840), .B2(new_n366), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n841), .A2(new_n365), .A3(new_n828), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n364), .A2(new_n254), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n830), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n390), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n397), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n844), .A2(new_n639), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT37), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n391), .A2(new_n822), .A3(new_n820), .A4(new_n397), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n402), .A2(new_n847), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT38), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT39), .B1(new_n837), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n822), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n402), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n391), .A2(new_n822), .A3(new_n397), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(KEYINPUT37), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n849), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT38), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n850), .A2(KEYINPUT38), .A3(new_n851), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT39), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n853), .A2(KEYINPUT103), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n607), .A2(new_n642), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n836), .B1(new_n834), .B2(new_n835), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n861), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT103), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n868), .A2(new_n869), .A3(KEYINPUT39), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n864), .A2(new_n866), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n611), .A2(new_n821), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n430), .A2(new_n433), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n435), .A2(G169), .A3(new_n432), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n440), .A2(new_n873), .A3(new_n427), .A4(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT101), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n415), .A2(new_n642), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n877), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n437), .A2(new_n440), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n876), .B1(new_n875), .B2(new_n877), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n342), .A2(new_n641), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n883), .B1(new_n792), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n872), .B1(new_n886), .B2(new_n868), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n871), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n613), .A2(new_n321), .ZN(new_n889));
  INV_X1    g0689(.A(new_n442), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n889), .B1(new_n890), .B2(new_n672), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n888), .B(new_n891), .Z(new_n892));
  AOI22_X1  g0692(.A1(new_n848), .A2(new_n849), .B1(new_n402), .B2(new_n847), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n859), .B1(KEYINPUT38), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n687), .A2(new_n688), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n675), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(new_n882), .A3(new_n789), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT40), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT40), .ZN(new_n899));
  INV_X1    g0699(.A(new_n878), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n881), .A2(new_n880), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n900), .A2(new_n901), .A3(new_n789), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n868), .A2(new_n899), .A3(new_n896), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n442), .B1(new_n675), .B2(new_n895), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n904), .A2(new_n905), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n907), .A2(new_n908), .A3(new_n781), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n819), .B1(new_n892), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n892), .B2(new_n910), .ZN(new_n912));
  INV_X1    g0712(.A(new_n510), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n459), .B(new_n221), .C1(new_n913), .C2(KEYINPUT35), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(KEYINPUT35), .B2(new_n913), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT36), .ZN(new_n916));
  OAI21_X1  g0716(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n661), .A2(new_n917), .B1(G50), .B2(new_n202), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(new_n634), .A3(new_n293), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT100), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n912), .A2(new_n921), .ZN(G367));
  OAI21_X1  g0722(.A(new_n759), .B1(new_n211), .B2(new_n330), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n238), .A2(new_n762), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n775), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n259), .A2(new_n708), .B1(new_n711), .B2(new_n797), .ZN(new_n926));
  INV_X1    g0726(.A(G137), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n279), .B1(new_n718), .B2(new_n927), .C1(new_n282), .C2(new_n723), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n803), .A2(new_n202), .B1(new_n721), .B2(new_n201), .ZN(new_n929));
  NOR3_X1   g0729(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  OAI221_X1 g0730(.A(new_n930), .B1(new_n215), .B2(new_n730), .C1(new_n744), .C2(new_n732), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n803), .A2(new_n335), .B1(new_n723), .B2(new_n419), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n760), .B(new_n932), .C1(G317), .C2(new_n719), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n933), .B1(new_n812), .B2(new_n730), .C1(new_n548), .C2(new_n732), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n721), .A2(new_n459), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n709), .A2(G303), .B1(KEYINPUT46), .B2(new_n935), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n936), .B1(KEYINPUT46), .B2(new_n935), .C1(new_n727), .C2(new_n711), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n931), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT47), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n925), .B1(new_n939), .B2(new_n703), .ZN(new_n940));
  OR3_X1    g0740(.A1(new_n615), .A2(new_n594), .A3(new_n642), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n615), .A2(new_n642), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n941), .B1(new_n665), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n940), .B1(new_n943), .B2(new_n757), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT109), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n772), .B(KEYINPUT108), .Z(new_n946));
  OR2_X1    g0746(.A1(new_n672), .A2(new_n697), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n654), .A2(new_n648), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n652), .B2(new_n654), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n647), .A2(KEYINPUT107), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT107), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n646), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n950), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n949), .B1(new_n646), .B2(new_n952), .ZN(new_n955));
  NOR3_X1   g0755(.A1(new_n947), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT105), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n518), .A2(new_n641), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n520), .A2(new_n522), .A3(new_n525), .A4(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n621), .A2(new_n641), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n655), .A2(new_n957), .A3(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT45), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n957), .B1(new_n655), .B2(new_n961), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n964), .B1(new_n963), .B2(new_n965), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n655), .A2(new_n961), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT44), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n653), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT106), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT106), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n970), .A2(new_n971), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n956), .A2(new_n974), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n977), .A2(new_n698), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n659), .B(KEYINPUT41), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n946), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n961), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(new_n948), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT42), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n981), .A2(new_n558), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n520), .A2(new_n522), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n642), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n983), .A2(new_n986), .B1(KEYINPUT43), .B2(new_n943), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n989), .A2(new_n971), .A3(new_n961), .A4(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT104), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n991), .A2(new_n992), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n989), .A2(new_n990), .B1(new_n971), .B2(new_n961), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n945), .B1(new_n980), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(G387));
  XNOR2_X1  g0798(.A(new_n646), .B(new_n952), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n955), .B1(new_n999), .B2(new_n949), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n659), .B1(new_n1000), .B2(new_n698), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n947), .B1(new_n954), .B2(new_n955), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n650), .A2(new_n651), .A3(new_n758), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n658), .A2(new_n766), .B1(G107), .B2(new_n211), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT111), .Z(new_n1005));
  OR2_X1    g0805(.A1(new_n243), .A2(new_n295), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n257), .A2(G50), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT50), .ZN(new_n1008));
  AOI211_X1 g0808(.A(G45), .B(new_n657), .C1(G68), .C2(G77), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n762), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1005), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n759), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n775), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n803), .A2(new_n330), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(G97), .B2(new_n724), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n282), .B2(new_n721), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(new_n328), .B2(new_n731), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n760), .B1(new_n259), .B2(new_n718), .C1(new_n711), .C2(new_n744), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G50), .B2(new_n709), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1017), .B(new_n1019), .C1(new_n202), .C2(new_n730), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n760), .B1(G326), .B2(new_n719), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n803), .A2(new_n812), .B1(new_n721), .B2(new_n548), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G317), .A2(new_n709), .B1(new_n712), .B2(G322), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n730), .B2(new_n807), .C1(new_n727), .C2(new_n732), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT48), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1022), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n1025), .B2(new_n1024), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT49), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1021), .B1(new_n459), .B2(new_n723), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1020), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1013), .B1(new_n1031), .B2(new_n703), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1001), .A2(new_n1002), .B1(new_n1003), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n999), .A2(new_n949), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n955), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n946), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(KEYINPUT110), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT110), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1000), .A2(new_n1039), .A3(new_n1036), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1033), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(KEYINPUT112), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT112), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1033), .A2(new_n1044), .A3(new_n1041), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1045), .ZN(G393));
  NAND3_X1  g0846(.A1(new_n976), .A2(new_n972), .A3(new_n1036), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n759), .B1(new_n419), .B2(new_n211), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n762), .A2(new_n251), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n775), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n259), .A2(new_n711), .B1(new_n708), .B2(new_n744), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT113), .Z(new_n1052));
  OR2_X1    g0852(.A1(new_n1052), .A2(KEYINPUT51), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(KEYINPUT51), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n215), .A2(new_n732), .B1(new_n730), .B2(new_n257), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n760), .B1(new_n718), .B2(new_n797), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n715), .A2(G77), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n202), .B2(new_n721), .C1(new_n746), .C2(new_n723), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n1055), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1053), .A2(new_n1054), .A3(new_n1059), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n279), .B(new_n748), .C1(G322), .C2(new_n719), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n812), .B2(new_n721), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT114), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G311), .A2(new_n709), .B1(new_n712), .B2(G317), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT52), .Z(new_n1065));
  OAI22_X1  g0865(.A1(new_n732), .A2(new_n807), .B1(new_n459), .B2(new_n803), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G294), .B2(new_n729), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1063), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1060), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1050), .B1(new_n1069), .B2(new_n703), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n961), .B2(new_n757), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1047), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n976), .A2(new_n972), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1000), .A2(new_n698), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n659), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1076), .A2(new_n977), .A3(KEYINPUT115), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(KEYINPUT115), .B1(new_n1076), .B2(new_n977), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1073), .B1(new_n1078), .B2(new_n1079), .ZN(G390));
  AOI21_X1  g0880(.A(new_n781), .B1(new_n675), .B2(new_n895), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n883), .B1(new_n1082), .B2(new_n790), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n885), .B1(new_n668), .B2(new_n790), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n696), .A2(G330), .A3(new_n789), .A4(new_n882), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1083), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT116), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n696), .A2(G330), .A3(new_n789), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n883), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n902), .A2(new_n1081), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n792), .A2(new_n885), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1088), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1089), .A2(new_n883), .B1(new_n902), .B2(new_n1081), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1093), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n1095), .A2(KEYINPUT116), .A3(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1087), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n890), .A2(new_n1081), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n891), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1091), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n866), .B1(new_n1093), .B2(new_n882), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n864), .B2(new_n870), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n866), .B(new_n894), .C1(new_n882), .C2(new_n1084), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1103), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n894), .A2(new_n866), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n1085), .B2(new_n883), .ZN(new_n1109));
  AOI211_X1 g0909(.A(KEYINPUT103), .B(new_n862), .C1(new_n867), .C2(new_n861), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n869), .B1(new_n868), .B2(KEYINPUT39), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1110), .B1(new_n1111), .B2(new_n863), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1109), .B(new_n1086), .C1(new_n1112), .C2(new_n1104), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1107), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1102), .A2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1098), .A2(new_n1107), .A3(new_n1113), .A4(new_n1101), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1115), .A2(new_n774), .A3(new_n1116), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1107), .A2(new_n1113), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n1112), .A2(new_n755), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n815), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n775), .B1(new_n1120), .B2(new_n328), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n721), .A2(new_n259), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT53), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT54), .B(G143), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n1123), .B1(new_n730), .B2(new_n1124), .C1(new_n927), .C2(new_n732), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G128), .A2(new_n712), .B1(new_n709), .B2(G132), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n723), .A2(new_n215), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n368), .B(new_n1127), .C1(G125), .C2(new_n719), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1126), .B(new_n1128), .C1(new_n744), .C2(new_n803), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(G116), .A2(new_n709), .B1(new_n712), .B2(G283), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n279), .B(new_n747), .C1(G294), .C2(new_n719), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1130), .A2(new_n1131), .A3(new_n802), .A4(new_n1057), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n419), .A2(new_n730), .B1(new_n732), .B2(new_n335), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n1125), .A2(new_n1129), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1121), .B1(new_n1134), .B2(new_n703), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1118), .A2(new_n1036), .B1(new_n1119), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1117), .A2(new_n1136), .ZN(G378));
  OAI21_X1  g0937(.A(new_n775), .B1(new_n1120), .B2(G50), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n761), .B(new_n294), .C1(new_n711), .C2(new_n459), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n724), .A2(G58), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n282), .B2(new_n721), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n803), .A2(new_n202), .B1(new_n812), .B2(new_n718), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(G97), .C2(new_n731), .ZN(new_n1143));
  OR2_X1    g0943(.A1(new_n730), .A2(new_n330), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1139), .B(new_n1145), .C1(G107), .C2(new_n709), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(G50), .B1(new_n276), .B2(new_n294), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n760), .B2(G41), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n709), .A2(G128), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1153), .B1(new_n259), .B2(new_n803), .C1(new_n721), .C2(new_n1124), .ZN(new_n1154));
  INV_X1    g0954(.A(G132), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n1155), .A2(new_n732), .B1(new_n730), .B2(new_n927), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1154), .B(new_n1156), .C1(G125), .C2(new_n712), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n724), .A2(G159), .ZN(new_n1161));
  AOI211_X1 g0961(.A(G33), .B(G41), .C1(new_n719), .C2(G124), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1152), .B1(new_n1159), .B2(new_n1163), .C1(new_n1148), .C2(new_n1147), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1138), .B1(new_n1164), .B2(new_n703), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n318), .A2(new_n821), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n315), .A2(new_n321), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1168), .B1(new_n315), .B2(new_n321), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1167), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1168), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n322), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1174), .A2(new_n1169), .A3(new_n1166), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n754), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1165), .A2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT118), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1179), .A2(KEYINPUT119), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(KEYINPUT119), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n902), .B(new_n896), .C1(new_n837), .C2(new_n859), .ZN(new_n1182));
  AND4_X1   g0982(.A1(new_n899), .A2(new_n896), .A3(new_n789), .A4(new_n882), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(KEYINPUT40), .A2(new_n1182), .B1(new_n1183), .B2(new_n868), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1176), .B1(new_n1184), .B2(new_n781), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1176), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n904), .A2(G330), .A3(new_n1186), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1185), .A2(new_n871), .A3(new_n887), .A4(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1186), .B1(new_n904), .B2(G330), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n781), .B(new_n1176), .C1(new_n898), .C2(new_n903), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n888), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1188), .A2(new_n1191), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1180), .A2(new_n1181), .B1(new_n1036), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1100), .A2(KEYINPUT120), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT120), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n891), .A2(new_n1195), .A3(new_n1099), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1116), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT57), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n1188), .B2(new_n1191), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n1199), .A2(KEYINPUT121), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT121), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1116), .A2(new_n1198), .B1(new_n1188), .B2(new_n1191), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n774), .B1(new_n1205), .B2(KEYINPUT57), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1193), .B1(new_n1204), .B2(new_n1206), .ZN(G375));
  XOR2_X1   g1007(.A(new_n946), .B(KEYINPUT122), .Z(new_n1208));
  NAND3_X1  g1008(.A1(new_n1092), .A2(new_n1088), .A3(new_n1093), .ZN(new_n1209));
  OAI21_X1  g1009(.A(KEYINPUT116), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1208), .B1(new_n1211), .B2(new_n1087), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n882), .A2(new_n755), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n368), .B1(new_n718), .B2(new_n807), .C1(new_n282), .C2(new_n723), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1014), .B(new_n1214), .C1(G97), .C2(new_n722), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G283), .A2(new_n709), .B1(new_n712), .B2(G294), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G107), .A2(new_n729), .B1(new_n731), .B2(G116), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT123), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n761), .B1(G128), .B2(new_n719), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n1155), .B2(new_n711), .C1(new_n927), .C2(new_n708), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1140), .B1(new_n744), .B2(new_n721), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G50), .B2(new_n715), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1223), .B1(new_n259), .B2(new_n730), .C1(new_n732), .C2(new_n1124), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1219), .B1(new_n1221), .B2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1218), .A2(KEYINPUT123), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n703), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1227), .B(new_n775), .C1(G68), .C2(new_n1120), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1213), .A2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(KEYINPUT124), .B1(new_n1212), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT124), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1229), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1083), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1231), .B(new_n1232), .C1(new_n1234), .C2(new_n1208), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1230), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n979), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1100), .B(new_n1087), .C1(new_n1094), .C2(new_n1097), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1102), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1236), .A2(new_n1239), .ZN(G381));
  NAND2_X1  g1040(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1192), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1241), .B1(new_n946), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT121), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1234), .A2(new_n1100), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1197), .B1(new_n1118), .B2(new_n1245), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n888), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1185), .A2(new_n1187), .B1(new_n871), .B2(new_n887), .ZN(new_n1248));
  OAI21_X1  g1048(.A(KEYINPUT57), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1244), .B1(new_n1246), .B2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1199), .A2(KEYINPUT121), .A3(new_n1201), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1199), .A2(new_n1192), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n659), .B1(new_n1253), .B2(new_n1200), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1243), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(G378), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1043), .A2(new_n783), .A3(new_n1045), .ZN(new_n1258));
  OR3_X1    g1058(.A1(new_n1258), .A2(G390), .A3(G384), .ZN(new_n1259));
  OR4_X1    g1059(.A1(G387), .A2(new_n1257), .A3(G381), .A4(new_n1259), .ZN(G407));
  OAI211_X1 g1060(.A(G407), .B(G213), .C1(G343), .C2(new_n1257), .ZN(G409));
  AND3_X1   g1061(.A1(new_n1033), .A2(new_n1044), .A3(new_n1041), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1044), .B1(new_n1033), .B2(new_n1041), .ZN(new_n1263));
  OAI21_X1  g1063(.A(G396), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1264), .A2(new_n1258), .A3(G390), .ZN(new_n1265));
  AOI21_X1  g1065(.A(G390), .B1(new_n1264), .B2(new_n1258), .ZN(new_n1266));
  OAI21_X1  g1066(.A(G387), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1264), .A2(new_n1258), .ZN(new_n1268));
  INV_X1    g1068(.A(G390), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1264), .A2(new_n1258), .A3(G390), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1270), .A2(new_n997), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1267), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n640), .A2(G213), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1117), .A2(new_n1136), .A3(new_n1179), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n979), .B1(new_n1116), .B2(new_n1198), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1208), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1192), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1275), .B1(new_n1277), .B2(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT126), .ZN(new_n1283));
  INV_X1    g1083(.A(G384), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(KEYINPUT125), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n796), .A2(KEYINPUT125), .A3(new_n817), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n659), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1234), .A2(KEYINPUT60), .A3(new_n1100), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT60), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1238), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1287), .A2(new_n1288), .A3(new_n1290), .ZN(new_n1291));
  AOI211_X1 g1091(.A(new_n1285), .B(new_n1286), .C1(new_n1236), .C2(new_n1291), .ZN(new_n1292));
  AND4_X1   g1092(.A1(KEYINPUT125), .A2(new_n1236), .A3(new_n1284), .A4(new_n1291), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1283), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1098), .A2(new_n1279), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1231), .B1(new_n1295), .B2(new_n1232), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1235), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1291), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1285), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1286), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1236), .A2(KEYINPUT125), .A3(new_n1284), .A4(new_n1291), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1301), .A2(KEYINPUT126), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1294), .A2(new_n1303), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1282), .A2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1273), .B1(new_n1305), .B2(KEYINPUT63), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT61), .ZN(new_n1307));
  INV_X1    g1107(.A(G2897), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1274), .B1(KEYINPUT127), .B2(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1309), .B1(KEYINPUT127), .B2(new_n1308), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1294), .A2(new_n1303), .A3(new_n1310), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1312), .A2(G2897), .A3(new_n1275), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1311), .A2(new_n1282), .A3(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT63), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1282), .B2(new_n1304), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1306), .A2(new_n1307), .A3(new_n1314), .A4(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(KEYINPUT62), .B1(new_n1282), .B2(new_n1304), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1280), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1274), .B1(new_n1319), .B2(new_n1276), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1320), .B1(G375), .B2(G378), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1301), .A2(KEYINPUT126), .A3(new_n1302), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT126), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT62), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1321), .A2(new_n1324), .A3(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1318), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1314), .A2(new_n1307), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1273), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1317), .A2(new_n1329), .ZN(G405));
  NAND2_X1  g1130(.A1(G375), .A2(G378), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1304), .A2(new_n1331), .A3(new_n1257), .ZN(new_n1332));
  AND2_X1   g1132(.A1(new_n1331), .A2(new_n1257), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1332), .B1(new_n1333), .B2(new_n1312), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1334), .A2(new_n1272), .A3(new_n1267), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1332), .B(new_n1273), .C1(new_n1333), .C2(new_n1312), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(G402));
endmodule


