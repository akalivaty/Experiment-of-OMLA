//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n816, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT71), .ZN(new_n203));
  XOR2_X1   g002(.A(G71gat), .B(G99gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G127gat), .B(G134gat), .ZN(new_n206));
  OR2_X1    g005(.A1(new_n206), .A2(KEYINPUT69), .ZN(new_n207));
  INV_X1    g006(.A(G113gat), .ZN(new_n208));
  INV_X1    g007(.A(G120gat), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT1), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G113gat), .A2(G120gat), .ZN(new_n211));
  AOI22_X1  g010(.A1(new_n206), .A2(KEYINPUT69), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n207), .B(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT27), .B(G183gat), .ZN(new_n215));
  INV_X1    g014(.A(G190gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT28), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT28), .B1(new_n215), .B2(new_n216), .ZN(new_n220));
  INV_X1    g019(.A(G169gat), .ZN(new_n221));
  INV_X1    g020(.A(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT26), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(KEYINPUT67), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n221), .A2(new_n222), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(new_n223), .B2(KEYINPUT26), .ZN(new_n228));
  OAI221_X1 g027(.A(new_n214), .B1(new_n219), .B2(new_n220), .C1(new_n225), .C2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT68), .ZN(new_n230));
  NOR2_X1   g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n231), .A2(KEYINPUT65), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n214), .A2(KEYINPUT24), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT24), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(G183gat), .A3(G190gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n231), .A2(KEYINPUT65), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT23), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n223), .B1(new_n226), .B2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT23), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n238), .A2(KEYINPUT25), .A3(new_n240), .A4(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT66), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n241), .B(KEYINPUT64), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n236), .B1(G183gat), .B2(G190gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(new_n240), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT25), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n213), .B1(new_n230), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G227gat), .ZN(new_n251));
  INV_X1    g050(.A(G233gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n229), .B(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n213), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n243), .A2(new_n248), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n250), .A2(new_n253), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT33), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n205), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n261), .A2(KEYINPUT70), .B1(KEYINPUT32), .B2(new_n259), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n205), .A2(new_n260), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n259), .A2(KEYINPUT32), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT34), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n250), .A2(new_n258), .ZN(new_n271));
  INV_X1    g070(.A(new_n253), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI211_X1 g072(.A(KEYINPUT34), .B(new_n253), .C1(new_n250), .C2(new_n258), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n263), .A2(new_n269), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n267), .B1(new_n261), .B2(new_n264), .ZN(new_n277));
  OAI22_X1  g076(.A1(new_n262), .A2(new_n277), .B1(new_n273), .B2(new_n274), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT31), .B(G50gat), .ZN(new_n280));
  INV_X1    g079(.A(G106gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G228gat), .A2(G233gat), .ZN(new_n284));
  XOR2_X1   g083(.A(new_n284), .B(KEYINPUT78), .Z(new_n285));
  XOR2_X1   g084(.A(KEYINPUT76), .B(G141gat), .Z(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G148gat), .ZN(new_n287));
  INV_X1    g086(.A(G148gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G141gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(G155gat), .A2(G162gat), .ZN(new_n290));
  OR3_X1    g089(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n287), .A2(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OR2_X1    g091(.A1(new_n288), .A2(G141gat), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT2), .B1(new_n293), .B2(new_n289), .ZN(new_n294));
  INV_X1    g093(.A(G155gat), .ZN(new_n295));
  INV_X1    g094(.A(G162gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(new_n296), .A3(KEYINPUT75), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT75), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(G155gat), .B2(G162gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n299), .A3(new_n290), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G197gat), .B(G204gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT22), .ZN(new_n304));
  INV_X1    g103(.A(G211gat), .ZN(new_n305));
  INV_X1    g104(.A(G218gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  XOR2_X1   g107(.A(G211gat), .B(G218gat), .Z(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(KEYINPUT73), .B(KEYINPUT29), .Z(new_n311));
  AOI21_X1  g110(.A(KEYINPUT79), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(KEYINPUT3), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n310), .A2(KEYINPUT79), .A3(new_n311), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n302), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OR3_X1    g114(.A1(new_n292), .A2(KEYINPUT3), .A3(new_n301), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n310), .B1(new_n316), .B2(new_n311), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n285), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT29), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT3), .B1(new_n310), .B2(new_n319), .ZN(new_n320));
  OAI211_X1 g119(.A(G228gat), .B(G233gat), .C1(new_n320), .C2(new_n302), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G22gat), .ZN(new_n325));
  INV_X1    g124(.A(G78gat), .ZN(new_n326));
  INV_X1    g125(.A(G22gat), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n318), .B(new_n327), .C1(new_n317), .C2(new_n321), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n325), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n326), .B1(new_n325), .B2(new_n328), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n283), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n325), .A2(new_n328), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G78gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n325), .A2(new_n326), .A3(new_n328), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n334), .A3(new_n282), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G8gat), .B(G36gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(G64gat), .B(G92gat), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n337), .B(new_n338), .Z(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n310), .ZN(new_n341));
  NAND2_X1  g140(.A1(G226gat), .A2(G233gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n230), .B2(new_n249), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT29), .B1(new_n257), .B2(new_n229), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n344), .B(KEYINPUT74), .C1(new_n343), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n255), .A2(new_n257), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n348), .A3(new_n343), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n341), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n311), .A2(new_n342), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n257), .A2(new_n229), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n343), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n352), .A2(new_n341), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n340), .B1(new_n350), .B2(new_n356), .ZN(new_n357));
  AOI211_X1 g156(.A(KEYINPUT74), .B(new_n342), .C1(new_n255), .C2(new_n257), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n348), .B1(new_n347), .B2(new_n343), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n342), .B1(new_n353), .B2(KEYINPUT29), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n339), .B(new_n355), .C1(new_n361), .C2(new_n341), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n357), .A2(KEYINPUT30), .A3(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n350), .A2(new_n356), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT30), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n365), .A3(new_n339), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n292), .A2(new_n301), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT3), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(new_n316), .A3(new_n256), .ZN(new_n370));
  NAND2_X1  g169(.A1(G225gat), .A2(G233gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n213), .A2(new_n302), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n213), .A2(new_n302), .A3(KEYINPUT4), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n370), .A2(new_n371), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n256), .A2(new_n368), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n371), .B1(new_n377), .B2(new_n372), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT5), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G1gat), .B(G29gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT0), .ZN(new_n382));
  XNOR2_X1  g181(.A(G57gat), .B(G85gat), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n382), .B(new_n383), .Z(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n374), .A2(new_n375), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n386), .A2(KEYINPUT5), .A3(new_n371), .A4(new_n370), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n380), .A2(KEYINPUT6), .A3(new_n385), .A4(new_n387), .ZN(new_n388));
  OR2_X1    g187(.A1(new_n388), .A2(KEYINPUT77), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(KEYINPUT77), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n380), .A2(new_n385), .A3(new_n387), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT6), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n380), .A2(new_n387), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n384), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n389), .A2(new_n390), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n279), .A2(new_n336), .A3(new_n367), .A4(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT35), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n331), .A2(new_n335), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n400), .B1(new_n276), .B2(new_n278), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT35), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n401), .A2(new_n402), .A3(new_n397), .A4(new_n367), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n370), .ZN(new_n405));
  INV_X1    g204(.A(new_n371), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n377), .A2(new_n371), .A3(new_n372), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(KEYINPUT39), .A3(new_n408), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n409), .B(new_n384), .C1(KEYINPUT39), .C2(new_n407), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT40), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n412), .A2(new_n391), .ZN(new_n413));
  OR2_X1    g212(.A1(new_n410), .A2(new_n411), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n413), .A2(new_n363), .A3(new_n366), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n336), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n355), .B1(new_n361), .B2(new_n341), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n340), .B1(new_n417), .B2(KEYINPUT37), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT38), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n310), .B1(new_n346), .B2(new_n349), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n352), .A2(new_n310), .A3(new_n354), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT37), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n419), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n396), .B(new_n362), .C1(new_n418), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n340), .A2(KEYINPUT37), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n357), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT37), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n426), .B1(new_n427), .B2(new_n364), .ZN(new_n428));
  AOI22_X1  g227(.A1(new_n424), .A2(KEYINPUT80), .B1(new_n428), .B2(KEYINPUT38), .ZN(new_n429));
  INV_X1    g228(.A(new_n423), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT80), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n431), .A2(new_n432), .A3(new_n396), .A4(new_n362), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n416), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n363), .A2(new_n366), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n400), .B1(new_n435), .B2(new_n396), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT36), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n437), .B1(new_n279), .B2(KEYINPUT72), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT72), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n276), .A2(new_n278), .A3(new_n439), .A4(KEYINPUT36), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n436), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n404), .B1(new_n434), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(G71gat), .A2(G78gat), .ZN(new_n443));
  NOR2_X1   g242(.A1(G71gat), .A2(G78gat), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT9), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(KEYINPUT90), .A2(G57gat), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(G64gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT91), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT91), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(G64gat), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n449), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n449), .B1(new_n451), .B2(new_n453), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n447), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AND2_X1   g255(.A1(G57gat), .A2(G64gat), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n445), .B(new_n443), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(KEYINPUT92), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT21), .ZN(new_n462));
  INV_X1    g261(.A(G8gat), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT87), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT86), .B(G1gat), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT16), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(G1gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT86), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT86), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(G1gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n472), .A2(KEYINPUT87), .A3(KEYINPUT16), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n467), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(G15gat), .B(G22gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n468), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n463), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n475), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n480), .B1(new_n467), .B2(new_n473), .ZN(new_n481));
  NOR3_X1   g280(.A1(new_n481), .A2(G8gat), .A3(new_n477), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n462), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT93), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n483), .A2(KEYINPUT93), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(new_n295), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n487), .B(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT21), .B1(new_n456), .B2(new_n459), .ZN(new_n491));
  NAND2_X1  g290(.A1(G231gat), .A2(G233gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(G127gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G183gat), .B(G211gat), .ZN(new_n496));
  XOR2_X1   g295(.A(new_n495), .B(new_n496), .Z(new_n497));
  XNOR2_X1  g296(.A(new_n490), .B(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G43gat), .B(G50gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT15), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT84), .ZN(new_n501));
  INV_X1    g300(.A(G29gat), .ZN(new_n502));
  INV_X1    g301(.A(G36gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT14), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT14), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(G29gat), .B2(G36gat), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n501), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n502), .A2(new_n503), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n504), .A2(new_n506), .A3(new_n501), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n500), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n504), .A2(new_n506), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n512), .A2(new_n508), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT85), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT15), .B1(new_n499), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT15), .ZN(new_n516));
  INV_X1    g315(.A(G43gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(G50gat), .ZN(new_n518));
  INV_X1    g317(.A(G50gat), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(G43gat), .ZN(new_n520));
  OAI211_X1 g319(.A(KEYINPUT85), .B(new_n516), .C1(new_n518), .C2(new_n520), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n513), .A2(new_n515), .A3(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n511), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G99gat), .B(G106gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(KEYINPUT96), .A2(G85gat), .A3(G92gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT7), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G99gat), .A2(G106gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT8), .ZN(new_n533));
  NAND2_X1  g332(.A1(G85gat), .A2(G92gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT95), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OR2_X1    g335(.A1(G85gat), .A2(G92gat), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n533), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n525), .B1(new_n531), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n526), .A2(new_n527), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(new_n526), .B2(new_n529), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n533), .A2(new_n536), .A3(new_n537), .ZN(new_n542));
  XOR2_X1   g341(.A(G99gat), .B(G106gat), .Z(new_n543));
  NOR3_X1   g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G232gat), .A2(G233gat), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n524), .A2(new_n545), .B1(KEYINPUT41), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT17), .B1(new_n511), .B2(new_n522), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT17), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n513), .A2(new_n515), .A3(new_n521), .ZN(new_n551));
  INV_X1    g350(.A(new_n510), .ZN(new_n552));
  NOR3_X1   g351(.A1(new_n552), .A2(new_n508), .A3(new_n507), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n550), .B(new_n551), .C1(new_n553), .C2(new_n500), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n545), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT97), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT97), .ZN(new_n558));
  AOI211_X1 g357(.A(new_n558), .B(new_n545), .C1(new_n549), .C2(new_n554), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n548), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G190gat), .B(G218gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT99), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n561), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n565), .B(new_n548), .C1(new_n557), .C2(new_n559), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n547), .A2(KEYINPUT41), .ZN(new_n567));
  XNOR2_X1  g366(.A(G134gat), .B(G162gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n560), .A2(KEYINPUT99), .A3(new_n561), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n564), .A2(new_n566), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n569), .B(KEYINPUT94), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n572), .B1(new_n562), .B2(new_n566), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n573), .A2(KEYINPUT98), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT98), .ZN(new_n575));
  AOI211_X1 g374(.A(new_n575), .B(new_n572), .C1(new_n562), .C2(new_n566), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n571), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G230gat), .A2(G233gat), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n443), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n580), .B1(KEYINPUT9), .B2(new_n444), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n451), .A2(new_n453), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n448), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n449), .A2(new_n451), .A3(new_n453), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n459), .ZN(new_n586));
  OAI22_X1  g385(.A1(new_n539), .A2(new_n544), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT10), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n531), .A2(new_n525), .A3(new_n538), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n543), .B1(new_n541), .B2(new_n542), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n589), .A2(new_n456), .A3(new_n590), .A4(new_n459), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n587), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT100), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT100), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n587), .A2(new_n594), .A3(new_n591), .A4(new_n588), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n556), .A2(new_n588), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n461), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n579), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n587), .A2(new_n591), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n599), .B1(new_n579), .B2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G120gat), .B(G148gat), .Z(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT101), .ZN(new_n603));
  XNOR2_X1  g402(.A(G176gat), .B(G204gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n600), .A2(new_n579), .ZN(new_n607));
  AOI22_X1  g406(.A1(new_n593), .A2(new_n595), .B1(new_n461), .B2(new_n597), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n607), .B(new_n605), .C1(new_n608), .C2(new_n579), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(KEYINPUT81), .B(KEYINPUT11), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT82), .ZN(new_n612));
  XOR2_X1   g411(.A(G113gat), .B(G141gat), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G169gat), .B(G197gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(KEYINPUT88), .B1(new_n479), .B2(new_n482), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n476), .A2(new_n463), .A3(new_n478), .ZN(new_n620));
  OAI21_X1  g419(.A(G8gat), .B1(new_n481), .B2(new_n477), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT88), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n619), .A2(new_n555), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G229gat), .A2(G233gat), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n524), .A2(new_n621), .A3(new_n620), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT18), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n523), .B1(new_n479), .B2(new_n482), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n625), .B(KEYINPUT13), .Z(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n624), .A2(KEYINPUT18), .A3(new_n625), .A4(new_n626), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT89), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n635), .A2(KEYINPUT89), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT83), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n618), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n636), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n635), .A2(KEYINPUT89), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI211_X1 g442(.A(KEYINPUT83), .B(new_n617), .C1(new_n643), .C2(new_n634), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NOR4_X1   g444(.A1(new_n498), .A2(new_n577), .A3(new_n610), .A4(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n442), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(new_n397), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(new_n468), .ZN(G1324gat));
  NOR2_X1   g448(.A1(new_n647), .A2(new_n367), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT16), .B(G8gat), .Z(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(KEYINPUT42), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT103), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n650), .A2(new_n463), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT102), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n650), .A2(new_n651), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n653), .B(new_n655), .C1(KEYINPUT42), .C2(new_n656), .ZN(G1325gat));
  NAND2_X1  g456(.A1(new_n438), .A2(new_n440), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(G15gat), .B1(new_n647), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(G15gat), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n279), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n660), .B1(new_n647), .B2(new_n662), .ZN(G1326gat));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n336), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT43), .B(G22gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1327gat));
  INV_X1    g465(.A(new_n577), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n436), .A2(new_n438), .A3(new_n440), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n423), .B1(new_n357), .B2(new_n425), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n389), .A2(new_n390), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n393), .A2(new_n395), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n670), .A2(new_n671), .A3(new_n362), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT80), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n428), .A2(KEYINPUT38), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n433), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n675), .A2(new_n336), .A3(new_n415), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n668), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n667), .B1(new_n677), .B2(new_n404), .ZN(new_n678));
  INV_X1    g477(.A(new_n498), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n679), .A2(new_n610), .A3(new_n645), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n681), .A2(new_n502), .A3(new_n396), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT45), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n442), .A2(new_n577), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n442), .A2(KEYINPUT44), .A3(new_n577), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n680), .B(KEYINPUT104), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(G29gat), .B1(new_n690), .B2(new_n397), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n683), .A2(new_n691), .ZN(G1328gat));
  AOI21_X1  g491(.A(G36gat), .B1(KEYINPUT105), .B2(KEYINPUT46), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n681), .A2(new_n435), .A3(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(G36gat), .B1(new_n690), .B2(new_n367), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(G1329gat));
  NAND4_X1  g497(.A1(new_n686), .A2(new_n658), .A3(new_n687), .A4(new_n689), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(G43gat), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n681), .A2(new_n517), .A3(new_n279), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1330gat));
  NAND4_X1  g503(.A1(new_n686), .A2(new_n400), .A3(new_n687), .A4(new_n689), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(G50gat), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n681), .A2(new_n519), .A3(new_n400), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT48), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1331gat));
  INV_X1    g509(.A(new_n645), .ZN(new_n711));
  INV_X1    g510(.A(new_n610), .ZN(new_n712));
  NOR4_X1   g511(.A1(new_n498), .A2(new_n711), .A3(new_n577), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT106), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n442), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n396), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(G57gat), .ZN(G1332gat));
  INV_X1    g516(.A(KEYINPUT49), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n435), .B1(new_n718), .B2(new_n450), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT107), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n718), .A2(new_n450), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1333gat));
  NAND2_X1  g522(.A1(new_n715), .A2(new_n658), .ZN(new_n724));
  AOI21_X1  g523(.A(G71gat), .B1(new_n276), .B2(new_n278), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n724), .A2(G71gat), .B1(new_n715), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g526(.A1(new_n715), .A2(new_n400), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g528(.A1(new_n679), .A2(new_n711), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n610), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n688), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733), .B2(new_n397), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n678), .A2(KEYINPUT108), .A3(KEYINPUT51), .A4(new_n730), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n442), .A2(KEYINPUT51), .A3(new_n577), .A4(new_n730), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT51), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n442), .A2(new_n577), .A3(new_n730), .ZN(new_n740));
  AOI22_X1  g539(.A1(new_n735), .A2(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OR3_X1    g540(.A1(new_n397), .A2(G85gat), .A3(new_n712), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n734), .B1(new_n741), .B2(new_n742), .ZN(G1336gat));
  OR3_X1    g542(.A1(new_n367), .A2(G92gat), .A3(new_n712), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n735), .A2(new_n738), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n442), .A2(KEYINPUT109), .A3(new_n577), .A4(new_n730), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n747), .A2(new_n739), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n744), .B1(new_n745), .B2(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n686), .A2(new_n435), .A3(new_n687), .A4(new_n732), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n751), .A2(G92gat), .ZN(new_n752));
  OAI21_X1  g551(.A(KEYINPUT52), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT52), .B1(new_n751), .B2(G92gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n740), .A2(new_n739), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n744), .B1(new_n745), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n756), .B2(KEYINPUT110), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n741), .A2(new_n758), .A3(new_n744), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n753), .B1(new_n757), .B2(new_n759), .ZN(G1337gat));
  OAI21_X1  g559(.A(G99gat), .B1(new_n733), .B2(new_n659), .ZN(new_n761));
  INV_X1    g560(.A(G99gat), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n279), .A2(new_n762), .A3(new_n610), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n741), .B2(new_n763), .ZN(G1338gat));
  NAND3_X1  g563(.A1(new_n400), .A2(new_n281), .A3(new_n610), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(new_n745), .B2(new_n749), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n686), .A2(new_n400), .A3(new_n687), .A4(new_n732), .ZN(new_n767));
  XNOR2_X1  g566(.A(KEYINPUT111), .B(G106gat), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT53), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT53), .B1(new_n767), .B2(new_n768), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n741), .B2(new_n765), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(G1339gat));
  NOR4_X1   g572(.A1(new_n498), .A2(new_n711), .A3(new_n577), .A4(new_n610), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n596), .A2(new_n579), .A3(new_n598), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n596), .A2(new_n598), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n578), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n608), .A2(KEYINPUT112), .A3(new_n579), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n777), .A2(new_n779), .A3(KEYINPUT54), .A4(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n605), .B1(new_n599), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT55), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785));
  AOI211_X1 g584(.A(new_n785), .B(new_n605), .C1(new_n599), .C2(new_n782), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n781), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n609), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT113), .ZN(new_n789));
  INV_X1    g588(.A(new_n609), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n786), .B2(new_n781), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n784), .B1(new_n789), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n638), .A2(new_n617), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n625), .B1(new_n624), .B2(new_n626), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n631), .A2(new_n632), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n616), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n794), .A2(new_n577), .A3(new_n800), .ZN(new_n801));
  AOI22_X1  g600(.A1(new_n794), .A2(new_n711), .B1(new_n610), .B2(new_n800), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n802), .B2(new_n577), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n774), .B1(new_n803), .B2(new_n498), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n400), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n435), .A2(new_n397), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(new_n279), .A3(new_n806), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n807), .A2(new_n208), .A3(new_n645), .ZN(new_n808));
  INV_X1    g607(.A(new_n401), .ZN(new_n809));
  NOR4_X1   g608(.A1(new_n804), .A2(new_n397), .A3(new_n435), .A4(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(G113gat), .B1(new_n810), .B2(new_n711), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n808), .A2(new_n811), .ZN(G1340gat));
  NOR3_X1   g611(.A1(new_n807), .A2(new_n209), .A3(new_n712), .ZN(new_n813));
  AOI21_X1  g612(.A(G120gat), .B1(new_n810), .B2(new_n610), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(G1341gat));
  OAI21_X1  g614(.A(G127gat), .B1(new_n807), .B2(new_n498), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n810), .A2(new_n494), .A3(new_n679), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XOR2_X1   g617(.A(new_n818), .B(KEYINPUT114), .Z(G1342gat));
  OAI21_X1  g618(.A(G134gat), .B1(new_n807), .B2(new_n667), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT115), .ZN(new_n821));
  INV_X1    g620(.A(G134gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n810), .A2(new_n822), .A3(new_n577), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n823), .B(KEYINPUT56), .Z(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n824), .ZN(G1343gat));
  NAND2_X1  g624(.A1(new_n659), .A2(new_n806), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n827), .B1(new_n804), .B2(new_n336), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n336), .A2(new_n827), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n679), .A2(new_n667), .A3(new_n712), .A4(new_n645), .ZN(new_n830));
  INV_X1    g629(.A(new_n784), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n792), .B1(new_n787), .B2(new_n609), .ZN(new_n832));
  AOI211_X1 g631(.A(KEYINPUT113), .B(new_n790), .C1(new_n786), .C2(new_n781), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n577), .B(new_n831), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n799), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n640), .A2(new_n644), .A3(new_n831), .A4(new_n791), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n610), .A2(new_n795), .A3(new_n798), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n577), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n498), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n830), .B1(new_n839), .B2(KEYINPUT116), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n836), .A2(new_n837), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n667), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n679), .B1(new_n842), .B2(new_n801), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n829), .B1(new_n840), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n826), .B1(new_n828), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n286), .B1(new_n847), .B2(new_n711), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n804), .A2(new_n397), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n658), .A2(new_n336), .A3(new_n435), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n645), .A2(G141gat), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT58), .B1(new_n848), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n857), .B1(new_n851), .B2(new_n853), .ZN(new_n858));
  INV_X1    g657(.A(new_n826), .ZN(new_n859));
  INV_X1    g658(.A(new_n829), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n774), .B1(new_n843), .B2(new_n844), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n839), .A2(KEYINPUT116), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n837), .B1(new_n864), .B2(new_n645), .ZN(new_n865));
  INV_X1    g664(.A(new_n834), .ZN(new_n866));
  AOI22_X1  g665(.A1(new_n865), .A2(new_n667), .B1(new_n866), .B2(new_n800), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n830), .B1(new_n867), .B2(new_n679), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT57), .B1(new_n868), .B2(new_n400), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n711), .B(new_n859), .C1(new_n863), .C2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n286), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n828), .A2(new_n846), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n873), .A2(KEYINPUT117), .A3(new_n711), .A4(new_n859), .ZN(new_n874));
  AOI211_X1 g673(.A(new_n856), .B(new_n858), .C1(new_n872), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n870), .A2(new_n871), .ZN(new_n876));
  INV_X1    g675(.A(new_n286), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n877), .A3(new_n874), .ZN(new_n878));
  INV_X1    g677(.A(new_n858), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT118), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n855), .B1(new_n875), .B2(new_n880), .ZN(G1344gat));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n834), .A2(KEYINPUT119), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n800), .B1(new_n834), .B2(KEYINPUT119), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n842), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n774), .B1(new_n885), .B2(new_n498), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n827), .B1(new_n886), .B2(new_n336), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n803), .A2(new_n498), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n336), .B1(new_n890), .B2(new_n830), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT57), .ZN(new_n892));
  OAI211_X1 g691(.A(KEYINPUT120), .B(new_n827), .C1(new_n886), .C2(new_n336), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n889), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n610), .A3(new_n859), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n882), .B1(new_n895), .B2(G148gat), .ZN(new_n896));
  AOI211_X1 g695(.A(KEYINPUT59), .B(new_n288), .C1(new_n847), .C2(new_n610), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n610), .A2(new_n288), .ZN(new_n898));
  OAI22_X1  g697(.A1(new_n896), .A2(new_n897), .B1(new_n851), .B2(new_n898), .ZN(G1345gat));
  AND2_X1   g698(.A1(new_n847), .A2(new_n679), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n679), .A2(new_n295), .ZN(new_n901));
  OAI22_X1  g700(.A1(new_n900), .A2(new_n295), .B1(new_n851), .B2(new_n901), .ZN(G1346gat));
  NOR2_X1   g701(.A1(new_n667), .A2(new_n296), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n849), .A2(new_n850), .A3(new_n577), .ZN(new_n904));
  AOI22_X1  g703(.A1(new_n847), .A2(new_n903), .B1(new_n904), .B2(new_n296), .ZN(G1347gat));
  NOR2_X1   g704(.A1(new_n367), .A2(new_n396), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT122), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n907), .A2(new_n279), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n805), .A2(new_n908), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n909), .A2(new_n221), .A3(new_n645), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n868), .A2(new_n397), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n911), .A2(KEYINPUT121), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(KEYINPUT121), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n809), .A2(new_n367), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n711), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n910), .B1(new_n918), .B2(new_n221), .ZN(G1348gat));
  OAI21_X1  g718(.A(G176gat), .B1(new_n909), .B2(new_n712), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n610), .A2(new_n222), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n916), .B2(new_n921), .ZN(G1349gat));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n923), .B1(new_n909), .B2(new_n498), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n805), .A2(KEYINPUT123), .A3(new_n679), .A4(new_n908), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(G183gat), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n679), .A2(new_n215), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n916), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT60), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT60), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n926), .B(new_n930), .C1(new_n916), .C2(new_n927), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1350gat));
  NAND3_X1  g731(.A1(new_n917), .A2(new_n216), .A3(new_n577), .ZN(new_n933));
  OAI21_X1  g732(.A(G190gat), .B1(new_n909), .B2(new_n667), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT61), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1351gat));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n937));
  XOR2_X1   g736(.A(KEYINPUT124), .B(G197gat), .Z(new_n938));
  NAND2_X1  g737(.A1(new_n907), .A2(new_n659), .ZN(new_n939));
  AOI22_X1  g738(.A1(new_n887), .A2(new_n888), .B1(KEYINPUT57), .B2(new_n891), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(new_n893), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n938), .B1(new_n941), .B2(new_n711), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n658), .A2(new_n336), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n435), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n944), .B1(new_n912), .B2(new_n913), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n945), .A2(new_n711), .A3(new_n938), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n937), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n945), .A2(new_n711), .A3(new_n938), .ZN(new_n948));
  AOI211_X1 g747(.A(new_n645), .B(new_n939), .C1(new_n940), .C2(new_n893), .ZN(new_n949));
  OAI211_X1 g748(.A(KEYINPUT125), .B(new_n948), .C1(new_n949), .C2(new_n938), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n947), .A2(new_n950), .ZN(G1352gat));
  NOR2_X1   g750(.A1(new_n712), .A2(G204gat), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n945), .A2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n953), .B(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(new_n941), .ZN(new_n956));
  OAI21_X1  g755(.A(G204gat), .B1(new_n956), .B2(new_n712), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(G1353gat));
  NAND3_X1  g757(.A1(new_n945), .A2(new_n305), .A3(new_n679), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n894), .A2(new_n659), .A3(new_n679), .A4(new_n907), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n960), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT63), .B1(new_n960), .B2(G211gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(G1354gat));
  INV_X1    g762(.A(new_n944), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n914), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n306), .B1(new_n965), .B2(new_n667), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(KEYINPUT126), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n968), .B(new_n306), .C1(new_n965), .C2(new_n667), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n577), .A2(G218gat), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n970), .B(KEYINPUT127), .ZN(new_n971));
  AOI22_X1  g770(.A1(new_n967), .A2(new_n969), .B1(new_n941), .B2(new_n971), .ZN(G1355gat));
endmodule


