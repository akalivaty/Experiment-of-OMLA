//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1274, new_n1275, new_n1276, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1350, new_n1351, new_n1352, new_n1353;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n211), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT67), .Z(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  AND2_X1   g0024(.A1(KEYINPUT66), .A2(G77), .ZN(new_n225));
  NOR2_X1   g0025(.A1(KEYINPUT66), .A2(G77), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n223), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT65), .B(G238), .Z(new_n231));
  INV_X1    g0031(.A(G68), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n229), .B(new_n230), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n213), .B1(new_n228), .B2(new_n233), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n216), .B(new_n221), .C1(new_n234), .C2(KEYINPUT1), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n234), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT68), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NOR2_X1   g0052(.A1(KEYINPUT73), .A2(KEYINPUT10), .ZN(new_n253));
  OAI21_X1  g0053(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n211), .A2(G33), .ZN(new_n256));
  OAI21_X1  g0056(.A(KEYINPUT70), .B1(G20), .B2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NOR3_X1   g0058(.A1(KEYINPUT70), .A2(G20), .A3(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G150), .ZN(new_n261));
  OAI221_X1 g0061(.A(new_n254), .B1(new_n255), .B2(new_n256), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT69), .ZN(new_n263));
  NAND3_X1  g0063(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n263), .B1(new_n264), .B2(new_n219), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(new_n263), .A3(new_n219), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n267), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n270), .A2(new_n272), .A3(new_n265), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n273), .B(G50), .C1(G1), .C2(new_n211), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n201), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n269), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT72), .ZN(new_n277));
  OR2_X1    g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n277), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(new_n279), .A3(KEYINPUT9), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G1), .A3(G13), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G274), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n282), .A2(new_n284), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n287), .A2(G226), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT3), .ZN(new_n289));
  INV_X1    g0089(.A(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(G222), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(G1698), .ZN(new_n296));
  INV_X1    g0096(.A(G223), .ZN(new_n297));
  OAI221_X1 g0097(.A(new_n295), .B1(new_n227), .B2(new_n293), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n299));
  AOI211_X1 g0099(.A(new_n285), .B(new_n288), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G200), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(G190), .ZN(new_n304));
  NAND2_X1  g0104(.A1(KEYINPUT73), .A2(KEYINPUT10), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n280), .A2(new_n303), .A3(new_n304), .A4(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(KEYINPUT9), .B1(new_n278), .B2(new_n279), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n253), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n309));
  INV_X1    g0109(.A(new_n307), .ZN(new_n310));
  INV_X1    g0110(.A(new_n253), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .A4(new_n280), .ZN(new_n312));
  INV_X1    g0112(.A(G179), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n300), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n314), .B(new_n276), .C1(G169), .C2(new_n300), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n308), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n255), .B1(new_n210), .B2(G20), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n273), .A2(new_n317), .B1(new_n255), .B2(new_n272), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT16), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n291), .A2(new_n211), .A3(new_n292), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT7), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n291), .A2(KEYINPUT7), .A3(new_n211), .A4(new_n292), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n232), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(G58), .B(G68), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G20), .ZN(new_n326));
  INV_X1    g0126(.A(G159), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n326), .B1(new_n260), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n319), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(KEYINPUT3), .A2(G33), .ZN(new_n330));
  NOR2_X1   g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT7), .B1(new_n332), .B2(new_n211), .ZN(new_n333));
  INV_X1    g0133(.A(new_n323), .ZN(new_n334));
  OAI21_X1  g0134(.A(G68), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n259), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n257), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n337), .A2(G159), .B1(new_n325), .B2(G20), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n335), .A2(KEYINPUT16), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n264), .A2(new_n219), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n329), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(G223), .B(new_n294), .C1(new_n330), .C2(new_n331), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT75), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n293), .A2(KEYINPUT75), .A3(G223), .A4(new_n294), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G33), .A2(G87), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n293), .A2(G226), .A3(G1698), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n344), .A2(new_n345), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n299), .ZN(new_n349));
  INV_X1    g0149(.A(G232), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n350), .A2(new_n286), .B1(new_n283), .B2(new_n284), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(G200), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  AOI211_X1 g0153(.A(G190), .B(new_n351), .C1(new_n348), .C2(new_n299), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n318), .B(new_n341), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT17), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G190), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n349), .A2(new_n358), .A3(new_n352), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n351), .B1(new_n348), .B2(new_n299), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n359), .B1(G200), .B2(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n361), .A2(KEYINPUT17), .A3(new_n318), .A4(new_n341), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n349), .A2(G179), .A3(new_n352), .ZN(new_n365));
  INV_X1    g0165(.A(G169), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n365), .B1(new_n366), .B2(new_n360), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n341), .A2(new_n318), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT18), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT76), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n367), .A2(new_n368), .A3(KEYINPUT18), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n372), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n364), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n260), .A2(new_n201), .ZN(new_n378));
  INV_X1    g0178(.A(G77), .ZN(new_n379));
  OAI22_X1  g0179(.A1(new_n256), .A2(new_n379), .B1(new_n211), .B2(G68), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n268), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT11), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n268), .B(KEYINPUT11), .C1(new_n378), .C2(new_n380), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT12), .B1(new_n271), .B2(G68), .ZN(new_n385));
  OR3_X1    g0185(.A1(new_n271), .A2(KEYINPUT12), .A3(G68), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n272), .A2(new_n340), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n232), .B1(new_n210), .B2(G20), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n385), .A2(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n383), .A2(new_n384), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT74), .ZN(new_n391));
  XNOR2_X1  g0191(.A(new_n390), .B(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT14), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n293), .A2(G232), .A3(G1698), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n293), .A2(G226), .A3(new_n294), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G97), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n299), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n285), .B1(G238), .B2(new_n287), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT13), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n400), .B1(new_n398), .B2(new_n399), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n393), .B(G169), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n398), .A2(new_n399), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT13), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(G179), .A3(new_n401), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n401), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n393), .B1(new_n409), .B2(G169), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n392), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(G200), .B1(new_n402), .B2(new_n403), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n406), .A2(G190), .A3(new_n401), .ZN(new_n413));
  INV_X1    g0213(.A(new_n390), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n340), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n271), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n379), .B1(new_n210), .B2(G20), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n227), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n418), .A2(new_n420), .B1(new_n421), .B2(new_n271), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n260), .A2(new_n255), .ZN(new_n423));
  XNOR2_X1  g0223(.A(KEYINPUT15), .B(G87), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n227), .A2(new_n211), .B1(new_n424), .B2(new_n256), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n340), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n426), .A2(KEYINPUT71), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(KEYINPUT71), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n422), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n293), .A2(G232), .A3(new_n294), .ZN(new_n431));
  OAI221_X1 g0231(.A(new_n431), .B1(new_n207), .B2(new_n293), .C1(new_n296), .C2(new_n231), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n299), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n285), .B1(G244), .B2(new_n287), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(new_n313), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n434), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n366), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n430), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(G200), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n429), .B(new_n439), .C1(new_n358), .C2(new_n436), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NOR4_X1   g0242(.A1(new_n316), .A2(new_n377), .A3(new_n416), .A4(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(G244), .B(new_n294), .C1(new_n330), .C2(new_n331), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT77), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n445), .A2(KEYINPUT4), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n293), .A2(G244), .A3(new_n294), .A4(new_n446), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n293), .A2(G250), .A3(G1698), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G283), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n448), .A2(new_n449), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n299), .ZN(new_n453));
  INV_X1    g0253(.A(G274), .ZN(new_n454));
  INV_X1    g0254(.A(new_n219), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(new_n281), .ZN(new_n456));
  INV_X1    g0256(.A(G41), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n210), .B(G45), .C1(new_n457), .C2(KEYINPUT5), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT5), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT78), .B1(new_n460), .B2(G41), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT78), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n462), .A2(new_n457), .A3(KEYINPUT5), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n456), .A2(new_n459), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n460), .A2(G41), .ZN(new_n465));
  OAI211_X1 g0265(.A(G257), .B(new_n282), .C1(new_n458), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n453), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n366), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT6), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n471), .A2(new_n206), .A3(G107), .ZN(new_n472));
  XNOR2_X1  g0272(.A(G97), .B(G107), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n472), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  OAI22_X1  g0274(.A1(new_n474), .A2(new_n211), .B1(new_n379), .B2(new_n260), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n207), .B1(new_n322), .B2(new_n323), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n340), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n210), .A2(G33), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n273), .A2(G97), .A3(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n271), .A2(G97), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n464), .A2(new_n313), .A3(new_n466), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n453), .A2(new_n483), .A3(KEYINPUT80), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT80), .B1(new_n453), .B2(new_n483), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n470), .B(new_n482), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT81), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n453), .A2(new_n483), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT80), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n453), .A2(new_n483), .A3(KEYINPUT80), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT81), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n492), .A2(new_n493), .A3(new_n470), .A4(new_n482), .ZN(new_n494));
  INV_X1    g0294(.A(new_n482), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n467), .B1(new_n452), .B2(new_n299), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G190), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT79), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n469), .B2(G200), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n496), .A2(KEYINPUT79), .A3(new_n301), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n495), .B(new_n497), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n487), .A2(new_n494), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G116), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n264), .A2(new_n219), .B1(G20), .B2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n451), .B(new_n211), .C1(G33), .C2(new_n206), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n504), .A2(KEYINPUT20), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT20), .B1(new_n504), .B2(new_n505), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n478), .A2(G116), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n418), .A2(new_n509), .B1(G116), .B2(new_n271), .ZN(new_n510));
  OAI21_X1  g0310(.A(G169), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n282), .B1(new_n458), .B2(new_n465), .ZN(new_n512));
  INV_X1    g0312(.A(G270), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n460), .A2(G41), .ZN(new_n514));
  INV_X1    g0314(.A(G45), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(G1), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n461), .A2(new_n463), .A3(new_n514), .A4(new_n516), .ZN(new_n517));
  OAI22_X1  g0317(.A1(new_n512), .A2(new_n513), .B1(new_n517), .B2(new_n283), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT85), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n299), .B1(new_n293), .B2(G303), .ZN(new_n520));
  INV_X1    g0320(.A(G257), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n294), .ZN(new_n522));
  INV_X1    g0322(.A(G264), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G1698), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n522), .A2(new_n524), .B1(new_n291), .B2(new_n292), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n519), .B1(new_n520), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(G303), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n282), .B1(new_n332), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n522), .A2(new_n524), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n293), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(KEYINPUT85), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n518), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n511), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n526), .A2(new_n531), .ZN(new_n534));
  INV_X1    g0334(.A(new_n518), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n534), .A2(G179), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n504), .A2(new_n505), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT20), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n504), .A2(KEYINPUT20), .A3(new_n505), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n509), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n387), .A2(new_n542), .B1(new_n503), .B2(new_n272), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n533), .A2(KEYINPUT21), .B1(new_n536), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n534), .A2(new_n535), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n544), .B1(new_n546), .B2(G200), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n358), .B2(new_n546), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n533), .A2(KEYINPUT86), .A3(KEYINPUT21), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT86), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n366), .B1(new_n541), .B2(new_n543), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT21), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n545), .B(new_n548), .C1(new_n549), .C2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n502), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(G33), .A2(G116), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(G20), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT23), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n211), .B2(G107), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n558), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n211), .B(G87), .C1(new_n330), .C2(new_n331), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n563), .A2(KEYINPUT22), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n563), .A2(KEYINPUT22), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT24), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT24), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n568), .B(new_n562), .C1(new_n564), .C2(new_n565), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n417), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n271), .A2(G107), .ZN(new_n571));
  XNOR2_X1  g0371(.A(new_n571), .B(KEYINPUT25), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n266), .A2(new_n271), .A3(new_n267), .A4(new_n478), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n572), .B1(new_n207), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT87), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n521), .A2(G1698), .ZN(new_n577));
  OAI221_X1 g0377(.A(new_n577), .B1(G250), .B2(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n578));
  NAND2_X1  g0378(.A1(G33), .A2(G294), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n282), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(G264), .B(new_n282), .C1(new_n458), .C2(new_n465), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n576), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(G250), .A2(G1698), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n521), .B2(G1698), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n585), .A2(new_n293), .B1(G33), .B2(G294), .ZN(new_n586));
  OAI211_X1 g0386(.A(KEYINPUT87), .B(new_n581), .C1(new_n586), .C2(new_n282), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n583), .A2(new_n464), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n588), .A2(KEYINPUT88), .A3(new_n301), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n581), .B1(new_n586), .B2(new_n282), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n517), .A2(new_n283), .ZN(new_n591));
  OR3_X1    g0391(.A1(new_n590), .A2(G190), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT88), .B1(new_n588), .B2(new_n301), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n575), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n591), .A2(new_n313), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n583), .A2(new_n587), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(G169), .B1(new_n590), .B2(new_n591), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n570), .B2(new_n574), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(G250), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n515), .B2(G1), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n210), .A2(new_n454), .A3(G45), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n282), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(G238), .A2(G1698), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n224), .B2(G1698), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n607), .A2(new_n293), .B1(G33), .B2(G116), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n313), .B(new_n605), .C1(new_n608), .C2(new_n282), .ZN(new_n609));
  INV_X1    g0409(.A(G238), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n294), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n224), .A2(G1698), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n611), .B(new_n612), .C1(new_n330), .C2(new_n331), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n282), .B1(new_n613), .B2(new_n557), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n282), .A2(new_n603), .A3(new_n604), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n366), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n609), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT19), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n211), .B1(new_n396), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(G87), .B2(new_n208), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n211), .B(G68), .C1(new_n330), .C2(new_n331), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n618), .B1(new_n256), .B2(new_n206), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n340), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n424), .A2(new_n272), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n624), .B(new_n625), .C1(new_n424), .C2(new_n573), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n617), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT83), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n613), .A2(new_n557), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n615), .B1(new_n629), .B2(new_n299), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n628), .B1(new_n630), .B2(G190), .ZN(new_n631));
  NOR4_X1   g0431(.A1(new_n614), .A2(KEYINPUT83), .A3(new_n615), .A4(new_n358), .ZN(new_n632));
  OAI22_X1  g0432(.A1(new_n631), .A2(new_n632), .B1(new_n301), .B2(new_n630), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT82), .ZN(new_n634));
  INV_X1    g0434(.A(G87), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n634), .B1(new_n573), .B2(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n273), .A2(KEYINPUT82), .A3(G87), .A4(new_n478), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n623), .A2(new_n340), .B1(new_n272), .B2(new_n424), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n627), .B1(new_n633), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT84), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n630), .A2(new_n301), .ZN(new_n644));
  OAI211_X1 g0444(.A(G190), .B(new_n605), .C1(new_n608), .C2(new_n282), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT83), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n630), .A2(new_n628), .A3(G190), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n624), .A2(new_n625), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n636), .B2(new_n637), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n651), .A2(KEYINPUT84), .A3(new_n627), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n643), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n443), .A2(new_n556), .A3(new_n601), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n654), .B(KEYINPUT89), .ZN(G372));
  NAND2_X1  g0455(.A1(new_n487), .A2(new_n494), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n656), .A2(new_n653), .A3(KEYINPUT26), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n486), .B2(new_n641), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n487), .A2(new_n494), .A3(new_n501), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n545), .B(new_n600), .C1(new_n549), .C2(new_n554), .ZN(new_n662));
  INV_X1    g0462(.A(new_n594), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n663), .A2(new_n592), .A3(new_n589), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n641), .B1(new_n664), .B2(new_n575), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n661), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n660), .A2(new_n627), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n443), .A2(new_n667), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n367), .A2(new_n368), .A3(KEYINPUT18), .ZN(new_n669));
  AOI21_X1  g0469(.A(KEYINPUT18), .B1(new_n367), .B2(new_n368), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n415), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n411), .B1(new_n672), .B2(new_n438), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n671), .B1(new_n673), .B2(new_n364), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n308), .A2(new_n312), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n315), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n668), .A2(new_n677), .ZN(G369));
  NAND3_X1  g0478(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT90), .ZN(new_n681));
  INV_X1    g0481(.A(G213), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n679), .B2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G343), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n601), .B1(new_n575), .B2(new_n686), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n600), .A2(new_n686), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n545), .B1(new_n549), .B2(new_n554), .ZN(new_n691));
  INV_X1    g0491(.A(new_n555), .ZN(new_n692));
  INV_X1    g0492(.A(new_n686), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n544), .ZN(new_n694));
  MUX2_X1   g0494(.A(new_n691), .B(new_n692), .S(new_n694), .Z(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G330), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n690), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n691), .A2(new_n595), .A3(new_n600), .A4(new_n686), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT91), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n600), .A2(new_n693), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n699), .B1(new_n698), .B2(new_n700), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n697), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT92), .ZN(G399));
  INV_X1    g0505(.A(new_n214), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n217), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n486), .A2(new_n641), .A3(new_n658), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n656), .A2(new_n653), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(new_n658), .ZN(new_n715));
  INV_X1    g0515(.A(new_n641), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n662), .A2(new_n595), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n627), .B1(new_n717), .B2(new_n502), .ZN(new_n718));
  OAI211_X1 g0518(.A(KEYINPUT29), .B(new_n686), .C1(new_n715), .C2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT93), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT29), .B1(new_n667), .B2(new_n686), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(G330), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n556), .A2(new_n601), .A3(new_n653), .A4(new_n686), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n583), .A2(new_n587), .A3(new_n630), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(new_n536), .A3(new_n496), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n725), .A2(new_n536), .A3(KEYINPUT30), .A4(new_n496), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n532), .A2(G179), .A3(new_n630), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(new_n469), .A3(new_n588), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n728), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n693), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(KEYINPUT31), .B1(new_n732), .B2(new_n693), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n723), .B1(new_n724), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(KEYINPUT26), .B1(new_n656), .B2(new_n653), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n666), .B(new_n627), .C1(new_n739), .C2(new_n713), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT93), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n740), .A2(new_n741), .A3(KEYINPUT29), .A4(new_n686), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n722), .A2(KEYINPUT94), .A3(new_n738), .A4(new_n742), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n738), .B(new_n742), .C1(new_n720), .C2(new_n721), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT94), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n712), .B1(new_n747), .B2(G1), .ZN(G364));
  INV_X1    g0548(.A(new_n696), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n211), .A2(G13), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n210), .B1(new_n750), .B2(G45), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n707), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(G330), .B2(new_n695), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n219), .B1(G20), .B2(new_n366), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR4_X1   g0557(.A1(new_n211), .A2(new_n301), .A3(G179), .A4(G190), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n207), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n211), .A2(new_n313), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G190), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR4_X1   g0564(.A1(new_n211), .A2(new_n358), .A3(new_n301), .A4(G179), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n764), .A2(new_n232), .B1(new_n635), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n762), .A2(new_n358), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n760), .B(new_n767), .C1(G50), .C2(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n358), .A2(G179), .A3(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n211), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT95), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G97), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G190), .A2(G200), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(G20), .A3(new_n313), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n327), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT32), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n761), .A2(G190), .A3(new_n301), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n293), .B1(new_n778), .B2(new_n202), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n761), .A2(new_n774), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n779), .B1(new_n421), .B2(new_n781), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n769), .A2(new_n773), .A3(new_n777), .A4(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n771), .ZN(new_n784));
  AOI22_X1  g0584(.A1(G294), .A2(new_n784), .B1(new_n768), .B2(G326), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT96), .ZN(new_n786));
  XNOR2_X1  g0586(.A(KEYINPUT33), .B(G317), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT97), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n764), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(new_n788), .B2(new_n787), .ZN(new_n790));
  INV_X1    g0590(.A(new_n778), .ZN(new_n791));
  INV_X1    g0591(.A(new_n775), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n791), .A2(G322), .B1(G329), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G311), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n793), .B(new_n332), .C1(new_n794), .C2(new_n780), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n766), .A2(new_n527), .B1(new_n759), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n786), .A2(new_n790), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n757), .B1(new_n783), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n706), .A2(new_n332), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G355), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(G116), .B2(new_n214), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n248), .A2(new_n515), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n706), .A2(new_n293), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n515), .B2(new_n218), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n803), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G13), .A2(G33), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(G20), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n756), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n753), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n800), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n811), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n695), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n755), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(G396));
  NAND2_X1  g0619(.A1(new_n441), .A2(new_n686), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n667), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n627), .ZN(new_n823));
  AND3_X1   g0623(.A1(new_n662), .A2(new_n595), .A3(new_n716), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n823), .B1(new_n824), .B2(new_n661), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n693), .B1(new_n825), .B2(new_n660), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n438), .A2(new_n693), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n440), .B1(new_n429), .B2(new_n686), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n827), .B1(new_n438), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n822), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n738), .ZN(new_n831));
  INV_X1    g0631(.A(new_n753), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n822), .B(new_n737), .C1(new_n826), .C2(new_n829), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n756), .A2(new_n809), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n832), .B1(new_n379), .B2(new_n835), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n791), .A2(G143), .B1(new_n781), .B2(G159), .ZN(new_n837));
  INV_X1    g0637(.A(new_n768), .ZN(new_n838));
  INV_X1    g0638(.A(G137), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n837), .B1(new_n838), .B2(new_n839), .C1(new_n261), .C2(new_n764), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT34), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n759), .A2(new_n232), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n845), .B1(new_n201), .B2(new_n766), .C1(new_n202), .C2(new_n771), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n332), .B1(new_n792), .B2(G132), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT99), .ZN(new_n848));
  NOR4_X1   g0648(.A1(new_n842), .A2(new_n843), .A3(new_n846), .A4(new_n848), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n780), .A2(new_n503), .B1(new_n775), .B2(new_n794), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n293), .B(new_n850), .C1(G294), .C2(new_n791), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n759), .A2(new_n635), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(G303), .B2(new_n768), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n763), .A2(G283), .B1(G107), .B2(new_n765), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n851), .A2(new_n773), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT98), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n855), .A2(new_n856), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n849), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n836), .B1(new_n757), .B2(new_n859), .C1(new_n829), .C2(new_n810), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n834), .A2(KEYINPUT100), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT100), .B1(new_n834), .B2(new_n860), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(G384));
  INV_X1    g0664(.A(new_n474), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n865), .A2(KEYINPUT35), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(KEYINPUT35), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n866), .A2(G116), .A3(new_n220), .A4(new_n867), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT36), .Z(new_n869));
  OAI211_X1 g0669(.A(new_n421), .B(new_n218), .C1(new_n202), .C2(new_n232), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n201), .A2(G68), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n210), .B(G13), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n329), .A2(new_n268), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n339), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n318), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT101), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(new_n685), .ZN(new_n878));
  INV_X1    g0678(.A(new_n318), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n874), .B2(new_n339), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT101), .B1(new_n880), .B2(new_n684), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n377), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n876), .A2(new_n367), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n878), .A2(new_n884), .A3(new_n881), .A4(new_n355), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(KEYINPUT37), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n368), .A2(new_n685), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n369), .A2(new_n887), .A3(new_n355), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n883), .A2(new_n890), .A3(KEYINPUT38), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n669), .A2(KEYINPUT76), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(new_n375), .A3(new_n371), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n894), .A2(new_n364), .B1(new_n878), .B2(new_n881), .ZN(new_n895));
  INV_X1    g0695(.A(new_n889), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n885), .B2(KEYINPUT37), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n892), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n891), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(G169), .B1(new_n402), .B2(new_n403), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(KEYINPUT14), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(new_n407), .A3(new_n404), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n392), .B(new_n693), .C1(new_n902), .C2(new_n672), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n392), .A2(new_n693), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n411), .A2(new_n415), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n829), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n724), .B2(new_n736), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n899), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT40), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n724), .A2(new_n736), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n828), .A2(new_n438), .ZN(new_n913));
  INV_X1    g0713(.A(new_n827), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n905), .B2(new_n903), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n912), .A2(new_n916), .A3(KEYINPUT40), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT102), .ZN(new_n919));
  INV_X1    g0719(.A(new_n887), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n671), .B2(new_n363), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n369), .A2(new_n887), .A3(new_n355), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT37), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n889), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n919), .B1(new_n925), .B2(new_n892), .ZN(new_n926));
  AOI211_X1 g0726(.A(KEYINPUT102), .B(KEYINPUT38), .C1(new_n921), .C2(new_n924), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n891), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n918), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n911), .A2(G330), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n443), .A2(new_n737), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT104), .Z(new_n933));
  AOI22_X1  g0733(.A1(new_n909), .A2(new_n910), .B1(new_n918), .B2(new_n928), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(new_n443), .A3(new_n912), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT105), .Z(new_n937));
  INV_X1    g0737(.A(KEYINPUT39), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n928), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n902), .A2(new_n392), .A3(new_n686), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n891), .A2(new_n898), .A3(KEYINPUT39), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n669), .A2(new_n670), .A3(new_n685), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n827), .B1(new_n667), .B2(new_n821), .ZN(new_n945));
  INV_X1    g0745(.A(new_n906), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n944), .B1(new_n947), .B2(new_n899), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT103), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n943), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n949), .B1(new_n943), .B2(new_n948), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n742), .B1(new_n720), .B2(new_n721), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n676), .B1(new_n953), .B2(new_n443), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n952), .B(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(KEYINPUT106), .B1(new_n937), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n937), .A2(new_n955), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n956), .B(new_n957), .C1(new_n210), .C2(new_n750), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n937), .A2(KEYINPUT106), .A3(new_n955), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n873), .B1(new_n958), .B2(new_n959), .ZN(G367));
  INV_X1    g0760(.A(new_n697), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n693), .A2(new_n482), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n487), .A2(new_n494), .A3(new_n501), .A4(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n486), .A2(new_n686), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n701), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n965), .B1(new_n966), .B2(new_n702), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT45), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g0769(.A(KEYINPUT45), .B(new_n965), .C1(new_n966), .C2(new_n702), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n965), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n703), .A2(new_n701), .A3(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT44), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n703), .A2(KEYINPUT44), .A3(new_n701), .A4(new_n972), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n961), .B1(new_n971), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n971), .A2(new_n977), .A3(new_n961), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n691), .A2(new_n686), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n698), .B1(new_n689), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(new_n696), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n747), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n707), .B(KEYINPUT41), .Z(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n752), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n650), .A2(new_n686), .ZN(new_n989));
  MUX2_X1   g0789(.A(new_n641), .B(new_n627), .S(new_n989), .Z(new_n990));
  INV_X1    g0790(.A(KEYINPUT43), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT107), .Z(new_n993));
  NOR2_X1   g0793(.A1(new_n972), .A2(new_n600), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n994), .A2(new_n656), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n995), .A2(new_n693), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n965), .A2(new_n601), .A3(new_n982), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT42), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n993), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n990), .A2(new_n991), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n961), .A2(new_n972), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n990), .A2(new_n811), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n812), .B1(new_n214), .B2(new_n424), .C1(new_n806), .C2(new_n243), .ZN(new_n1005));
  INV_X1    g0805(.A(G294), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n764), .A2(new_n1006), .B1(new_n206), .B2(new_n759), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n791), .A2(G303), .B1(new_n781), .B2(G283), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n765), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1009));
  XOR2_X1   g0809(.A(KEYINPUT108), .B(G317), .Z(new_n1010));
  AOI21_X1  g0810(.A(new_n293), .B1(new_n792), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n838), .A2(new_n794), .B1(new_n207), .B2(new_n771), .ZN(new_n1013));
  AOI21_X1  g0813(.A(KEYINPUT46), .B1(new_n765), .B2(G116), .ZN(new_n1014));
  OR4_X1    g0814(.A1(new_n1007), .A2(new_n1012), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n778), .A2(new_n261), .B1(new_n780), .B2(new_n201), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(KEYINPUT109), .B(G137), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n332), .B(new_n1016), .C1(new_n792), .C2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n772), .A2(G68), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n768), .A2(G143), .B1(new_n421), .B2(new_n758), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n763), .A2(G159), .B1(G58), .B2(new_n765), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1015), .A2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT47), .Z(new_n1025));
  OAI211_X1 g0825(.A(new_n753), .B(new_n1005), .C1(new_n1025), .C2(new_n757), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n988), .A2(new_n1003), .B1(new_n1004), .B2(new_n1026), .ZN(G387));
  AOI21_X1  g0827(.A(new_n984), .B1(new_n743), .B2(new_n746), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1028), .A2(new_n708), .ZN(new_n1029));
  AND3_X1   g0829(.A1(new_n743), .A2(new_n746), .A3(new_n984), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n984), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n690), .A2(new_n811), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n255), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n201), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT50), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n709), .ZN(new_n1039));
  AOI211_X1 g0839(.A(G45), .B(new_n1039), .C1(G68), .C2(G77), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n806), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1041), .A2(KEYINPUT110), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(KEYINPUT110), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(new_n515), .C2(new_n240), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n801), .A2(new_n1039), .B1(new_n207), .B2(new_n706), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1044), .A2(KEYINPUT111), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n812), .ZN(new_n1047));
  AOI21_X1  g0847(.A(KEYINPUT111), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n753), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n772), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1050), .A2(new_n424), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n778), .A2(new_n201), .B1(new_n780), .B2(new_n232), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n332), .B(new_n1052), .C1(G150), .C2(new_n792), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n768), .A2(G159), .B1(G97), .B2(new_n758), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n766), .A2(new_n227), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n1035), .B2(new_n763), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1051), .A2(new_n1053), .A3(new_n1054), .A4(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n293), .B1(new_n792), .B2(G326), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n766), .A2(new_n1006), .B1(new_n796), .B2(new_n771), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n791), .A2(new_n1010), .B1(new_n781), .B2(G303), .ZN(new_n1060));
  INV_X1    g0860(.A(G322), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1060), .B1(new_n838), .B2(new_n1061), .C1(new_n794), .C2(new_n764), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT48), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1059), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n1063), .B2(new_n1062), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT49), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1058), .B1(new_n503), .B2(new_n759), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1057), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT112), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1049), .B1(new_n1070), .B2(new_n756), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1033), .A2(new_n752), .B1(new_n1034), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1032), .A2(new_n1072), .ZN(G393));
  INV_X1    g0873(.A(new_n980), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1074), .A2(new_n978), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n708), .B1(new_n1028), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT113), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n979), .A2(new_n1077), .A3(new_n980), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1074), .B1(new_n978), .B2(KEYINPUT113), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1076), .B1(new_n1028), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n972), .A2(new_n811), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n812), .B1(new_n206), .B2(new_n214), .C1(new_n806), .C2(new_n251), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n753), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n766), .A2(new_n232), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n852), .B(new_n1085), .C1(G50), .C2(new_n763), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n772), .A2(G77), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n781), .A2(new_n1035), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n332), .B1(new_n792), .B2(G143), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G150), .A2(new_n768), .B1(new_n791), .B2(G159), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT51), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n332), .B1(new_n775), .B2(new_n1061), .C1(new_n780), .C2(new_n1006), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n760), .B(new_n1093), .C1(G283), .C2(new_n765), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(G116), .A2(new_n784), .B1(new_n763), .B2(G303), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1095), .A2(KEYINPUT114), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(KEYINPUT114), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1094), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(G317), .A2(new_n768), .B1(new_n791), .B2(G311), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT52), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1090), .A2(new_n1092), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1084), .B1(new_n1101), .B2(new_n756), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1080), .A2(new_n752), .B1(new_n1082), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1081), .A2(new_n1103), .ZN(G390));
  NAND3_X1  g0904(.A1(new_n737), .A2(new_n829), .A3(new_n906), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n820), .B1(new_n825), .B2(new_n660), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n906), .B1(new_n1106), .B2(new_n827), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n939), .A2(new_n942), .B1(new_n940), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n928), .A2(new_n940), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n686), .B(new_n913), .C1(new_n715), .C2(new_n718), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n946), .B1(new_n1110), .B2(new_n914), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(KEYINPUT115), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n940), .B1(new_n945), .B2(new_n946), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n357), .B(new_n362), .C1(new_n669), .C2(new_n670), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1115), .A2(new_n920), .B1(new_n923), .B2(new_n889), .ZN(new_n1116));
  OAI21_X1  g0916(.A(KEYINPUT102), .B1(new_n1116), .B2(KEYINPUT38), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n925), .A2(new_n919), .A3(new_n892), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(KEYINPUT39), .B1(new_n1119), .B2(new_n891), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n891), .A2(new_n898), .A3(KEYINPUT39), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1114), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1110), .A2(new_n914), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n928), .B(new_n940), .C1(new_n1123), .C2(new_n946), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT115), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1122), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1105), .B1(new_n1113), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1105), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1128), .B1(new_n1129), .B2(KEYINPUT115), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n1127), .A2(new_n751), .A3(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n809), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n778), .A2(new_n503), .B1(new_n780), .B2(new_n206), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n845), .B1(new_n207), .B2(new_n764), .C1(new_n796), .C2(new_n838), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1133), .B(new_n1134), .C1(G294), .C2(new_n792), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n293), .B1(new_n765), .B2(G87), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT117), .Z(new_n1137));
  NAND3_X1  g0937(.A1(new_n1135), .A2(new_n1087), .A3(new_n1137), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n764), .A2(new_n1017), .B1(new_n201), .B2(new_n759), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(G128), .B2(new_n768), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT54), .B(G143), .ZN(new_n1141));
  INV_X1    g0941(.A(G125), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n780), .A2(new_n1141), .B1(new_n775), .B2(new_n1142), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n332), .B(new_n1143), .C1(G132), .C2(new_n791), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n772), .A2(G159), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n765), .A2(G150), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT53), .Z(new_n1147));
  NAND4_X1  g0947(.A1(new_n1140), .A2(new_n1144), .A3(new_n1145), .A4(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n757), .B1(new_n1138), .B2(new_n1148), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n832), .B(new_n1149), .C1(new_n255), .C2(new_n835), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT118), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1132), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1131), .A2(new_n1152), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n1108), .A2(new_n1112), .A3(KEYINPUT115), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1125), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1128), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1130), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n953), .A2(new_n443), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1158), .A2(new_n677), .A3(new_n931), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n641), .A2(new_n642), .ZN(new_n1160));
  AOI21_X1  g0960(.A(KEYINPUT84), .B1(new_n651), .B2(new_n627), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n595), .B(new_n600), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  NOR4_X1   g0962(.A1(new_n1162), .A2(new_n502), .A3(new_n555), .A4(new_n693), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n735), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n733), .ZN(new_n1165));
  OAI211_X1 g0965(.A(G330), .B(new_n829), .C1(new_n1163), .C2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n946), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1123), .A2(new_n1167), .A3(new_n1105), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n945), .B1(new_n1167), .B2(new_n1105), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1159), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1156), .A2(new_n1157), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT116), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(new_n1173), .A3(new_n707), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1171), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1173), .B1(new_n1172), .B2(new_n707), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1153), .B1(new_n1177), .B2(new_n1178), .ZN(G378));
  OAI22_X1  g0979(.A1(new_n206), .A2(new_n764), .B1(new_n838), .B2(new_n503), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n759), .A2(new_n202), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1180), .A2(new_n1055), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n332), .A2(new_n457), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n778), .A2(new_n207), .B1(new_n780), .B2(new_n424), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(G283), .C2(new_n792), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1182), .A2(new_n1020), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT58), .ZN(new_n1187));
  AOI21_X1  g0987(.A(G50), .B1(new_n290), .B2(new_n457), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1186), .A2(new_n1187), .B1(new_n1183), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(G128), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n778), .A2(new_n1190), .B1(new_n780), .B2(new_n839), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G132), .B2(new_n763), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1141), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n768), .A2(G125), .B1(new_n765), .B2(new_n1193), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1192), .B(new_n1194), .C1(new_n1050), .C2(new_n261), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1195), .A2(KEYINPUT59), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(KEYINPUT59), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n758), .A2(G159), .ZN(new_n1198));
  AOI211_X1 g0998(.A(G33), .B(G41), .C1(new_n792), .C2(G124), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1189), .B1(new_n1187), .B2(new_n1186), .C1(new_n1196), .C2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n756), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n832), .B1(new_n201), .B2(new_n835), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n684), .B1(new_n278), .B2(new_n279), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n316), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n316), .A2(new_n1204), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1205), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1202), .B(new_n1203), .C1(new_n1212), .C2(new_n810), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT119), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n943), .A2(new_n948), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(KEYINPUT103), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n943), .A2(new_n948), .A3(new_n949), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1212), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n930), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1212), .B1(new_n934), .B2(G330), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1216), .B(new_n1217), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n934), .A2(G330), .A3(new_n1212), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n930), .A2(new_n1218), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(new_n950), .C2(new_n951), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1221), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1214), .B1(new_n1225), .B2(new_n752), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1113), .A2(new_n1126), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1130), .B1(new_n1227), .B2(new_n1128), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1159), .B1(new_n1228), .B2(new_n1171), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1225), .A2(KEYINPUT57), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n707), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1159), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1172), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT57), .B1(new_n1233), .B2(new_n1225), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1226), .B1(new_n1231), .B2(new_n1234), .ZN(G375));
  OR2_X1    g1035(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1236), .A2(new_n931), .A3(new_n954), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1159), .A2(new_n1170), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n987), .A3(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n946), .A2(new_n809), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n764), .A2(new_n1141), .B1(new_n327), .B2(new_n766), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1181), .B(new_n1241), .C1(G132), .C2(new_n768), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n780), .A2(new_n261), .B1(new_n775), .B2(new_n1190), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n332), .B(new_n1243), .C1(new_n791), .C2(new_n1018), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1242), .B(new_n1244), .C1(new_n201), .C2(new_n1050), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n778), .A2(new_n796), .B1(new_n780), .B2(new_n207), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n293), .B(new_n1246), .C1(G303), .C2(new_n792), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n768), .A2(G294), .B1(G77), .B2(new_n758), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n763), .A2(G116), .B1(G97), .B2(new_n765), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1051), .A2(new_n1247), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n757), .B1(new_n1245), .B2(new_n1250), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n832), .B(new_n1251), .C1(new_n232), .C2(new_n835), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1240), .A2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n1170), .B2(new_n751), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1239), .A2(new_n1255), .ZN(G381));
  INV_X1    g1056(.A(G375), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1026), .A2(new_n1004), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n744), .B(KEYINPUT94), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n1033), .B2(new_n1075), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n751), .B1(new_n1260), .B2(new_n986), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1002), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1001), .B(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1258), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1153), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n708), .B1(new_n1228), .B2(new_n1171), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1175), .B1(new_n1266), .B2(new_n1173), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1127), .A2(new_n1237), .A3(new_n1130), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT116), .B1(new_n1268), .B2(new_n708), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1265), .B1(new_n1267), .B2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1032), .A2(new_n818), .A3(new_n1072), .ZN(new_n1271));
  NOR4_X1   g1071(.A1(G390), .A2(new_n1271), .A3(G384), .A4(G381), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1257), .A2(new_n1264), .A3(new_n1270), .A4(new_n1272), .ZN(G407));
  NOR2_X1   g1073(.A1(new_n682), .A2(G343), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1257), .A2(new_n1270), .A3(new_n1274), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1275), .B(KEYINPUT120), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(G213), .A3(G407), .ZN(G409));
  NOR3_X1   g1077(.A1(new_n1030), .A2(new_n1028), .A3(new_n708), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1072), .ZN(new_n1279));
  OAI21_X1  g1079(.A(G396), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1271), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1264), .B2(G390), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1081), .A2(new_n1103), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1283), .A2(G387), .ZN(new_n1284));
  OAI21_X1  g1084(.A(KEYINPUT125), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(G387), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1264), .A2(G390), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT125), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1286), .A2(new_n1287), .A3(new_n1288), .A4(new_n1281), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT124), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1290), .B1(new_n1264), .B2(G390), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1283), .A2(G387), .A3(KEYINPUT124), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n1292), .A3(new_n1287), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1281), .ZN(new_n1294));
  AOI22_X1  g1094(.A1(new_n1285), .A2(new_n1289), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1269), .A2(new_n1176), .A3(new_n1174), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n987), .B(new_n1225), .C1(new_n1268), .C2(new_n1159), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1226), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1296), .A2(new_n1298), .A3(new_n1153), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(G375), .B2(new_n1270), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1274), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1159), .A2(new_n1170), .A3(KEYINPUT60), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1302), .A2(new_n707), .ZN(new_n1303));
  OAI21_X1  g1103(.A(KEYINPUT60), .B1(new_n1159), .B2(new_n1170), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1238), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(G384), .B1(new_n1306), .B2(new_n1255), .ZN(new_n1307));
  AOI211_X1 g1107(.A(new_n863), .B(new_n1254), .C1(new_n1303), .C2(new_n1305), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1300), .A2(new_n1301), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(KEYINPUT121), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1233), .A2(KEYINPUT57), .A3(new_n1225), .ZN(new_n1312));
  AOI22_X1  g1112(.A1(new_n1172), .A2(new_n1232), .B1(new_n1224), .B2(new_n1221), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1312), .B(new_n707), .C1(KEYINPUT57), .C2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1314), .A2(G378), .A3(new_n1226), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1274), .B1(new_n1315), .B2(new_n1299), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT121), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1316), .A2(new_n1317), .A3(new_n1309), .ZN(new_n1318));
  AOI21_X1  g1118(.A(KEYINPUT62), .B1(new_n1311), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1310), .A2(KEYINPUT62), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1274), .A2(G2897), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1309), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(KEYINPUT122), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT122), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1309), .A2(new_n1325), .A3(new_n1322), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1324), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1322), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1328), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(KEYINPUT123), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT123), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1331), .B(new_n1328), .C1(new_n1307), .C2(new_n1308), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1330), .A2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1321), .A2(new_n1327), .A3(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT61), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1320), .A2(new_n1335), .A3(new_n1336), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1295), .B1(new_n1319), .B2(new_n1337), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1300), .A2(KEYINPUT63), .A3(new_n1301), .A4(new_n1309), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT126), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1316), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(new_n1309), .ZN(new_n1342));
  AND2_X1   g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1333), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1344));
  AOI211_X1 g1144(.A(KEYINPUT61), .B(new_n1295), .C1(new_n1344), .C2(new_n1327), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT63), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1311), .A2(new_n1318), .A3(new_n1346), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1343), .A2(new_n1345), .A3(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1338), .A2(new_n1348), .ZN(G405));
  NAND2_X1  g1149(.A1(G375), .A2(new_n1270), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1350), .A2(new_n1315), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1309), .A2(KEYINPUT127), .ZN(new_n1352));
  XNOR2_X1  g1152(.A(new_n1351), .B(new_n1352), .ZN(new_n1353));
  XOR2_X1   g1153(.A(new_n1353), .B(new_n1295), .Z(G402));
endmodule


