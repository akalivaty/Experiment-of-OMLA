//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1244, new_n1245, new_n1246, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G244), .ZN(new_n205));
  INV_X1    g0005(.A(G116), .ZN(new_n206));
  INV_X1    g0006(.A(G270), .ZN(new_n207));
  OAI22_X1  g0007(.A1(new_n202), .A2(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  INV_X1    g0010(.A(G97), .ZN(new_n211));
  INV_X1    g0011(.A(G257), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI211_X1 g0013(.A(new_n208), .B(new_n213), .C1(G68), .C2(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G50), .ZN(new_n215));
  INV_X1    g0015(.A(G226), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(KEYINPUT65), .ZN(new_n218));
  AND2_X1   g0018(.A1(new_n217), .A2(KEYINPUT65), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G20), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT66), .Z(new_n223));
  AND2_X1   g0023(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n221), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT64), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  OAI21_X1  g0029(.A(G50), .B1(G58), .B2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NOR4_X1   g0033(.A1(new_n224), .A2(new_n225), .A3(new_n229), .A4(new_n233), .ZN(G361));
  XOR2_X1   g0034(.A(KEYINPUT67), .B(G232), .Z(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n207), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G97), .B(G107), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G87), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n206), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n258));
  OAI21_X1  g0058(.A(KEYINPUT68), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n255), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT68), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G232), .A3(G1698), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G97), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n265), .B(new_n266), .C1(new_n268), .C2(new_n216), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n232), .B1(G33), .B2(G41), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n254), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT13), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  OAI211_X1 g0073(.A(G1), .B(G13), .C1(new_n257), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n252), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G238), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n271), .A2(new_n272), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n272), .B1(new_n271), .B2(new_n277), .ZN(new_n280));
  OAI21_X1  g0080(.A(G169), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT14), .ZN(new_n282));
  INV_X1    g0082(.A(new_n280), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G179), .A3(new_n278), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT14), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n285), .B(G169), .C1(new_n279), .C2(new_n280), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n282), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT69), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(new_n221), .B2(new_n257), .ZN(new_n289));
  NAND4_X1  g0089(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(new_n232), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n291), .B1(new_n251), .B2(G20), .ZN(new_n292));
  INV_X1    g0092(.A(G68), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G20), .ZN(new_n294));
  INV_X1    g0094(.A(G13), .ZN(new_n295));
  NOR3_X1   g0095(.A1(new_n294), .A2(G1), .A3(new_n295), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n292), .A2(G68), .B1(KEYINPUT12), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(KEYINPUT12), .B2(new_n296), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT74), .ZN(new_n299));
  NOR2_X1   g0099(.A1(G20), .A2(G33), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n257), .A2(G20), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OAI221_X1 g0103(.A(new_n294), .B1(new_n301), .B2(new_n215), .C1(new_n303), .C2(new_n202), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n291), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT11), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n287), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n307), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n283), .A2(G190), .A3(new_n278), .ZN(new_n310));
  OAI21_X1  g0110(.A(G200), .B1(new_n279), .B2(new_n280), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n264), .A2(G238), .A3(G1698), .ZN(new_n313));
  OR2_X1    g0113(.A1(KEYINPUT72), .A2(G107), .ZN(new_n314));
  NAND2_X1  g0114(.A1(KEYINPUT72), .A2(G107), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n313), .B1(new_n264), .B2(new_n316), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n262), .B1(new_n260), .B2(new_n261), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G232), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n320), .A2(new_n321), .A3(G1698), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n270), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n254), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n276), .A2(G244), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G190), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT8), .B(G58), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT73), .ZN(new_n330));
  XOR2_X1   g0130(.A(KEYINPUT15), .B(G87), .Z(new_n331));
  AOI22_X1  g0131(.A1(new_n330), .A2(new_n300), .B1(new_n302), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n231), .B2(new_n202), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n295), .A2(new_n231), .A3(G1), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n333), .A2(new_n291), .B1(new_n202), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n292), .A2(G77), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G200), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n328), .B(new_n338), .C1(new_n339), .C2(new_n327), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n308), .A2(new_n312), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G150), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n329), .A2(new_n303), .B1(new_n342), .B2(new_n301), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT70), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI221_X1 g0145(.A(KEYINPUT70), .B1(new_n342), .B2(new_n301), .C1(new_n329), .C2(new_n303), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n345), .B(new_n346), .C1(new_n231), .C2(new_n201), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n291), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT71), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n347), .A2(KEYINPUT71), .A3(new_n291), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n334), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(G50), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n292), .A2(G50), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n352), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT9), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n352), .A2(KEYINPUT9), .A3(new_n355), .A4(new_n356), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n264), .A2(G223), .A3(G1698), .ZN(new_n361));
  INV_X1    g0161(.A(G222), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n361), .B1(new_n202), .B2(new_n264), .C1(new_n268), .C2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n254), .B1(new_n363), .B2(new_n270), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n276), .A2(G226), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(G190), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n365), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(G200), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n359), .A2(new_n360), .A3(new_n366), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT10), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n360), .A2(new_n368), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT10), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n371), .A2(new_n372), .A3(new_n366), .A4(new_n359), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G169), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n367), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G179), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n364), .A2(new_n377), .A3(new_n365), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(new_n357), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT16), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT7), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(new_n264), .B2(G20), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n256), .A2(KEYINPUT76), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT76), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n260), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n261), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n387), .A2(KEYINPUT7), .A3(new_n231), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n293), .B1(new_n383), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G58), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n390), .A2(new_n293), .ZN(new_n391));
  NOR2_X1   g0191(.A1(G58), .A2(G68), .ZN(new_n392));
  OAI21_X1  g0192(.A(G20), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT75), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n300), .A2(G159), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT75), .B(G20), .C1(new_n391), .C2(new_n392), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n381), .B1(new_n389), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n291), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n260), .A2(new_n261), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n401), .A2(new_n382), .A3(new_n231), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n231), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n293), .B1(new_n403), .B2(KEYINPUT7), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n398), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n400), .B1(new_n405), .B2(KEYINPUT16), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n399), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n329), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n408), .A2(new_n334), .ZN(new_n409));
  INV_X1    g0209(.A(new_n292), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n409), .B1(new_n410), .B2(new_n408), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n256), .A2(new_n258), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n216), .A2(G1698), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n413), .B(new_n414), .C1(G223), .C2(G1698), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G33), .A2(G87), .ZN(new_n416));
  XOR2_X1   g0216(.A(new_n416), .B(KEYINPUT77), .Z(new_n417));
  AOI21_X1  g0217(.A(new_n274), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n275), .A2(new_n321), .ZN(new_n419));
  NOR3_X1   g0219(.A1(new_n418), .A2(new_n419), .A3(new_n254), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G200), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(G190), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n407), .A2(new_n412), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT17), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n411), .B1(new_n399), .B2(new_n406), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT17), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n426), .A2(new_n427), .A3(new_n422), .A4(new_n423), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n420), .A2(G179), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n375), .B2(new_n420), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n399), .A2(new_n406), .ZN(new_n431));
  OAI211_X1 g0231(.A(KEYINPUT18), .B(new_n430), .C1(new_n431), .C2(new_n411), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT18), .ZN(new_n433));
  NOR4_X1   g0233(.A1(new_n418), .A2(new_n419), .A3(new_n377), .A4(new_n254), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(new_n421), .B2(G169), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n433), .B1(new_n426), .B2(new_n435), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n425), .A2(new_n428), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n337), .B1(new_n326), .B2(G179), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n327), .A2(G169), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n341), .A2(new_n380), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n259), .A2(G303), .A3(new_n263), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT81), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n413), .A2(new_n445), .A3(G264), .A4(G1698), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n413), .A2(G257), .A3(new_n267), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n260), .A2(new_n261), .A3(G264), .A4(G1698), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT81), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n444), .A2(new_n446), .A3(new_n447), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n270), .ZN(new_n451));
  INV_X1    g0251(.A(G45), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(G1), .ZN(new_n453));
  AND2_X1   g0253(.A1(KEYINPUT5), .A2(G41), .ZN(new_n454));
  NOR2_X1   g0254(.A1(KEYINPUT5), .A2(G41), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OR2_X1    g0256(.A1(new_n456), .A2(new_n253), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n274), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(new_n207), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n451), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT20), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n206), .A2(G20), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n291), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n231), .B1(new_n211), .B2(G33), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G283), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT79), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT79), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(G33), .A3(G283), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n465), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n462), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n470), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n472), .A2(KEYINPUT20), .A3(new_n291), .A4(new_n463), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n463), .A2(G1), .A3(new_n295), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n257), .A2(G1), .ZN(new_n477));
  NOR4_X1   g0277(.A1(new_n291), .A2(new_n206), .A3(new_n334), .A4(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n474), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n461), .A2(new_n480), .A3(G169), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT21), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n461), .A2(new_n480), .A3(KEYINPUT21), .A4(G169), .ZN(new_n484));
  INV_X1    g0284(.A(new_n457), .ZN(new_n485));
  AOI211_X1 g0285(.A(new_n485), .B(new_n459), .C1(new_n450), .C2(new_n270), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(G179), .A3(new_n480), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n451), .A2(G190), .A3(new_n457), .A4(new_n460), .ZN(new_n488));
  AOI211_X1 g0288(.A(new_n475), .B(new_n478), .C1(new_n471), .C2(new_n473), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n488), .B(new_n489), .C1(new_n486), .C2(new_n339), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n483), .A2(new_n484), .A3(new_n487), .A4(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT82), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT24), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT23), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G116), .ZN(new_n495));
  NAND2_X1  g0295(.A1(KEYINPUT22), .A2(G87), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n494), .B(new_n495), .C1(new_n401), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n231), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G20), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n316), .B2(new_n494), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT22), .B1(new_n264), .B2(G87), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n492), .B(new_n493), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT22), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(new_n320), .B2(new_n209), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n501), .B1(new_n497), .B2(new_n231), .ZN(new_n508));
  NAND2_X1  g0308(.A1(KEYINPUT82), .A2(KEYINPUT24), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n492), .A2(new_n493), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n507), .A2(new_n508), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n505), .A2(new_n291), .A3(new_n511), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n291), .A2(new_n334), .A3(new_n477), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G107), .ZN(new_n514));
  INV_X1    g0314(.A(G107), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n334), .A2(new_n515), .ZN(new_n516));
  XOR2_X1   g0316(.A(new_n516), .B(KEYINPUT25), .Z(new_n517));
  NAND3_X1  g0317(.A1(new_n512), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n210), .A2(new_n267), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n212), .A2(G1698), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n260), .A2(new_n519), .A3(new_n261), .A4(new_n520), .ZN(new_n521));
  XNOR2_X1  g0321(.A(KEYINPUT83), .B(G294), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n521), .B1(new_n257), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n270), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n456), .A2(new_n274), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G264), .ZN(new_n526));
  INV_X1    g0326(.A(G190), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n524), .A2(new_n526), .A3(new_n527), .A4(new_n457), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(KEYINPUT84), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n524), .A2(new_n526), .A3(new_n457), .ZN(new_n530));
  OAI211_X1 g0330(.A(KEYINPUT84), .B(new_n528), .C1(new_n530), .C2(G200), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n518), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n491), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n530), .A2(G169), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n377), .B2(new_n530), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n518), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n513), .A2(G87), .ZN(new_n538));
  AOI21_X1  g0338(.A(G87), .B1(new_n314), .B2(new_n315), .ZN(new_n539));
  NAND3_X1  g0339(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n539), .A2(new_n211), .B1(new_n231), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n231), .A2(G33), .A3(G97), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT19), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n293), .A2(G20), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n544), .B1(new_n401), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n291), .B1(new_n541), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n353), .A2(new_n331), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n538), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n260), .A2(new_n261), .A3(G238), .A4(new_n267), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n260), .A2(new_n261), .A3(G244), .A4(G1698), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n554), .A3(new_n495), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n270), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n270), .A2(new_n453), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n557), .A2(G250), .B1(G274), .B2(new_n453), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n339), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n552), .A2(KEYINPUT80), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT80), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n551), .B2(new_n559), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n556), .A2(new_n558), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G190), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n561), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n316), .A2(new_n209), .A3(new_n211), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n540), .A2(new_n231), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n413), .A2(new_n545), .B1(new_n543), .B2(new_n542), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n549), .B1(new_n572), .B2(new_n291), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n513), .A2(new_n331), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n573), .A2(new_n574), .B1(new_n565), .B2(new_n377), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(G169), .B2(new_n565), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n567), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n537), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT4), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(new_n205), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n267), .B(new_n580), .C1(new_n318), .C2(new_n319), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT78), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n264), .A2(KEYINPUT78), .A3(new_n267), .A4(new_n580), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n264), .A2(G250), .A3(G1698), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n260), .A2(new_n261), .A3(G244), .A4(new_n267), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n586), .A2(new_n579), .B1(new_n469), .B2(new_n467), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n583), .A2(new_n584), .A3(new_n585), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n270), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n457), .B1(new_n458), .B2(new_n212), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(G179), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n590), .B1(new_n588), .B2(new_n270), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n375), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n353), .A2(G97), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n513), .A2(G97), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n316), .B1(new_n383), .B2(new_n388), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n301), .A2(new_n202), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT6), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n247), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n515), .A2(KEYINPUT6), .A3(G97), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G20), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n598), .A2(new_n599), .A3(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n596), .B(new_n597), .C1(new_n606), .C2(new_n400), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n594), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n589), .A2(new_n591), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(G200), .ZN(new_n610));
  INV_X1    g0410(.A(new_n316), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT7), .B1(new_n320), .B2(new_n231), .ZN(new_n612));
  INV_X1    g0412(.A(new_n388), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n599), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(new_n615), .A3(new_n604), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n595), .B1(new_n616), .B2(new_n291), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n593), .A2(G190), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n610), .A2(new_n617), .A3(new_n597), .A4(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n608), .A2(new_n619), .ZN(new_n620));
  AND4_X1   g0420(.A1(new_n443), .A2(new_n534), .A3(new_n578), .A4(new_n620), .ZN(G372));
  NAND2_X1  g0421(.A1(new_n558), .A2(KEYINPUT85), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n558), .A2(KEYINPUT85), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n556), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n375), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n575), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n594), .A2(new_n576), .A3(new_n567), .A4(new_n607), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n628), .B1(new_n629), .B2(KEYINPUT26), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT86), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n375), .B1(new_n589), .B2(new_n591), .ZN(new_n632));
  AOI211_X1 g0432(.A(new_n377), .B(new_n590), .C1(new_n588), .C2(new_n270), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n592), .B(KEYINPUT86), .C1(new_n375), .C2(new_n593), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT26), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n625), .A2(G200), .B1(G190), .B2(new_n565), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n638), .A2(new_n552), .B1(new_n575), .B2(new_n626), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n636), .A2(new_n637), .A3(new_n607), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n630), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT87), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n483), .A2(new_n484), .A3(new_n487), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n639), .B1(new_n537), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n608), .A2(new_n619), .ZN(new_n645));
  OR3_X1    g0445(.A1(new_n644), .A2(new_n645), .A3(new_n533), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT87), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n630), .A2(new_n640), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n642), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n443), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n379), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n432), .A2(new_n436), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n287), .A2(new_n307), .B1(new_n312), .B2(new_n440), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n425), .A2(new_n428), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n652), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n651), .B1(new_n656), .B2(new_n374), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n650), .A2(new_n657), .ZN(G369));
  NAND3_X1  g0458(.A1(new_n251), .A2(new_n231), .A3(G13), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT88), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n660), .A2(KEYINPUT88), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n661), .A2(G213), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n489), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n643), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n491), .B2(new_n668), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(KEYINPUT89), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT89), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n537), .A2(new_n667), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  OR3_X1    g0477(.A1(new_n518), .A2(new_n529), .A3(new_n532), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n518), .A2(new_n666), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n537), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n675), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  INV_X1    g0483(.A(new_n537), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n643), .A2(new_n667), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n677), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n682), .A2(new_n688), .ZN(G399));
  NOR2_X1   g0489(.A1(new_n568), .A2(G116), .ZN(new_n690));
  INV_X1    g0490(.A(new_n226), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(G41), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n690), .A2(G1), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n230), .B2(new_n693), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n630), .A2(new_n640), .A3(new_n647), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n647), .B1(new_n630), .B2(new_n640), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n666), .B1(new_n699), .B2(new_n646), .ZN(new_n700));
  OAI21_X1  g0500(.A(KEYINPUT91), .B1(new_n700), .B2(KEYINPUT29), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n629), .A2(KEYINPUT26), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n636), .A2(new_n607), .A3(new_n639), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n627), .B(new_n702), .C1(new_n703), .C2(new_n637), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n644), .A2(new_n645), .A3(new_n533), .ZN(new_n705));
  OAI211_X1 g0505(.A(KEYINPUT29), .B(new_n667), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n649), .A2(new_n667), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT91), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT29), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n701), .A2(new_n706), .A3(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n620), .A2(new_n534), .A3(new_n578), .A4(new_n667), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n593), .A2(new_n565), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n524), .A2(new_n526), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n461), .A2(new_n377), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n714), .A2(KEYINPUT30), .A3(new_n715), .A4(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT30), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n715), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n718), .B1(new_n719), .B2(new_n713), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n625), .A2(new_n461), .A3(new_n377), .ZN(new_n721));
  OR3_X1    g0521(.A1(new_n721), .A2(new_n530), .A3(new_n593), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n717), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n666), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n724), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n724), .A2(KEYINPUT31), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(G330), .A3(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT90), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n725), .A2(new_n726), .A3(KEYINPUT90), .A4(G330), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n711), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n696), .B1(new_n734), .B2(G1), .ZN(G364));
  NOR2_X1   g0535(.A1(new_n295), .A2(G20), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G45), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n737), .A2(KEYINPUT92), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(KEYINPUT92), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n738), .A2(G1), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n692), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G330), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n671), .A2(new_n743), .A3(new_n673), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n675), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G190), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  XOR2_X1   g0548(.A(KEYINPUT33), .B(G317), .Z(new_n749));
  NOR2_X1   g0549(.A1(G179), .A2(G200), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n231), .B1(new_n750), .B2(G190), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n748), .A2(new_n749), .B1(new_n522), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n231), .A2(G190), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n750), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G329), .ZN(new_n756));
  INV_X1    g0556(.A(G311), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n377), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G322), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n231), .A2(new_n527), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n758), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n756), .B1(new_n757), .B2(new_n759), .C1(new_n760), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n339), .A2(G179), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n753), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n752), .B(new_n763), .C1(G283), .C2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n746), .A2(new_n527), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G326), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n761), .A2(new_n764), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n264), .B1(G303), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT93), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n767), .A2(new_n769), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n759), .A2(new_n202), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n751), .A2(new_n211), .ZN(new_n776));
  INV_X1    g0576(.A(G159), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n754), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT32), .ZN(new_n779));
  INV_X1    g0579(.A(new_n768), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n778), .A2(new_n779), .B1(new_n215), .B2(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n776), .B(new_n781), .C1(new_n779), .C2(new_n778), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n320), .B1(G68), .B2(new_n747), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n765), .A2(new_n515), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n770), .A2(new_n209), .ZN(new_n785));
  INV_X1    g0585(.A(new_n762), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n784), .B(new_n785), .C1(G58), .C2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n782), .A2(new_n783), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n774), .B1(new_n775), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n232), .B1(G20), .B2(new_n375), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n246), .A2(G45), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n413), .A2(new_n691), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n791), .B(new_n792), .C1(G45), .C2(new_n230), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n264), .A2(G355), .A3(new_n226), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n793), .B(new_n794), .C1(G116), .C2(new_n226), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G13), .A2(G33), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n790), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n789), .A2(new_n790), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n798), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n741), .B(new_n800), .C1(new_n674), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n745), .A2(new_n802), .ZN(G396));
  INV_X1    g0603(.A(new_n340), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n441), .A2(KEYINPUT95), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT95), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n804), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n649), .A2(new_n667), .A3(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT95), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n440), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n340), .B1(new_n811), .B2(new_n806), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n338), .A2(new_n667), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n812), .A2(new_n813), .B1(new_n441), .B2(new_n667), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n809), .B1(new_n700), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n732), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n731), .B(new_n809), .C1(new_n700), .C2(new_n814), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n816), .A2(new_n817), .A3(new_n742), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n770), .A2(new_n515), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n759), .A2(new_n206), .B1(new_n754), .B2(new_n757), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n819), .B(new_n820), .C1(G294), .C2(new_n786), .ZN(new_n821));
  INV_X1    g0621(.A(G303), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n780), .A2(new_n822), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n776), .B(new_n823), .C1(G283), .C2(new_n747), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n766), .A2(G87), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n821), .A2(new_n824), .A3(new_n320), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n766), .A2(G68), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n215), .B2(new_n770), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(KEYINPUT94), .ZN(new_n829));
  INV_X1    g0629(.A(new_n751), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n401), .B(new_n829), .C1(G58), .C2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n759), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n832), .A2(G159), .B1(G137), .B2(new_n768), .ZN(new_n833));
  INV_X1    g0633(.A(G143), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n833), .B1(new_n834), .B2(new_n762), .C1(new_n342), .C2(new_n748), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT34), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n828), .A2(KEYINPUT94), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n831), .A2(new_n837), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(G132), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n754), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n826), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n790), .A2(new_n796), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n843), .A2(new_n790), .B1(new_n202), .B2(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n741), .B(new_n845), .C1(new_n814), .C2(new_n797), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT96), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n818), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT97), .Z(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G384));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  INV_X1    g0651(.A(new_n664), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n431), .A2(new_n411), .B1(new_n430), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT37), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n853), .A2(new_n854), .A3(new_n424), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n854), .B1(new_n853), .B2(new_n424), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n852), .B1(new_n431), .B2(new_n411), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n654), .B2(new_n652), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n851), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT39), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n853), .A2(new_n854), .A3(new_n424), .ZN(new_n862));
  INV_X1    g0662(.A(new_n398), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n404), .A2(new_n402), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(KEYINPUT16), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n291), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n405), .A2(KEYINPUT16), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n412), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n430), .B2(new_n852), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n869), .A2(new_n424), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n862), .B1(new_n870), .B2(new_n854), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n868), .A2(new_n852), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n871), .B(KEYINPUT38), .C1(new_n437), .C2(new_n872), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n860), .A2(new_n861), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n854), .B1(new_n869), .B2(new_n424), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n855), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n872), .B1(new_n654), .B2(new_n652), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n851), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n861), .B1(new_n878), .B2(new_n873), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT98), .B1(new_n874), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT98), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n860), .A2(new_n873), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n881), .B1(new_n882), .B2(KEYINPUT39), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n308), .A2(new_n666), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n652), .A2(new_n852), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n307), .A2(new_n666), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n308), .A2(new_n312), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n312), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n307), .B(new_n666), .C1(new_n890), .C2(new_n287), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n805), .A2(new_n667), .A3(new_n807), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n892), .B1(new_n809), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n878), .A2(new_n873), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n887), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n886), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n701), .A2(new_n443), .A3(new_n706), .A4(new_n710), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n657), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n897), .B(new_n899), .Z(new_n900));
  NAND2_X1  g0700(.A1(new_n725), .A2(new_n726), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n889), .A2(new_n891), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n902), .A2(new_n814), .A3(new_n882), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT40), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT40), .B1(new_n878), .B2(new_n873), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n902), .A2(new_n906), .A3(new_n814), .A4(new_n903), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n443), .A2(new_n902), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n908), .B(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(G330), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n900), .B(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n251), .B2(new_n736), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n206), .B1(new_n603), .B2(KEYINPUT35), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n232), .A2(new_n231), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n914), .B(new_n915), .C1(KEYINPUT35), .C2(new_n603), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT36), .ZN(new_n917));
  OAI21_X1  g0717(.A(G77), .B1(new_n390), .B2(new_n293), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n918), .A2(new_n230), .B1(G50), .B2(new_n293), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(G1), .A3(new_n295), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n913), .A2(new_n917), .A3(new_n920), .ZN(G367));
  INV_X1    g0721(.A(new_n740), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT45), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n607), .A2(new_n666), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n620), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n636), .A2(new_n607), .A3(new_n666), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n676), .B1(new_n680), .B2(new_n686), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n927), .A2(new_n928), .A3(KEYINPUT101), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT101), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n925), .A2(new_n926), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n930), .B1(new_n688), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n923), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT101), .B1(new_n927), .B2(new_n928), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n688), .A2(new_n930), .A3(new_n931), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(KEYINPUT45), .A3(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT44), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n688), .B2(new_n931), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n927), .A2(new_n928), .A3(KEYINPUT44), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n933), .A2(new_n936), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n681), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n682), .A2(new_n933), .A3(new_n936), .A4(new_n940), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n680), .A2(new_n677), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(new_n686), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT102), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n675), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n949), .A2(new_n675), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n732), .B(new_n711), .C1(new_n944), .C2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT103), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n692), .B(KEYINPUT41), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n954), .B1(new_n953), .B2(new_n955), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n922), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n931), .A2(new_n945), .A3(new_n687), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT42), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n608), .B1(new_n927), .B2(new_n684), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n960), .B1(new_n667), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n552), .A2(new_n667), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n627), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n639), .B2(new_n963), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT99), .Z(new_n966));
  XNOR2_X1  g0766(.A(KEYINPUT100), .B(KEYINPUT43), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n962), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT43), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n970), .B1(new_n971), .B2(new_n966), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n962), .A2(new_n969), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n682), .A2(new_n927), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n958), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n966), .A2(new_n798), .ZN(new_n978));
  INV_X1    g0778(.A(new_n331), .ZN(new_n979));
  INV_X1    g0779(.A(new_n792), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n799), .B1(new_n226), .B2(new_n979), .C1(new_n242), .C2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n832), .A2(G50), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n765), .A2(new_n202), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(G150), .B2(new_n786), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n390), .B2(new_n770), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n751), .A2(new_n293), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(new_n768), .B2(G143), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n777), .B2(new_n748), .ZN(new_n988));
  INV_X1    g0788(.A(G137), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n264), .B1(new_n989), .B2(new_n754), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n985), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n765), .A2(new_n211), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G283), .B2(new_n832), .ZN(new_n993));
  INV_X1    g0793(.A(G317), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n993), .B1(new_n994), .B2(new_n754), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n771), .A2(KEYINPUT46), .A3(G116), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n768), .A2(G311), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n830), .A2(new_n611), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT46), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n770), .B2(new_n206), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n996), .A2(new_n997), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n401), .B1(new_n748), .B2(new_n522), .ZN(new_n1002));
  NOR3_X1   g0802(.A1(new_n995), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n786), .A2(G303), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n982), .A2(new_n991), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT47), .Z(new_n1006));
  AOI21_X1  g0806(.A(new_n742), .B1(new_n1006), .B2(new_n790), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n978), .A2(new_n981), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n977), .A2(new_n1008), .ZN(G387));
  INV_X1    g0809(.A(new_n952), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n734), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n733), .A2(new_n952), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1011), .A2(new_n692), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(new_n740), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n979), .A2(new_n751), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n992), .B(new_n1015), .C1(G159), .C2(new_n768), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n771), .A2(G77), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n759), .A2(new_n293), .B1(new_n754), .B2(new_n342), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G50), .B2(new_n786), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n401), .B1(new_n408), .B2(new_n747), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n762), .A2(new_n994), .B1(new_n759), .B2(new_n822), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n1022), .A2(KEYINPUT104), .B1(G311), .B2(new_n747), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(KEYINPUT104), .B2(new_n1022), .C1(new_n760), .C2(new_n780), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT105), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT48), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n770), .A2(new_n522), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n830), .A2(G283), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT49), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n413), .B1(new_n755), .B2(G326), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n765), .A2(new_n206), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1021), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n330), .A2(new_n215), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1039), .A2(KEYINPUT50), .ZN(new_n1040));
  AOI211_X1 g0840(.A(G116), .B(new_n568), .C1(G68), .C2(G77), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(KEYINPUT50), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n452), .A4(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n980), .B1(new_n239), .B2(G45), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n690), .A2(new_n320), .A3(new_n691), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(G107), .B2(new_n226), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n1038), .A2(new_n790), .B1(new_n799), .B2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1048), .B(new_n741), .C1(new_n945), .C2(new_n801), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT106), .Z(new_n1050));
  NAND3_X1  g0850(.A1(new_n1013), .A2(new_n1014), .A3(new_n1050), .ZN(G393));
  INV_X1    g0851(.A(new_n944), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n740), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n799), .B1(new_n211), .B2(new_n226), .C1(new_n249), .C2(new_n980), .ZN(new_n1054));
  INV_X1    g0854(.A(G294), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n320), .B1(new_n1055), .B2(new_n759), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n748), .A2(new_n822), .B1(new_n751), .B2(new_n206), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n1056), .A2(new_n784), .A3(new_n1057), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n780), .A2(new_n994), .B1(new_n762), .B2(new_n757), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT52), .ZN(new_n1060));
  INV_X1    g0860(.A(G283), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n770), .A2(new_n1061), .B1(new_n754), .B2(new_n760), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT107), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1058), .A2(new_n1060), .A3(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n751), .A2(new_n202), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n825), .B(new_n413), .C1(new_n834), .C2(new_n754), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(G50), .C2(new_n747), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n780), .A2(new_n342), .B1(new_n762), .B2(new_n777), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT51), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n330), .A2(new_n832), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1067), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n770), .A2(new_n293), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1064), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n742), .B1(new_n1073), .B2(new_n790), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1054), .B(new_n1074), .C1(new_n931), .C2(new_n801), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1053), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n693), .B1(new_n1011), .B2(new_n944), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n734), .A2(new_n1052), .A3(new_n1010), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(G390));
  INV_X1    g0880(.A(new_n814), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1081), .B(new_n892), .C1(new_n729), .C2(new_n730), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n885), .B1(new_n860), .B2(new_n873), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n808), .B(new_n667), .C1(new_n704), .C2(new_n705), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1084), .A2(new_n893), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1083), .B1(new_n1085), .B2(new_n892), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n809), .A2(new_n893), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n885), .B1(new_n1087), .B2(new_n903), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1082), .B(new_n1086), .C1(new_n1088), .C2(new_n884), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n902), .A2(G330), .A3(new_n814), .A4(new_n903), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n880), .B(new_n883), .C1(new_n894), .C2(new_n885), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1092), .B1(new_n1093), .B2(new_n1086), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1081), .B1(new_n729), .B2(new_n730), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1091), .B1(new_n1096), .B2(new_n903), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n1087), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n903), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n727), .A2(KEYINPUT108), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT108), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n725), .A2(new_n726), .A3(new_n1101), .A4(G330), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1100), .A2(new_n814), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n892), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1099), .A2(new_n1104), .A3(new_n1085), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1098), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n443), .A2(G330), .A3(new_n902), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n898), .A2(new_n657), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1095), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n898), .A2(new_n657), .A3(new_n1107), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n1098), .B2(new_n1105), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1086), .B1(new_n1088), .B2(new_n884), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n1091), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n1089), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT109), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1112), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1116), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n692), .B(new_n1110), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n762), .A2(new_n206), .B1(new_n754), .B2(new_n1055), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n785), .B(new_n1120), .C1(G97), .C2(new_n832), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n780), .A2(new_n1061), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1065), .B(new_n1122), .C1(new_n611), .C2(new_n747), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1121), .A2(new_n1123), .A3(new_n320), .A4(new_n827), .ZN(new_n1124));
  XOR2_X1   g0924(.A(new_n1124), .B(KEYINPUT111), .Z(new_n1125));
  OAI21_X1  g0925(.A(new_n264), .B1(new_n215), .B2(new_n765), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT110), .Z(new_n1127));
  OAI21_X1  g0927(.A(KEYINPUT53), .B1(new_n770), .B2(new_n342), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n748), .B2(new_n989), .ZN(new_n1129));
  XOR2_X1   g0929(.A(KEYINPUT54), .B(G143), .Z(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(G125), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n1131), .A2(new_n759), .B1(new_n1132), .B2(new_n754), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n770), .A2(KEYINPUT53), .A3(new_n342), .ZN(new_n1134));
  INV_X1    g0934(.A(G128), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n780), .A2(new_n1135), .B1(new_n751), .B2(new_n777), .ZN(new_n1136));
  NOR4_X1   g0936(.A1(new_n1129), .A2(new_n1133), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1127), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G132), .B2(new_n786), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n790), .B1(new_n1125), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n741), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n884), .A2(new_n797), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(new_n329), .C2(new_n844), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n1115), .B2(new_n740), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1119), .A2(new_n1144), .ZN(G378));
  AND2_X1   g0945(.A1(new_n357), .A2(new_n852), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n374), .B2(new_n379), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT55), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n374), .A2(new_n379), .A3(new_n1147), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n651), .B(new_n1146), .C1(new_n370), .C2(new_n373), .ZN(new_n1153));
  OAI21_X1  g0953(.A(KEYINPUT55), .B1(new_n1148), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT56), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1152), .A2(new_n1154), .A3(KEYINPUT56), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1157), .A2(new_n796), .A3(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n832), .A2(new_n331), .B1(G97), .B2(new_n747), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT112), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1017), .B(new_n273), .C1(new_n206), .C2(new_n780), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1162), .A2(new_n413), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n762), .A2(new_n515), .B1(new_n754), .B2(new_n1061), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n986), .B(new_n1164), .C1(G58), .C2(new_n766), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1161), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT113), .ZN(new_n1167));
  OR2_X1    g0967(.A1(new_n1167), .A2(KEYINPUT58), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n762), .A2(new_n1135), .B1(new_n759), .B2(new_n989), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n771), .B2(new_n1130), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G125), .A2(new_n768), .B1(new_n747), .B2(G132), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(new_n342), .C2(new_n751), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT59), .Z(new_n1173));
  AOI21_X1  g0973(.A(G41), .B1(new_n755), .B2(G124), .ZN(new_n1174));
  AOI21_X1  g0974(.A(G33), .B1(new_n766), .B2(G159), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1167), .A2(KEYINPUT58), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n273), .B1(new_n255), .B2(new_n257), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n215), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1168), .A2(new_n1176), .A3(new_n1177), .A4(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n790), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1181), .B(KEYINPUT114), .Z(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n215), .B2(new_n844), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1159), .A2(new_n741), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n892), .A2(new_n1081), .A3(new_n901), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1187), .A2(new_n906), .B1(new_n904), .B2(KEYINPUT40), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1186), .B1(new_n1188), .B2(new_n743), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n908), .A2(G330), .A3(new_n1158), .A4(new_n1157), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(new_n1190), .A3(KEYINPUT115), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n897), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1191), .B(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1185), .B1(new_n1193), .B2(new_n740), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1108), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT57), .B1(new_n1195), .B2(new_n1193), .ZN(new_n1196));
  OAI21_X1  g0996(.A(KEYINPUT109), .B1(new_n1095), .B2(new_n1109), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1112), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1111), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1189), .A2(new_n1190), .A3(new_n897), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n897), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1202));
  OAI21_X1  g1002(.A(KEYINPUT57), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n692), .B1(new_n1199), .B2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1194), .B1(new_n1196), .B2(new_n1204), .ZN(G375));
  NAND3_X1  g1005(.A1(new_n1111), .A2(new_n1098), .A3(new_n1105), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1109), .A2(new_n955), .A3(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT116), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n770), .A2(new_n211), .B1(new_n754), .B2(new_n822), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n983), .B(new_n1209), .C1(new_n611), .C2(new_n832), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n768), .A2(G294), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1015), .B1(new_n747), .B2(G116), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n264), .B1(G283), .B2(new_n786), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G159), .A2(new_n771), .B1(new_n755), .B2(G128), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(new_n390), .B2(new_n765), .C1(new_n342), .C2(new_n759), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n401), .B(new_n1216), .C1(G50), .C2(new_n830), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT118), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1130), .A2(new_n747), .B1(G132), .B2(new_n768), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n762), .A2(new_n989), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1214), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1224), .A2(new_n790), .B1(new_n293), .B2(new_n844), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n741), .B(new_n1225), .C1(new_n903), .C2(new_n797), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n740), .B(KEYINPUT117), .Z(new_n1228));
  AOI21_X1  g1028(.A(new_n1227), .B1(new_n1106), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1208), .A2(new_n1229), .ZN(G381));
  INV_X1    g1030(.A(new_n1203), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n693), .B1(new_n1195), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT57), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1191), .B(new_n897), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1233), .B1(new_n1199), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(G378), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(new_n1237), .A3(new_n1194), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1238), .A2(G384), .A3(G381), .ZN(new_n1239));
  INV_X1    g1039(.A(G396), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1013), .A2(new_n1050), .A3(new_n1240), .A4(new_n1014), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(G387), .A2(G390), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1239), .A2(new_n1242), .ZN(G407));
  NAND2_X1  g1043(.A1(new_n665), .A2(G213), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n1244), .B(KEYINPUT119), .Z(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  OAI211_X1 g1046(.A(G407), .B(G213), .C1(new_n1238), .C2(new_n1246), .ZN(G409));
  INV_X1    g1047(.A(KEYINPUT125), .ZN(new_n1248));
  AOI21_X1  g1048(.A(G390), .B1(new_n977), .B2(new_n1008), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1008), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1250), .B(new_n1079), .C1(new_n958), .C2(new_n976), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1248), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G393), .A2(G396), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT124), .ZN(new_n1254));
  AND3_X1   g1054(.A1(new_n1253), .A2(new_n1254), .A3(new_n1241), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1254), .B1(new_n1253), .B2(new_n1241), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1252), .A2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1257), .B(new_n1248), .C1(new_n1251), .C2(new_n1249), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1245), .A2(G2897), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT60), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n693), .B1(new_n1206), .B2(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1111), .A2(new_n1098), .A3(KEYINPUT60), .A4(new_n1105), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1266), .A2(KEYINPUT120), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1266), .A2(KEYINPUT120), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1109), .B(new_n1265), .C1(new_n1267), .C2(new_n1268), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1269), .A2(new_n849), .A3(new_n1229), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n849), .B1(new_n1269), .B2(new_n1229), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1263), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(KEYINPUT121), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT120), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1266), .B(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1265), .A2(new_n1109), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1229), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(G384), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1269), .A2(new_n849), .A3(new_n1229), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT121), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1280), .A2(new_n1281), .A3(new_n1263), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1263), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1278), .A2(new_n1279), .A3(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT122), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1278), .A2(KEYINPUT122), .A3(new_n1279), .A4(new_n1283), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1273), .A2(new_n1282), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT126), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1237), .B1(new_n1236), .B2(new_n1194), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1195), .A2(new_n955), .A3(new_n1193), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1228), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1119), .A2(new_n1144), .A3(new_n1184), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1246), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1289), .B1(new_n1290), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G375), .A2(G378), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1292), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1234), .B1(new_n1299), .B2(new_n1108), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1298), .B1(new_n1300), .B2(new_n955), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1119), .A2(new_n1144), .A3(new_n1184), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1245), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1297), .A2(KEYINPUT126), .A3(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1288), .A2(new_n1296), .A3(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT61), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT62), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1297), .A2(new_n1303), .A3(new_n1307), .A4(new_n1280), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1305), .A2(new_n1306), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1296), .A2(new_n1304), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1307), .B1(new_n1310), .B2(new_n1280), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1262), .B1(new_n1309), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1297), .A2(new_n1303), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1273), .A2(new_n1282), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1314), .A2(KEYINPUT123), .A3(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(KEYINPUT123), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1313), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1297), .A2(new_n1280), .A3(new_n1303), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT63), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1321), .A2(new_n1306), .A3(new_n1261), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1310), .A2(KEYINPUT63), .A3(new_n1280), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1318), .A2(new_n1322), .A3(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1312), .A2(new_n1324), .ZN(G405));
  INV_X1    g1125(.A(new_n1238), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1280), .B1(new_n1326), .B2(new_n1290), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1297), .A2(new_n1238), .A3(new_n1279), .A4(new_n1278), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(KEYINPUT127), .B1(new_n1329), .B2(new_n1262), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1262), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT127), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1327), .A2(new_n1261), .A3(new_n1332), .A4(new_n1328), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1330), .A2(new_n1331), .A3(new_n1333), .ZN(G402));
endmodule


