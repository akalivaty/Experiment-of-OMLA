//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1222, new_n1223, new_n1224;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  OR4_X1    g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  NAND2_X1  g032(.A1(G113), .A2(G2104), .ZN(new_n458));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n465), .C1(new_n459), .C2(new_n460), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n466), .A2(KEYINPUT67), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(KEYINPUT67), .B1(new_n466), .B2(new_n469), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT68), .ZN(G160));
  NOR2_X1   g048(.A1(new_n461), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n461), .A2(new_n465), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(new_n465), .B2(G112), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n475), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT69), .ZN(G162));
  INV_X1    g056(.A(new_n468), .ZN(new_n482));
  INV_X1    g057(.A(G102), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(G114), .A2(G2104), .ZN(new_n485));
  INV_X1    g060(.A(G126), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n485), .B1(new_n461), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n484), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(G138), .B(new_n465), .C1(new_n459), .C2(new_n460), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  XNOR2_X1  g065(.A(KEYINPUT3), .B(G2104), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n491), .A2(new_n492), .A3(G138), .A4(new_n465), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  NAND2_X1  g071(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n497));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n501), .A2(G62), .ZN(new_n502));
  NAND2_X1  g077(.A1(G75), .A2(G543), .ZN(new_n503));
  XOR2_X1   g078(.A(new_n503), .B(KEYINPUT73), .Z(new_n504));
  OAI21_X1  g079(.A(G651), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(KEYINPUT6), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT70), .A3(G651), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n508), .A2(new_n510), .B1(KEYINPUT6), .B2(new_n507), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(G88), .A3(new_n501), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(new_n510), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n513), .A2(G50), .A3(G543), .A4(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n516));
  AND3_X1   g091(.A1(new_n512), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n516), .B1(new_n512), .B2(new_n515), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n505), .B1(new_n517), .B2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND3_X1  g095(.A1(new_n511), .A2(G51), .A3(G543), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n511), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n524));
  AND3_X1   g099(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n525));
  AOI21_X1  g100(.A(G543), .B1(KEYINPUT71), .B2(KEYINPUT5), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n521), .B(new_n523), .C1(new_n524), .C2(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  NAND3_X1  g104(.A1(new_n511), .A2(G90), .A3(new_n501), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n511), .A2(G52), .A3(G543), .ZN(new_n531));
  INV_X1    g106(.A(G64), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n532), .B1(new_n499), .B2(new_n500), .ZN(new_n533));
  AND2_X1   g108(.A1(G77), .A2(G543), .ZN(new_n534));
  OAI21_X1  g109(.A(G651), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n530), .A2(new_n531), .A3(new_n535), .ZN(G171));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n537));
  INV_X1    g112(.A(G56), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n538), .B1(new_n499), .B2(new_n500), .ZN(new_n539));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n537), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g117(.A(G56), .B1(new_n525), .B2(new_n526), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n543), .A2(KEYINPUT74), .A3(new_n540), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n542), .A2(G651), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n511), .A2(G43), .A3(G543), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n511), .A2(G81), .A3(new_n501), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  NAND3_X1  g130(.A1(new_n513), .A2(new_n501), .A3(new_n514), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n527), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n557), .A2(G91), .B1(new_n560), .B2(G651), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n513), .A2(G53), .A3(G543), .A4(new_n514), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n511), .A2(new_n564), .A3(G53), .A4(G543), .ZN(new_n565));
  AND3_X1   g140(.A1(new_n563), .A2(KEYINPUT75), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g141(.A(KEYINPUT75), .B1(new_n563), .B2(new_n565), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n561), .B1(new_n566), .B2(new_n567), .ZN(G299));
  NAND3_X1  g143(.A1(new_n530), .A2(new_n531), .A3(new_n535), .ZN(G301));
  NAND3_X1  g144(.A1(new_n511), .A2(G49), .A3(G543), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n511), .A2(G87), .A3(new_n501), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n513), .A2(G543), .A3(new_n514), .ZN(new_n575));
  INV_X1    g150(.A(G48), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n511), .A2(KEYINPUT76), .A3(G48), .A4(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n557), .A2(G86), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n501), .A2(G61), .ZN(new_n581));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n507), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n579), .A2(new_n580), .A3(new_n584), .ZN(G305));
  AOI22_X1  g160(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n586), .A2(new_n507), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n511), .A2(G85), .A3(new_n501), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n513), .A2(G47), .A3(G543), .A4(new_n514), .ZN(new_n589));
  AND3_X1   g164(.A1(new_n588), .A2(new_n589), .A3(KEYINPUT77), .ZN(new_n590));
  AOI21_X1  g165(.A(KEYINPUT77), .B1(new_n588), .B2(new_n589), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n587), .B1(new_n590), .B2(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  XOR2_X1   g168(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G92), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n556), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n527), .A2(new_n598), .ZN(new_n599));
  AND2_X1   g174(.A1(G79), .A2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n511), .A2(G92), .A3(new_n501), .A4(new_n594), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n511), .A2(G54), .A3(G543), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n597), .A2(new_n601), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n593), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n593), .B1(new_n605), .B2(G868), .ZN(G321));
  NAND2_X1  g182(.A1(G286), .A2(G868), .ZN(new_n608));
  INV_X1    g183(.A(G299), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(G297));
  OAI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n605), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n491), .A2(new_n468), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT79), .B(G2100), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n619), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n474), .A2(G135), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n623), .A2(KEYINPUT80), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n623), .A2(KEYINPUT80), .B1(G123), .B2(new_n476), .ZN(new_n625));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n626), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n627));
  AND3_X1   g202(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT81), .ZN(new_n629));
  AND2_X1   g204(.A1(new_n629), .A2(G2096), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n629), .A2(G2096), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n622), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT82), .ZN(G156));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2435), .ZN(new_n641));
  XOR2_X1   g216(.A(G2427), .B(G2438), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n639), .B(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(G14), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n645), .A2(new_n646), .ZN(G401));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  XNOR2_X1  g223(.A(G2072), .B(G2078), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT83), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n648), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n649), .B(KEYINPUT17), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n653), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT84), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n648), .A2(new_n651), .A3(new_n649), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT18), .Z(new_n660));
  NAND3_X1  g235(.A1(new_n655), .A2(new_n648), .A3(new_n652), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2096), .ZN(new_n663));
  INV_X1    g238(.A(G2100), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n662), .A2(G2096), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n662), .A2(G2096), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(G2100), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n668), .ZN(G227));
  INV_X1    g244(.A(KEYINPUT20), .ZN(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT85), .ZN(new_n672));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n670), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n672), .A2(new_n673), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n678), .A2(new_n676), .A3(new_n674), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n672), .A2(KEYINPUT20), .A3(new_n673), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n677), .B(new_n679), .C1(new_n681), .C2(new_n676), .ZN(new_n682));
  XOR2_X1   g257(.A(G1991), .B(G1996), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1981), .B(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G229));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G4), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(new_n605), .B2(new_n689), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT90), .B(G1348), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n468), .A2(G103), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT25), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n474), .A2(G139), .ZN(new_n697));
  AOI22_X1  g272(.A1(new_n491), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n696), .B(new_n697), .C1(new_n465), .C2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT91), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G29), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G29), .B2(G33), .ZN(new_n705));
  INV_X1    g280(.A(G2072), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT92), .Z(new_n708));
  NOR2_X1   g283(.A1(G29), .A2(G35), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G162), .B2(G29), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G2090), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n705), .A2(new_n706), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G27), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G164), .B2(new_n714), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT95), .B(G2078), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(G26), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n474), .A2(G140), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n476), .A2(G128), .ZN(new_n721));
  OR2_X1    g296(.A1(G104), .A2(G2105), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n722), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n720), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n719), .B1(new_n725), .B2(new_n714), .ZN(new_n726));
  MUX2_X1   g301(.A(new_n719), .B(new_n726), .S(KEYINPUT28), .Z(new_n727));
  NOR2_X1   g302(.A1(G16), .A2(G21), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G168), .B2(G16), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n727), .A2(G2067), .B1(G1966), .B2(new_n729), .ZN(new_n730));
  AND4_X1   g305(.A1(new_n712), .A2(new_n713), .A3(new_n718), .A4(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n711), .A2(G2090), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n727), .A2(G2067), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n708), .A2(new_n731), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n689), .A2(G20), .ZN(new_n735));
  OAI211_X1 g310(.A(KEYINPUT23), .B(new_n735), .C1(new_n609), .C2(new_n689), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(KEYINPUT23), .B2(new_n735), .ZN(new_n737));
  INV_X1    g312(.A(G1956), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G5), .A2(G16), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G171), .B2(G16), .ZN(new_n741));
  OAI22_X1  g316(.A1(new_n729), .A2(G1966), .B1(new_n741), .B2(G1961), .ZN(new_n742));
  OR2_X1    g317(.A1(G29), .A2(G32), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n474), .A2(G141), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n476), .A2(G129), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT26), .Z(new_n747));
  NAND3_X1  g322(.A1(new_n744), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n468), .A2(G105), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT94), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n743), .B1(new_n752), .B2(new_n714), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT27), .B(G1996), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n714), .B1(new_n757), .B2(G28), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n757), .B2(G28), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n628), .B2(G29), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n755), .A2(new_n756), .A3(new_n760), .ZN(new_n761));
  AOI211_X1 g336(.A(new_n742), .B(new_n761), .C1(G1961), .C2(new_n741), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT31), .B(G11), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT93), .B(G34), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT24), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n765), .A2(G29), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G160), .B2(G29), .ZN(new_n767));
  INV_X1    g342(.A(G2084), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n689), .A2(G19), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n549), .B2(new_n689), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(G1341), .Z(new_n772));
  NAND4_X1  g347(.A1(new_n762), .A2(new_n763), .A3(new_n769), .A4(new_n772), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n734), .A2(new_n739), .A3(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G24), .ZN(new_n775));
  OAI21_X1  g350(.A(KEYINPUT87), .B1(new_n775), .B2(G16), .ZN(new_n776));
  OR3_X1    g351(.A1(new_n775), .A2(KEYINPUT87), .A3(G16), .ZN(new_n777));
  INV_X1    g352(.A(G290), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n776), .B(new_n777), .C1(new_n778), .C2(new_n689), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(G1986), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(G1986), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n714), .A2(G25), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n474), .A2(G131), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n476), .A2(G119), .ZN(new_n784));
  OR2_X1    g359(.A1(G95), .A2(G2105), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n785), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n783), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n782), .B1(new_n788), .B2(new_n714), .ZN(new_n789));
  MUX2_X1   g364(.A(new_n782), .B(new_n789), .S(KEYINPUT86), .Z(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT35), .B(G1991), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n780), .A2(new_n781), .A3(new_n792), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n689), .A2(G6), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G305), .B2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT32), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1981), .ZN(new_n797));
  OAI21_X1  g372(.A(KEYINPUT88), .B1(G16), .B2(G23), .ZN(new_n798));
  OR3_X1    g373(.A1(KEYINPUT88), .A2(G16), .A3(G23), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n798), .B(new_n799), .C1(G288), .C2(new_n689), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT33), .B(G1976), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n689), .A2(G22), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G166), .B2(new_n689), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT89), .B(G1971), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n797), .A2(new_n802), .A3(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT34), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n797), .A2(KEYINPUT34), .A3(new_n802), .A4(new_n806), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n793), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n790), .A2(new_n791), .ZN(new_n813));
  AND3_X1   g388(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n812), .B1(new_n811), .B2(new_n813), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n693), .B(new_n774), .C1(new_n814), .C2(new_n815), .ZN(G150));
  NAND2_X1  g391(.A1(G150), .A2(KEYINPUT96), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n809), .A2(new_n810), .ZN(new_n818));
  INV_X1    g393(.A(new_n793), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n818), .A2(new_n813), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT36), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT96), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n823), .A2(new_n824), .A3(new_n693), .A4(new_n774), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n817), .A2(new_n825), .ZN(G311));
  INV_X1    g401(.A(KEYINPUT97), .ZN(new_n827));
  INV_X1    g402(.A(G67), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n499), .B2(new_n500), .ZN(new_n829));
  NAND2_X1  g404(.A1(G80), .A2(G543), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n827), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  OAI211_X1 g407(.A(KEYINPUT97), .B(new_n830), .C1(new_n527), .C2(new_n828), .ZN(new_n833));
  AND3_X1   g408(.A1(new_n832), .A2(new_n833), .A3(G651), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n511), .A2(G55), .A3(G543), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n511), .A2(G93), .A3(new_n501), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(G860), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  INV_X1    g414(.A(new_n548), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n542), .A2(G651), .A3(new_n544), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n840), .B(new_n841), .C1(new_n834), .C2(new_n837), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n836), .A2(new_n835), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n832), .A2(new_n833), .A3(G651), .ZN(new_n844));
  OAI211_X1 g419(.A(new_n843), .B(new_n844), .C1(new_n545), .C2(new_n548), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT39), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n605), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n847), .B(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n839), .B1(new_n850), .B2(G860), .ZN(G145));
  NAND2_X1  g426(.A1(new_n701), .A2(new_n702), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(new_n725), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n724), .B1(new_n701), .B2(new_n702), .ZN(new_n854));
  OAI21_X1  g429(.A(G164), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n853), .A2(G164), .A3(new_n854), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n752), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n474), .A2(G142), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n476), .A2(G130), .ZN(new_n860));
  NOR2_X1   g435(.A1(G106), .A2(G2105), .ZN(new_n861));
  OAI21_X1  g436(.A(G2104), .B1(new_n465), .B2(G118), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n859), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(new_n619), .Z(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(new_n787), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n787), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(KEYINPUT98), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT98), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n853), .ZN(new_n871));
  INV_X1    g446(.A(new_n854), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(new_n872), .A3(new_n495), .ZN(new_n873));
  INV_X1    g448(.A(new_n752), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n873), .A2(new_n855), .A3(new_n874), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n858), .A2(new_n867), .A3(new_n870), .A4(new_n875), .ZN(new_n876));
  XOR2_X1   g451(.A(G160), .B(new_n628), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G162), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n880));
  INV_X1    g455(.A(new_n875), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n874), .B1(new_n873), .B2(new_n855), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n858), .A2(KEYINPUT99), .A3(new_n875), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n876), .B(new_n879), .C1(new_n885), .C2(new_n868), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n870), .A2(new_n867), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(new_n881), .B2(new_n882), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n876), .ZN(new_n889));
  AOI21_X1  g464(.A(G37), .B1(new_n889), .B2(new_n878), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT40), .ZN(G395));
  NOR3_X1   g467(.A1(new_n834), .A2(G868), .A3(new_n837), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT101), .ZN(new_n894));
  XOR2_X1   g469(.A(G290), .B(KEYINPUT100), .Z(new_n895));
  INV_X1    g470(.A(G288), .ZN(new_n896));
  NAND2_X1  g471(.A1(G303), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n505), .B(G288), .C1(new_n517), .C2(new_n518), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G305), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n898), .A3(G305), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n895), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(G290), .B(KEYINPUT100), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n897), .A2(new_n898), .A3(G305), .ZN(new_n905));
  AOI21_X1  g480(.A(G305), .B1(new_n897), .B2(new_n898), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT42), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n846), .B(new_n614), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n563), .A2(new_n565), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT75), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n563), .A2(KEYINPUT75), .A3(new_n565), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n604), .B1(new_n915), .B2(new_n561), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n604), .B(new_n561), .C1(new_n566), .C2(new_n567), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n910), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT41), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(new_n916), .B2(new_n918), .ZN(new_n922));
  NAND2_X1  g497(.A1(G299), .A2(new_n605), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n923), .A2(KEYINPUT41), .A3(new_n917), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n920), .B1(new_n925), .B2(new_n910), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n894), .B1(new_n909), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n909), .A2(new_n926), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n927), .B(new_n928), .Z(new_n929));
  AOI21_X1  g504(.A(new_n893), .B1(new_n929), .B2(G868), .ZN(G295));
  AOI21_X1  g505(.A(new_n893), .B1(new_n929), .B2(G868), .ZN(G331));
  NAND2_X1  g506(.A1(new_n511), .A2(G89), .ZN(new_n932));
  NAND2_X1  g507(.A1(G63), .A2(G651), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n501), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n935), .A2(G301), .A3(new_n521), .A4(new_n523), .ZN(new_n936));
  NAND2_X1  g511(.A1(G286), .A2(G171), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n846), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n842), .A2(new_n845), .A3(new_n936), .A4(new_n937), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(KEYINPUT102), .A3(new_n940), .ZN(new_n941));
  OR3_X1    g516(.A1(new_n846), .A2(new_n938), .A3(KEYINPUT102), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n923), .A2(KEYINPUT41), .A3(new_n917), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT41), .B1(new_n923), .B2(new_n917), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n941), .B(new_n942), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT103), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n939), .A2(new_n940), .ZN(new_n948));
  OR2_X1    g523(.A1(new_n948), .A2(new_n919), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n925), .A2(KEYINPUT103), .A3(new_n942), .A4(new_n941), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n947), .A2(new_n908), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n952));
  INV_X1    g527(.A(G37), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n903), .A2(new_n907), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n922), .A2(new_n924), .B1(new_n940), .B2(new_n939), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n919), .B1(new_n941), .B2(new_n942), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT104), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n956), .A2(new_n955), .ZN(new_n961));
  AOI21_X1  g536(.A(G37), .B1(new_n961), .B2(new_n954), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n962), .A2(KEYINPUT104), .A3(new_n952), .A4(new_n951), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n954), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n966), .A2(new_n953), .A3(new_n951), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT44), .B1(new_n964), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n967), .A2(new_n952), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n962), .A2(KEYINPUT43), .A3(new_n951), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT105), .B1(new_n969), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n968), .A2(new_n960), .A3(new_n963), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n970), .ZN(new_n976));
  INV_X1    g551(.A(new_n973), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n974), .A2(new_n979), .ZN(G397));
  INV_X1    g555(.A(G1986), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n778), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT108), .ZN(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n491), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n985));
  OAI22_X1  g560(.A1(new_n985), .A2(new_n465), .B1(new_n483), .B2(new_n482), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n490), .A2(new_n493), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  XOR2_X1   g566(.A(KEYINPUT107), .B(G40), .Z(new_n992));
  OAI211_X1 g567(.A(new_n464), .B(new_n992), .C1(new_n470), .C2(new_n471), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n778), .A2(new_n981), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n983), .B(new_n994), .C1(new_n997), .C2(new_n982), .ZN(new_n998));
  INV_X1    g573(.A(G1996), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n874), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G2067), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n724), .B(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n752), .A2(G1996), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1000), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n787), .B(new_n791), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n994), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n998), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT49), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n583), .B1(new_n577), .B2(new_n578), .ZN(new_n1009));
  INV_X1    g584(.A(G1981), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n1009), .A2(new_n1010), .A3(new_n580), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n1009), .B2(new_n580), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1008), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(G305), .A2(G1981), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1009), .A2(new_n1010), .A3(new_n580), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(KEYINPUT49), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n988), .A2(new_n993), .ZN(new_n1017));
  INV_X1    g592(.A(G8), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1013), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1013), .A2(new_n1016), .A3(KEYINPUT113), .A4(new_n1019), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n993), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1384), .B1(new_n488), .B2(new_n494), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n896), .A2(KEYINPUT111), .A3(G1976), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n1029));
  INV_X1    g604(.A(G1976), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(G288), .B2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1027), .A2(new_n1028), .A3(G8), .A4(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n896), .A2(G1976), .ZN(new_n1033));
  OR3_X1    g608(.A1(new_n1032), .A2(KEYINPUT52), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(KEYINPUT52), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT112), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1032), .A2(KEYINPUT112), .A3(KEYINPUT52), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1024), .A2(new_n1034), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1022), .A2(new_n1023), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(KEYINPUT118), .A3(new_n1034), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G303), .A2(G8), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1046), .B(KEYINPUT55), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1026), .A2(KEYINPUT50), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT50), .ZN(new_n1050));
  AOI211_X1 g625(.A(new_n1050), .B(G1384), .C1(new_n488), .C2(new_n494), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1025), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G2090), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n495), .A2(KEYINPUT45), .A3(new_n984), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT110), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1026), .A2(KEYINPUT110), .A3(KEYINPUT45), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n993), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n988), .A2(KEYINPUT109), .A3(new_n990), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT109), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n1026), .B2(new_n989), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(G1971), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1048), .B(G8), .C1(new_n1056), .C2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1052), .A2(KEYINPUT116), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1071), .B(new_n1025), .C1(new_n1049), .C2(new_n1051), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1070), .A2(new_n1054), .A3(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1069), .B1(new_n1073), .B2(new_n1066), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1066), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1070), .A2(new_n1054), .A3(new_n1072), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(new_n1076), .A3(KEYINPUT117), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(G8), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1068), .B1(new_n1078), .B2(new_n1047), .ZN(new_n1079));
  INV_X1    g654(.A(G1966), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1025), .B1(new_n988), .B2(new_n990), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1026), .A2(KEYINPUT45), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n768), .B(new_n1025), .C1(new_n1049), .C2(new_n1051), .ZN(new_n1084));
  AOI211_X1 g659(.A(new_n1018), .B(G286), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1045), .A2(new_n1079), .A3(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT119), .B(KEYINPUT63), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1089), .A2(new_n1065), .A3(new_n1025), .ZN(new_n1090));
  INV_X1    g665(.A(G1971), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1090), .A2(new_n1091), .B1(new_n1054), .B2(new_n1053), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1047), .B1(new_n1092), .B2(new_n1018), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1043), .A2(new_n1093), .A3(new_n1034), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1067), .A2(KEYINPUT63), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1094), .A2(KEYINPUT120), .A3(new_n1096), .A4(new_n1085), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1043), .A2(new_n1093), .A3(new_n1034), .A4(new_n1085), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1098), .B1(new_n1099), .B2(new_n1095), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1088), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G2078), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1089), .A2(new_n1065), .A3(new_n1103), .A4(new_n1025), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n1105));
  INV_X1    g680(.A(G1961), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1104), .A2(new_n1105), .B1(new_n1106), .B2(new_n1052), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1105), .A2(G2078), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(G171), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1083), .A2(G168), .A3(new_n1084), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(G8), .A3(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1120), .A2(G8), .A3(G286), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1118), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1113), .A2(G8), .A3(new_n1116), .A4(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1119), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1112), .B1(new_n1124), .B2(KEYINPUT62), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT62), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1119), .A2(new_n1126), .A3(new_n1121), .A4(new_n1123), .ZN(new_n1127));
  AND4_X1   g702(.A1(new_n1045), .A2(new_n1079), .A3(new_n1125), .A4(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(G288), .A2(G1976), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1024), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(KEYINPUT115), .A3(new_n1015), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT115), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1129), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1133), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1132), .B1(new_n1134), .B2(new_n1011), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1019), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1136), .A2(KEYINPUT114), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(KEYINPUT114), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1131), .A2(new_n1135), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(new_n1040), .B2(new_n1067), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1128), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1102), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1052), .A2(new_n1106), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1143), .A2(G301), .A3(new_n1144), .A4(new_n1110), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT124), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n472), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1147), .A2(G40), .A3(new_n991), .A4(new_n1109), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1143), .A2(new_n1144), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(G171), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1107), .A2(new_n1151), .A3(G301), .A4(new_n1110), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1146), .A2(new_n1150), .A3(KEYINPUT54), .A4(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT54), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1107), .A2(G301), .A3(new_n1148), .ZN(new_n1155));
  AOI21_X1  g730(.A(G301), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1158), .A2(new_n1124), .A3(new_n1045), .A4(new_n1079), .ZN(new_n1159));
  XNOR2_X1  g734(.A(KEYINPUT56), .B(G2072), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1061), .A2(new_n1065), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1052), .A2(new_n738), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT57), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n561), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n911), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1167), .B1(KEYINPUT57), .B2(G299), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1163), .A2(new_n1169), .ZN(new_n1170));
  OAI22_X1  g745(.A1(new_n1053), .A2(G1348), .B1(G2067), .B2(new_n1027), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1170), .B1(new_n604), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1161), .A2(new_n1168), .A3(new_n1162), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(KEYINPUT121), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1161), .A2(new_n1176), .A3(new_n1168), .A4(new_n1162), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1173), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1175), .A2(new_n1170), .A3(new_n1177), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1170), .A2(KEYINPUT61), .A3(new_n1174), .ZN(new_n1182));
  XNOR2_X1  g757(.A(KEYINPUT58), .B(G1341), .ZN(new_n1183));
  OAI22_X1  g758(.A1(new_n1090), .A2(G1996), .B1(new_n1017), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT59), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1184), .A2(new_n1185), .A3(new_n549), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1185), .B1(new_n1184), .B2(new_n549), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1182), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(KEYINPUT122), .B1(new_n1181), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1172), .A2(KEYINPUT60), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(new_n605), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1191), .B1(KEYINPUT60), .B2(new_n1172), .ZN(new_n1192));
  OR2_X1    g767(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT122), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .A4(new_n1182), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1189), .A2(new_n1192), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1159), .B1(new_n1178), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1007), .B1(new_n1142), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(new_n994), .ZN(new_n1200));
  OR3_X1    g775(.A1(new_n1004), .A2(new_n791), .A3(new_n787), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n725), .A2(new_n1001), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1200), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n994), .A2(new_n999), .ZN(new_n1204));
  XOR2_X1   g779(.A(new_n1204), .B(KEYINPUT46), .Z(new_n1205));
  NAND2_X1  g780(.A1(new_n1002), .A2(new_n874), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1206), .A2(new_n994), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1207), .B(KEYINPUT125), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(KEYINPUT47), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1200), .A2(new_n995), .ZN(new_n1211));
  XOR2_X1   g786(.A(new_n1211), .B(KEYINPUT48), .Z(new_n1212));
  AOI211_X1 g787(.A(new_n1203), .B(new_n1210), .C1(new_n1006), .C2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1199), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g789(.A(G229), .B1(new_n886), .B2(new_n890), .ZN(new_n1216));
  NAND3_X1  g790(.A1(new_n665), .A2(G319), .A3(new_n668), .ZN(new_n1217));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n1218));
  OAI22_X1  g792(.A1(new_n1217), .A2(new_n1218), .B1(new_n646), .B2(new_n645), .ZN(new_n1219));
  AOI21_X1  g793(.A(new_n1219), .B1(new_n1218), .B2(new_n1217), .ZN(new_n1220));
  NAND3_X1  g794(.A1(new_n1216), .A2(new_n975), .A3(new_n1220), .ZN(G225));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n1222));
  NAND2_X1  g796(.A1(G225), .A2(new_n1222), .ZN(new_n1223));
  NAND4_X1  g797(.A1(new_n1216), .A2(new_n975), .A3(new_n1220), .A4(KEYINPUT127), .ZN(new_n1224));
  NAND2_X1  g798(.A1(new_n1223), .A2(new_n1224), .ZN(G308));
endmodule


