//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 0 0 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT0), .A2(G128), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n188), .A2(new_n190), .A3(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G143), .B(G146), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT0), .B(G128), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n192), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G137), .ZN(new_n198));
  INV_X1    g012(.A(G137), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT11), .A3(G134), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(G137), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n198), .A2(new_n200), .A3(new_n201), .A4(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n198), .A2(new_n200), .A3(new_n202), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G131), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n195), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n189), .A2(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n187), .A2(G143), .ZN(new_n209));
  OAI211_X1 g023(.A(G128), .B(new_n207), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n197), .A2(G137), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n199), .A2(G134), .ZN(new_n212));
  OAI21_X1  g026(.A(G131), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n188), .B(new_n190), .C1(KEYINPUT1), .C2(new_n214), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n210), .A2(new_n203), .A3(new_n213), .A4(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n206), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT64), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT2), .ZN(new_n220));
  INV_X1    g034(.A(G113), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT64), .B1(KEYINPUT2), .B2(G113), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT2), .A2(G113), .ZN(new_n225));
  XNOR2_X1  g039(.A(G116), .B(G119), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n226), .B1(new_n224), .B2(new_n225), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT28), .B1(new_n218), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n205), .A2(new_n203), .ZN(new_n232));
  INV_X1    g046(.A(new_n195), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n234), .A2(new_n229), .A3(new_n216), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n229), .B1(new_n234), .B2(new_n216), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT28), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n231), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(G237), .A2(G953), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G210), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n240), .B(KEYINPUT27), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT26), .B(G101), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n238), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n234), .A2(new_n229), .A3(new_n216), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT65), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n247), .A2(new_n248), .A3(new_n243), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT30), .B1(new_n206), .B2(new_n217), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT30), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n234), .A2(new_n251), .A3(new_n216), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n229), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n248), .B1(new_n247), .B2(new_n243), .ZN(new_n254));
  NOR3_X1   g068(.A1(new_n249), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT66), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT31), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n250), .A2(new_n252), .ZN(new_n258));
  INV_X1    g072(.A(new_n228), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n247), .A2(new_n243), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT65), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n247), .A2(new_n243), .A3(new_n248), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n262), .A2(new_n264), .A3(new_n256), .A4(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT31), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n246), .B1(new_n257), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT32), .ZN(new_n270));
  NOR2_X1   g084(.A1(G472), .A2(G902), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n266), .A2(new_n267), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n249), .A2(new_n253), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n274), .A2(new_n256), .A3(KEYINPUT31), .A4(new_n264), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n273), .A2(new_n275), .B1(new_n238), .B2(new_n245), .ZN(new_n276));
  INV_X1    g090(.A(new_n271), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT32), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n261), .B1(new_n206), .B2(new_n217), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n279), .B1(new_n280), .B2(new_n247), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT68), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n230), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n237), .A2(KEYINPUT68), .ZN(new_n284));
  INV_X1    g098(.A(new_n243), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT29), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n283), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT69), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n288), .A2(KEYINPUT69), .A3(new_n289), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n285), .B1(new_n253), .B2(new_n235), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n294), .B(new_n286), .C1(new_n238), .C2(new_n245), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n292), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n272), .A2(new_n278), .B1(new_n296), .B2(G472), .ZN(new_n297));
  INV_X1    g111(.A(G110), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT24), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT24), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G110), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT70), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n302), .B1(new_n299), .B2(new_n301), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n214), .A2(G119), .ZN(new_n305));
  INV_X1    g119(.A(G119), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(G128), .ZN(new_n307));
  OAI22_X1  g121(.A1(new_n303), .A2(new_n304), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n306), .A2(G128), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n214), .A2(KEYINPUT23), .A3(G119), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n310), .B(new_n311), .C1(new_n307), .C2(KEYINPUT23), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n309), .B1(new_n312), .B2(G110), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT23), .B1(new_n214), .B2(G119), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(new_n305), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n315), .A2(KEYINPUT73), .A3(new_n298), .A4(new_n311), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n308), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(G125), .B(G140), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n187), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n321), .A2(KEYINPUT16), .A3(G140), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n322), .B1(new_n318), .B2(KEYINPUT16), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n320), .B1(new_n323), .B2(G146), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n317), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n303), .A2(new_n304), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n305), .A2(new_n307), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n312), .A2(KEYINPUT71), .A3(G110), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT71), .B1(new_n312), .B2(G110), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G140), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G125), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n321), .A2(G140), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT16), .ZN(new_n335));
  OR3_X1    g149(.A1(new_n321), .A2(KEYINPUT16), .A3(G140), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT72), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n335), .A2(new_n336), .A3(new_n337), .A4(G146), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(new_n323), .B2(G146), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n337), .B1(new_n323), .B2(G146), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n325), .B1(new_n331), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT22), .B(G137), .ZN(new_n343));
  INV_X1    g157(.A(G953), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(G221), .A3(G234), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n343), .B(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n325), .B(new_n346), .C1(new_n341), .C2(new_n331), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n289), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT25), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n348), .A2(KEYINPUT25), .A3(new_n289), .A4(new_n349), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n352), .A2(KEYINPUT74), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT74), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n350), .A2(new_n355), .A3(new_n351), .ZN(new_n356));
  INV_X1    g170(.A(G217), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(G234), .B2(new_n289), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n348), .A2(new_n349), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n358), .A2(G902), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  OAI22_X1  g176(.A1(new_n354), .A2(new_n359), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n297), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(G210), .B1(G237), .B2(G902), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n195), .A2(G125), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n210), .A2(new_n215), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n367), .B1(new_n368), .B2(G125), .ZN(new_n369));
  INV_X1    g183(.A(G224), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(G953), .ZN(new_n371));
  XOR2_X1   g185(.A(new_n369), .B(new_n371), .Z(new_n372));
  NAND2_X1  g186(.A1(new_n226), .A2(KEYINPUT5), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n306), .A2(G116), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n373), .B(G113), .C1(KEYINPUT5), .C2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G104), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT3), .B1(new_n376), .B2(G107), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT3), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(G104), .ZN(new_n380));
  INV_X1    g194(.A(G101), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n376), .A2(G107), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n377), .A2(new_n380), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n376), .A2(G107), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n379), .A2(G104), .ZN(new_n385));
  OAI21_X1  g199(.A(G101), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n375), .A2(new_n387), .A3(new_n260), .ZN(new_n388));
  XNOR2_X1  g202(.A(G110), .B(G122), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n377), .A2(new_n380), .A3(new_n382), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G101), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT75), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(KEYINPUT75), .A3(G101), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n393), .A2(KEYINPUT4), .A3(new_n383), .A4(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  XOR2_X1   g210(.A(KEYINPUT76), .B(KEYINPUT4), .Z(new_n397));
  NAND3_X1  g211(.A1(new_n390), .A2(G101), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n261), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n388), .B(new_n389), .C1(new_n396), .C2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT6), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n388), .B1(new_n396), .B2(new_n399), .ZN(new_n402));
  INV_X1    g216(.A(new_n389), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n403), .A2(KEYINPUT77), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n402), .A2(KEYINPUT6), .A3(new_n404), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n372), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT7), .B1(new_n370), .B2(G953), .ZN(new_n409));
  OR2_X1    g223(.A1(new_n369), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n369), .A2(new_n409), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n375), .A2(new_n260), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n383), .A2(new_n386), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n414), .A2(new_n388), .ZN(new_n415));
  XOR2_X1   g229(.A(new_n389), .B(KEYINPUT8), .Z(new_n416));
  OAI211_X1 g230(.A(new_n410), .B(new_n411), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n400), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n289), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n366), .B1(new_n408), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n372), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n400), .A2(KEYINPUT6), .B1(new_n402), .B2(new_n404), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n402), .A2(KEYINPUT6), .A3(new_n404), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n410), .A2(new_n411), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n416), .B1(new_n414), .B2(new_n388), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(G902), .B1(new_n427), .B2(new_n400), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n424), .A2(new_n365), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n420), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(KEYINPUT9), .B(G234), .ZN(new_n431));
  OAI21_X1  g245(.A(G221), .B1(new_n431), .B2(G902), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G469), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(new_n289), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n233), .A2(new_n398), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n395), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n232), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT10), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n368), .A2(new_n387), .A3(new_n439), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n210), .A2(new_n383), .A3(new_n386), .A4(new_n215), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT10), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n437), .A2(new_n438), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n210), .A2(new_n215), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n413), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n441), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n447), .A2(KEYINPUT12), .A3(new_n232), .ZN(new_n448));
  AOI21_X1  g262(.A(KEYINPUT12), .B1(new_n447), .B2(new_n232), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n444), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(G110), .B(G140), .ZN(new_n451));
  INV_X1    g265(.A(G227), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(G953), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n451), .B(new_n453), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n395), .A2(new_n436), .B1(new_n440), .B2(new_n442), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n454), .B1(new_n455), .B2(new_n438), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n437), .A2(new_n443), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n232), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n450), .A2(new_n454), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n435), .B1(new_n459), .B2(G469), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n437), .A2(new_n438), .A3(new_n443), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n438), .B1(new_n437), .B2(new_n443), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n454), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n454), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n444), .B(new_n464), .C1(new_n448), .C2(new_n449), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n434), .A3(new_n289), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n433), .B1(new_n460), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(G214), .B1(G237), .B2(G902), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n430), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n239), .A2(G143), .A3(G214), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(G143), .B1(new_n239), .B2(G214), .ZN(new_n474));
  OAI21_X1  g288(.A(G131), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT17), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT80), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n474), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n201), .B1(new_n478), .B2(new_n472), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT80), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(new_n480), .A3(KEYINPUT17), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n478), .A2(new_n201), .A3(new_n472), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n475), .A2(new_n483), .A3(new_n476), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n341), .A3(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(G113), .B(G122), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(new_n376), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n478), .A2(KEYINPUT18), .A3(G131), .A4(new_n472), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT18), .ZN(new_n489));
  OAI22_X1  g303(.A1(new_n473), .A2(new_n474), .B1(new_n489), .B2(new_n201), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n333), .A2(new_n334), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G146), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT78), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n493), .A2(new_n319), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n494), .B1(new_n493), .B2(new_n319), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n491), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n485), .A2(new_n487), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n487), .B1(new_n485), .B2(new_n497), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n289), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(G475), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n475), .A2(new_n483), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n318), .A2(KEYINPUT19), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n318), .A2(KEYINPUT19), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n187), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n323), .A2(G146), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n503), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT79), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n497), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n487), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n509), .B1(new_n497), .B2(new_n508), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n498), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT20), .ZN(new_n515));
  NOR2_X1   g329(.A1(G475), .A2(G902), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n515), .B1(new_n514), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n502), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n431), .A2(new_n357), .A3(G953), .ZN(new_n520));
  XOR2_X1   g334(.A(new_n520), .B(KEYINPUT89), .Z(new_n521));
  INV_X1    g335(.A(KEYINPUT85), .ZN(new_n522));
  INV_X1    g336(.A(G122), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n522), .B(KEYINPUT14), .C1(new_n523), .C2(G116), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(G116), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G116), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(G122), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n522), .B1(new_n528), .B2(KEYINPUT14), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT86), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT14), .B1(new_n523), .B2(G116), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT85), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT86), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n532), .A2(new_n533), .A3(new_n525), .A4(new_n524), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT14), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n527), .A3(G122), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT87), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n535), .A2(new_n527), .A3(KEYINPUT87), .A4(G122), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n530), .A2(new_n534), .A3(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n541), .A2(KEYINPUT88), .A3(G107), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT88), .B1(new_n541), .B2(G107), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n525), .A2(new_n528), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT81), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n525), .A2(new_n528), .A3(KEYINPUT81), .ZN(new_n547));
  AOI21_X1  g361(.A(G107), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n189), .A2(G128), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n214), .A2(G143), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT84), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT84), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(new_n197), .ZN(new_n557));
  AOI21_X1  g371(.A(G134), .B1(new_n554), .B2(new_n555), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n549), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n542), .A2(new_n543), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n558), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n546), .A2(G107), .A3(new_n547), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n561), .B1(new_n563), .B2(new_n548), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT82), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n189), .A2(G128), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT13), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n565), .B(new_n550), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n568), .A2(G134), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n550), .B1(new_n566), .B2(new_n567), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n570), .B(KEYINPUT82), .C1(new_n567), .C2(new_n550), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT83), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n571), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT83), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n564), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n521), .B1(new_n560), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT90), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n575), .A2(new_n573), .ZN(new_n579));
  INV_X1    g393(.A(new_n564), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n521), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n556), .B(new_n197), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n538), .A2(new_n539), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n532), .A2(new_n525), .A3(new_n524), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n584), .B1(new_n585), .B2(KEYINPUT86), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n379), .B1(new_n586), .B2(new_n534), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n549), .B(new_n583), .C1(new_n587), .C2(KEYINPUT88), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n581), .B(new_n582), .C1(new_n588), .C2(new_n542), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n577), .A2(new_n578), .A3(new_n589), .ZN(new_n590));
  OAI211_X1 g404(.A(KEYINPUT90), .B(new_n521), .C1(new_n560), .C2(new_n576), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n289), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT91), .ZN(new_n593));
  INV_X1    g407(.A(G478), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(KEYINPUT15), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT91), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n590), .A2(new_n596), .A3(new_n289), .A4(new_n591), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n593), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n595), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n590), .A2(new_n289), .A3(new_n599), .A4(new_n591), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n600), .A2(KEYINPUT92), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT92), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n593), .A2(new_n603), .A3(new_n595), .A4(new_n597), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n519), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT93), .ZN(new_n606));
  NAND2_X1  g420(.A1(G234), .A2(G237), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(G952), .A3(new_n344), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(G902), .A3(G953), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT21), .B(G898), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n605), .A2(new_n606), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n606), .B1(new_n605), .B2(new_n614), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n364), .B(new_n471), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G101), .ZN(G3));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n590), .A2(new_n619), .A3(new_n591), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n577), .A2(KEYINPUT33), .A3(new_n589), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n594), .A2(G902), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT94), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n593), .A2(new_n594), .A3(new_n597), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT94), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n620), .A2(new_n626), .A3(new_n621), .A4(new_n622), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n469), .ZN(new_n629));
  AOI211_X1 g443(.A(new_n613), .B(new_n629), .C1(new_n420), .C2(new_n429), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n628), .A2(new_n519), .A3(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(G472), .B1(new_n276), .B2(G902), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n633), .B1(new_n276), .B2(new_n277), .ZN(new_n634));
  INV_X1    g448(.A(new_n468), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n634), .A2(new_n363), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT34), .B(G104), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT95), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n637), .B(new_n639), .ZN(G6));
  INV_X1    g454(.A(new_n519), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n602), .A2(new_n630), .A3(new_n604), .A4(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n636), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT96), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT35), .B(G107), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G9));
  OR2_X1    g461(.A1(new_n347), .A2(KEYINPUT36), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n342), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n342), .A2(new_n648), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n361), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n356), .A2(new_n358), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n352), .A2(KEYINPUT74), .A3(new_n353), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n634), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n471), .B(new_n657), .C1(new_n615), .C2(new_n616), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT37), .B(G110), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT97), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n658), .B(new_n660), .ZN(G12));
  NOR3_X1   g475(.A1(new_n297), .A2(new_n470), .A3(new_n656), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n344), .A2(G900), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(G902), .A3(new_n607), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n664), .A2(KEYINPUT98), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n664), .A2(KEYINPUT98), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n665), .A2(new_n666), .A3(new_n609), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n667), .B(KEYINPUT99), .Z(new_n668));
  AND4_X1   g482(.A1(new_n602), .A2(new_n604), .A3(new_n641), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n662), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  XNOR2_X1  g485(.A(new_n430), .B(KEYINPUT38), .ZN(new_n672));
  AND4_X1   g486(.A1(new_n519), .A2(new_n672), .A3(new_n469), .A4(new_n656), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n602), .A2(new_n604), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n272), .A2(new_n278), .ZN(new_n675));
  NAND2_X1  g489(.A1(G472), .A2(G902), .ZN(new_n676));
  INV_X1    g490(.A(new_n245), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n235), .A2(new_n236), .ZN(new_n678));
  OAI21_X1  g492(.A(G472), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n676), .B1(new_n679), .B2(new_n255), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT100), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n668), .B(KEYINPUT39), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n468), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n684), .B(KEYINPUT40), .Z(new_n685));
  NAND4_X1  g499(.A1(new_n673), .A2(new_n674), .A3(new_n682), .A4(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT101), .B(G143), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G45));
  AND3_X1   g502(.A1(new_n628), .A2(new_n519), .A3(new_n668), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n662), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  NAND2_X1  g505(.A1(new_n296), .A2(G472), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n675), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n363), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n466), .A2(new_n289), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(G469), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n467), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n433), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n693), .A2(new_n694), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n631), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT41), .B(G113), .Z(new_n701));
  XOR2_X1   g515(.A(new_n701), .B(KEYINPUT102), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n700), .B(new_n702), .ZN(G15));
  NOR2_X1   g517(.A1(new_n699), .A2(new_n642), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n527), .ZN(G18));
  AOI21_X1  g519(.A(new_n434), .B1(new_n466), .B2(new_n289), .ZN(new_n706));
  AOI211_X1 g520(.A(G469), .B(G902), .C1(new_n463), .C2(new_n465), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n430), .A2(new_n708), .A3(new_n469), .A4(new_n432), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n297), .A2(new_n709), .A3(new_n656), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n710), .B1(new_n615), .B2(new_n616), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G119), .ZN(G21));
  AND2_X1   g526(.A1(new_n283), .A2(new_n284), .ZN(new_n713));
  OAI22_X1  g527(.A1(new_n257), .A2(new_n268), .B1(new_n713), .B2(new_n677), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n271), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n633), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n697), .A2(new_n613), .A3(new_n433), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n717), .A3(new_n694), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n408), .A2(new_n366), .A3(new_n419), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n365), .B1(new_n424), .B2(new_n428), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n519), .B(new_n469), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n602), .A3(new_n604), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n523), .ZN(G24));
  OAI21_X1  g539(.A(new_n652), .B1(new_n354), .B2(new_n359), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n633), .A2(new_n715), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n709), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(new_n519), .A3(new_n628), .A4(new_n668), .ZN(new_n729));
  XOR2_X1   g543(.A(KEYINPUT103), .B(G125), .Z(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G27));
  INV_X1    g545(.A(KEYINPUT104), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n270), .B1(new_n269), .B2(new_n271), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n276), .A2(KEYINPUT32), .A3(new_n277), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n272), .A2(new_n278), .A3(KEYINPUT104), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n692), .A3(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n468), .A2(new_n469), .A3(new_n420), .A4(new_n429), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT42), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n689), .A2(new_n694), .A3(new_n737), .A4(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n738), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n693), .A2(new_n742), .A3(new_n694), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n628), .A2(new_n519), .A3(new_n668), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n739), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G131), .ZN(G33));
  NAND3_X1  g561(.A1(new_n669), .A2(new_n364), .A3(new_n742), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  NAND2_X1  g563(.A1(new_n459), .A2(KEYINPUT45), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT105), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n459), .A2(KEYINPUT45), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n434), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT106), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT106), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n752), .A2(new_n757), .A3(new_n754), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n435), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  OR3_X1    g573(.A1(new_n759), .A2(KEYINPUT107), .A3(KEYINPUT46), .ZN(new_n760));
  OAI21_X1  g574(.A(KEYINPUT107), .B1(new_n759), .B2(KEYINPUT46), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n707), .B1(new_n759), .B2(KEYINPUT46), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n432), .ZN(new_n764));
  INV_X1    g578(.A(new_n683), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n420), .A2(new_n469), .A3(new_n429), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n628), .A2(new_n641), .ZN(new_n769));
  XOR2_X1   g583(.A(new_n769), .B(KEYINPUT43), .Z(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n634), .A3(new_n726), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n766), .A2(new_n768), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G137), .ZN(G39));
  INV_X1    g590(.A(KEYINPUT47), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n764), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n763), .A2(KEYINPUT47), .A3(new_n432), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR4_X1   g594(.A1(new_n744), .A2(new_n693), .A3(new_n694), .A4(new_n767), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(KEYINPUT108), .B(G140), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(G42));
  NOR2_X1   g598(.A1(new_n682), .A2(new_n363), .ZN(new_n785));
  INV_X1    g599(.A(new_n698), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n786), .A2(new_n767), .A3(new_n608), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n628), .A2(new_n519), .ZN(new_n789));
  OAI211_X1 g603(.A(G952), .B(new_n344), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n716), .A2(new_n694), .A3(new_n609), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n770), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n709), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n770), .A2(new_n787), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT118), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n737), .A2(new_n694), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n798), .A2(KEYINPUT48), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(KEYINPUT48), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n794), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n796), .A2(new_n727), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n788), .A2(new_n519), .A3(new_n628), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n697), .A2(new_n432), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n780), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n792), .A2(new_n768), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n804), .B(KEYINPUT51), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT51), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n672), .A2(new_n469), .A3(new_n786), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n770), .A2(new_n791), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT50), .B1(new_n814), .B2(KEYINPUT115), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n815), .B1(KEYINPUT115), .B2(new_n814), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n816), .A2(KEYINPUT116), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(KEYINPUT116), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n792), .A2(KEYINPUT50), .A3(new_n813), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n801), .B1(new_n812), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n780), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT114), .B1(new_n778), .B2(new_n779), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n823), .A2(new_n805), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n804), .B1(new_n825), .B2(new_n807), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n820), .A2(new_n809), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n810), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n821), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n617), .A2(new_n658), .A3(new_n637), .A4(new_n644), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  OAI22_X1  g645(.A1(new_n699), .A2(new_n631), .B1(new_n723), .B2(new_n718), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n704), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(new_n711), .A3(new_n746), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n727), .A2(new_n738), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n689), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n668), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n738), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n605), .A2(new_n838), .A3(new_n693), .A4(new_n726), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n748), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n834), .A2(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n722), .A2(new_n602), .A3(new_n604), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT109), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n450), .A2(new_n454), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n456), .A2(new_n458), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n844), .A2(G469), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n435), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n432), .B(new_n668), .C1(new_n848), .C2(new_n707), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n843), .B1(new_n849), .B2(new_n726), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n656), .A2(new_n468), .A3(KEYINPUT109), .A4(new_n668), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n850), .A2(new_n851), .B1(new_n675), .B2(new_n681), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n842), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n690), .A2(new_n670), .A3(new_n729), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT52), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n662), .B1(new_n689), .B2(new_n669), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n857), .A3(new_n729), .A4(new_n853), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n831), .A2(new_n841), .A3(new_n855), .A4(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g675(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT54), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n859), .A2(new_n862), .ZN(new_n866));
  AND4_X1   g680(.A1(KEYINPUT53), .A2(new_n748), .A3(new_n836), .A4(new_n839), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n855), .A2(new_n858), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n830), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n834), .A2(KEYINPUT111), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT111), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n833), .A2(new_n711), .A3(new_n746), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT112), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n869), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n874), .B1(new_n869), .B2(new_n873), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n865), .B(new_n866), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n864), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT113), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n829), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(G952), .A2(G953), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n629), .B(new_n433), .C1(new_n697), .C2(KEYINPUT49), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(KEYINPUT49), .B2(new_n697), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(new_n672), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n785), .ZN(new_n885));
  OAI22_X1  g699(.A1(new_n880), .A2(new_n881), .B1(new_n769), .B2(new_n885), .ZN(G75));
  NOR2_X1   g700(.A1(new_n344), .A2(G952), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n866), .B1(new_n875), .B2(new_n876), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n888), .A2(G902), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(G210), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT56), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n422), .A2(new_n423), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n372), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n424), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT55), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n887), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n890), .A2(KEYINPUT119), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n889), .A2(new_n899), .A3(G210), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n896), .A2(KEYINPUT56), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n897), .A2(new_n902), .ZN(G51));
  NAND2_X1  g717(.A1(new_n888), .A2(KEYINPUT54), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n904), .A2(KEYINPUT120), .A3(new_n877), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT120), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n888), .A2(new_n906), .A3(KEYINPUT54), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n435), .B(KEYINPUT57), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n905), .A2(KEYINPUT121), .A3(new_n907), .A4(new_n908), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n911), .A2(new_n466), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n889), .A2(new_n758), .A3(new_n756), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n887), .B1(new_n913), .B2(new_n914), .ZN(G54));
  NAND3_X1  g729(.A1(new_n889), .A2(KEYINPUT58), .A3(G475), .ZN(new_n916));
  INV_X1    g730(.A(new_n514), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n887), .ZN(G60));
  XOR2_X1   g734(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n921));
  NOR2_X1   g735(.A1(new_n594), .A2(new_n289), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  AOI22_X1  g738(.A1(new_n879), .A2(new_n924), .B1(new_n620), .B2(new_n621), .ZN(new_n925));
  INV_X1    g739(.A(new_n887), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n905), .A2(new_n907), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n620), .A2(new_n621), .A3(new_n924), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n925), .A2(new_n929), .ZN(G63));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT60), .Z(new_n932));
  NAND2_X1  g746(.A1(new_n888), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n360), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n888), .A2(new_n651), .A3(new_n932), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n934), .A2(new_n926), .A3(new_n935), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g751(.A(G953), .B1(new_n612), .B2(new_n370), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n831), .A2(new_n711), .A3(new_n833), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n938), .B1(new_n939), .B2(G953), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n893), .B1(G898), .B2(new_n344), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(G69));
  XOR2_X1   g756(.A(new_n258), .B(KEYINPUT123), .Z(new_n943));
  NOR2_X1   g757(.A1(new_n504), .A2(new_n505), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n943), .B(new_n944), .Z(new_n945));
  NAND2_X1  g759(.A1(new_n674), .A2(new_n641), .ZN(new_n946));
  AOI211_X1 g760(.A(new_n765), .B(new_n743), .C1(new_n946), .C2(new_n789), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n782), .A2(new_n775), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n856), .A2(new_n729), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT124), .Z(new_n951));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n951), .A2(new_n952), .A3(new_n686), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n952), .B1(new_n951), .B2(new_n686), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n949), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n945), .B1(new_n956), .B2(G953), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n663), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n766), .A2(new_n694), .A3(new_n842), .A4(new_n737), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n782), .A2(new_n960), .A3(new_n746), .A4(new_n748), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n775), .A2(new_n951), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(KEYINPUT126), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n775), .A2(new_n964), .A3(new_n951), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n961), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n945), .A2(G953), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OAI211_X1 g782(.A(KEYINPUT125), .B(new_n959), .C1(new_n966), .C2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n958), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n663), .B1(new_n452), .B2(G953), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(G72));
  NOR2_X1   g786(.A1(new_n253), .A2(new_n235), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n956), .A2(new_n939), .ZN(new_n974));
  XNOR2_X1  g788(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(new_n676), .ZN(new_n976));
  AOI211_X1 g790(.A(new_n285), .B(new_n973), .C1(new_n974), .C2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n973), .A2(new_n285), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n966), .A2(new_n939), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n978), .B1(new_n979), .B2(new_n976), .ZN(new_n980));
  INV_X1    g794(.A(new_n294), .ZN(new_n981));
  OAI221_X1 g795(.A(new_n976), .B1(new_n255), .B2(new_n981), .C1(new_n861), .C2(new_n863), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n926), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n977), .A2(new_n980), .A3(new_n983), .ZN(G57));
endmodule


