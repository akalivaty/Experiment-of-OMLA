//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n996, new_n997;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G8gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(KEYINPUT97), .A3(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n203), .B1(new_n202), .B2(KEYINPUT97), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n202), .A2(new_n207), .ZN(new_n208));
  OAI22_X1  g007(.A1(new_n205), .A2(new_n206), .B1(new_n208), .B2(G1gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n206), .ZN(new_n210));
  AOI21_X1  g009(.A(G1gat), .B1(new_n202), .B2(new_n207), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(new_n211), .A3(new_n204), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G43gat), .B(G50gat), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(KEYINPUT15), .ZN(new_n217));
  XOR2_X1   g016(.A(G43gat), .B(G50gat), .Z(new_n218));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G29gat), .ZN(new_n221));
  INV_X1    g020(.A(G36gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT14), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT14), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G29gat), .B2(G36gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT96), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n223), .A2(new_n225), .A3(KEYINPUT96), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n217), .A2(new_n220), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  OAI211_X1 g029(.A(KEYINPUT15), .B(new_n216), .C1(new_n226), .C2(new_n215), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT17), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n232), .B1(new_n230), .B2(new_n231), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n213), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n230), .A2(new_n231), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(new_n212), .A3(new_n209), .ZN(new_n237));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n235), .A2(KEYINPUT18), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n230), .A2(new_n231), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n213), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n237), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n238), .B(KEYINPUT13), .Z(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n239), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT18), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G141gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(G197gat), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT11), .B(G169gat), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT12), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT95), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n249), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n253), .B(KEYINPUT12), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n248), .A2(new_n244), .A3(new_n239), .A4(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n259), .A2(KEYINPUT98), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT98), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n255), .B1(new_n247), .B2(new_n246), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n261), .B1(new_n245), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n257), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(KEYINPUT91), .B(KEYINPUT38), .Z(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT37), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT75), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT22), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G211gat), .A2(G218gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(KEYINPUT75), .A2(KEYINPUT22), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G197gat), .B(G204gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G211gat), .B(G218gat), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n274), .A2(new_n277), .A3(new_n275), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G226gat), .ZN(new_n283));
  INV_X1    g082(.A(G233gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT26), .ZN(new_n288));
  OR2_X1    g087(.A1(new_n287), .A2(KEYINPUT26), .ZN(new_n289));
  INV_X1    g088(.A(G169gat), .ZN(new_n290));
  INV_X1    g089(.A(G176gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n286), .B(new_n288), .C1(new_n289), .C2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n294));
  INV_X1    g093(.A(G190gat), .ZN(new_n295));
  INV_X1    g094(.A(G183gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(KEYINPUT27), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n295), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT27), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G183gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n296), .A2(KEYINPUT27), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT69), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n294), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT28), .A4(new_n295), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n293), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n286), .A2(KEYINPUT24), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT24), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n309), .A2(G183gat), .A3(G190gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n312));
  OR3_X1    g111(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AND4_X1   g113(.A1(KEYINPUT65), .A2(new_n290), .A3(new_n291), .A4(KEYINPUT23), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT65), .B1(new_n287), .B2(KEYINPUT23), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n287), .ZN(new_n318));
  OAI22_X1  g117(.A1(new_n290), .A2(new_n291), .B1(KEYINPUT66), .B2(KEYINPUT23), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT66), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT23), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n318), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n314), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT25), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n287), .A2(KEYINPUT23), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n323), .A2(KEYINPUT25), .A3(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n296), .A2(KEYINPUT24), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n329), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n286), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT67), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(new_n296), .A3(new_n295), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT68), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n333), .ZN(new_n336));
  NOR3_X1   g135(.A1(KEYINPUT67), .A2(G183gat), .A3(G190gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT68), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n339), .A3(new_n311), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n328), .B1(new_n335), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n307), .B1(new_n326), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n285), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n335), .A2(new_n340), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n327), .A2(KEYINPUT25), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n320), .A2(new_n321), .B1(G169gat), .B2(G176gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n347), .B1(new_n320), .B2(new_n321), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n346), .B1(new_n348), .B2(new_n318), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n345), .A2(new_n349), .B1(new_n324), .B2(new_n325), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n285), .B1(new_n350), .B2(new_n306), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n282), .B1(new_n344), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n285), .ZN(new_n354));
  NOR3_X1   g153(.A1(new_n330), .A2(new_n334), .A3(KEYINPUT68), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n339), .B1(new_n338), .B2(new_n311), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n349), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n324), .A2(new_n325), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n306), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n354), .B1(new_n359), .B2(KEYINPUT29), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(new_n281), .A3(new_n351), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n268), .B1(new_n353), .B2(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(G8gat), .B(G36gat), .Z(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT76), .ZN(new_n364));
  XNOR2_X1  g163(.A(G64gat), .B(G92gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT93), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n361), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n368), .B1(KEYINPUT37), .B2(new_n369), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n362), .A2(KEYINPUT93), .A3(new_n367), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n267), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G113gat), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n373), .A2(KEYINPUT71), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(KEYINPUT71), .ZN(new_n375));
  OAI21_X1  g174(.A(G120gat), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G120gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G127gat), .B(G134gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT72), .B(KEYINPUT1), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n376), .A2(new_n378), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(KEYINPUT70), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT1), .B1(G113gat), .B2(G120gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G127gat), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n385), .A2(KEYINPUT70), .A3(G134gat), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n382), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n381), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n390));
  INV_X1    g189(.A(G148gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n390), .B1(new_n391), .B2(G141gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(G141gat), .ZN(new_n393));
  INV_X1    g192(.A(G141gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(KEYINPUT77), .A3(G148gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(G155gat), .ZN(new_n397));
  INV_X1    g196(.A(G162gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G155gat), .A2(G162gat), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(KEYINPUT78), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT78), .ZN(new_n402));
  AND2_X1   g201(.A1(G155gat), .A2(G162gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(G155gat), .A2(G162gat), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n400), .A2(KEYINPUT2), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n396), .A2(new_n401), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT3), .ZN(new_n408));
  XNOR2_X1  g207(.A(G141gat), .B(G148gat), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n400), .B(new_n399), .C1(new_n409), .C2(KEYINPUT2), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n407), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  AND2_X1   g210(.A1(new_n389), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n407), .A2(new_n410), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT79), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n407), .A2(new_n415), .A3(new_n410), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n412), .B1(new_n417), .B2(new_n408), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n381), .A2(new_n388), .A3(new_n407), .A4(new_n410), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT4), .ZN(new_n420));
  NAND2_X1  g219(.A1(G225gat), .A2(G233gat), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  OR2_X1    g221(.A1(new_n422), .A2(KEYINPUT5), .ZN(new_n423));
  INV_X1    g222(.A(new_n421), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n407), .A2(new_n415), .A3(new_n410), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n415), .B1(new_n407), .B2(new_n410), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n379), .A2(new_n380), .A3(new_n378), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n386), .B1(new_n379), .B2(KEYINPUT70), .ZN(new_n428));
  AOI22_X1  g227(.A1(new_n427), .A2(new_n376), .B1(new_n428), .B2(new_n384), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n425), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n419), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n424), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT80), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(KEYINPUT80), .B(new_n424), .C1(new_n430), .C2(new_n431), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n434), .A2(new_n422), .A3(KEYINPUT5), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n423), .A2(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(G1gat), .B(G29gat), .Z(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G57gat), .B(G85gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n443));
  OR2_X1    g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(new_n443), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n437), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n423), .A2(new_n436), .A3(new_n443), .A4(new_n442), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n360), .A2(new_n281), .A3(new_n351), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n281), .B1(new_n360), .B2(new_n351), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n448), .B1(new_n367), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n362), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT90), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n366), .B(new_n266), .C1(new_n369), .C2(KEYINPUT37), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n362), .A2(KEYINPUT90), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT92), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT92), .ZN(new_n461));
  NOR4_X1   g260(.A1(new_n455), .A2(new_n457), .A3(new_n458), .A4(new_n461), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n372), .B(new_n452), .C1(new_n460), .C2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n366), .B1(new_n449), .B2(new_n450), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n353), .A2(new_n367), .A3(new_n361), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT30), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT30), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n467), .A3(new_n367), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT89), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n466), .A2(KEYINPUT89), .A3(new_n468), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n421), .B1(new_n418), .B2(new_n420), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT39), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n442), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n419), .B1(new_n417), .B2(new_n429), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT39), .B1(new_n477), .B2(new_n424), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n476), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n479), .B(KEYINPUT40), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n437), .A2(new_n442), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n473), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(G228gat), .A2(G233gat), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n274), .A2(new_n277), .A3(new_n275), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n277), .B1(new_n274), .B2(new_n275), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n343), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n486), .A2(new_n408), .B1(new_n410), .B2(new_n407), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n281), .B1(new_n411), .B2(new_n343), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n483), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT83), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g290(.A(KEYINPUT83), .B(new_n483), .C1(new_n487), .C2(new_n488), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n486), .A2(new_n408), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n493), .A2(new_n414), .A3(new_n416), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n488), .A2(new_n483), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n491), .A2(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(G22gat), .B1(new_n496), .B2(KEYINPUT86), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n491), .A2(new_n492), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n495), .A2(new_n494), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n498), .A2(KEYINPUT86), .A3(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT87), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n498), .A2(new_n499), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT86), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT87), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n496), .A2(KEYINPUT86), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n504), .A2(new_n505), .A3(G22gat), .A4(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(KEYINPUT84), .B(G22gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n496), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G78gat), .B(G106gat), .ZN(new_n510));
  INV_X1    g309(.A(G50gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n512), .B(new_n513), .Z(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n509), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n507), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT85), .ZN(new_n519));
  INV_X1    g318(.A(new_n508), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n509), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n519), .B1(new_n522), .B2(new_n514), .ZN(new_n523));
  AOI211_X1 g322(.A(KEYINPUT85), .B(new_n515), .C1(new_n521), .C2(new_n509), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n518), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n463), .A2(new_n482), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n429), .B1(new_n350), .B2(new_n306), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n307), .B(new_n389), .C1(new_n326), .C2(new_n341), .ZN(new_n528));
  INV_X1    g327(.A(G227gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n529), .A2(new_n284), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(G71gat), .B(G99gat), .Z(new_n532));
  XNOR2_X1  g331(.A(G15gat), .B(G43gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT33), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(KEYINPUT32), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT73), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT73), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n531), .A2(new_n538), .A3(KEYINPUT32), .A4(new_n535), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n531), .A2(KEYINPUT32), .ZN(new_n541));
  INV_X1    g340(.A(new_n531), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n541), .B(new_n534), .C1(new_n542), .C2(KEYINPUT33), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT34), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n528), .ZN(new_n546));
  INV_X1    g345(.A(new_n530), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI211_X1 g347(.A(KEYINPUT34), .B(new_n530), .C1(new_n527), .C2(new_n528), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n544), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n540), .A2(new_n550), .A3(new_n543), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT36), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n554), .B1(KEYINPUT74), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(KEYINPUT74), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n448), .A2(new_n469), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT88), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n525), .B(new_n560), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n526), .B(new_n558), .C1(new_n559), .C2(new_n561), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n540), .A2(new_n550), .A3(new_n543), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n550), .B1(new_n540), .B2(new_n543), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT35), .B1(new_n446), .B2(new_n447), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n565), .A2(new_n472), .A3(new_n471), .A4(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n497), .A2(new_n500), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n516), .B1(new_n568), .B2(new_n505), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n498), .A2(new_n499), .A3(new_n508), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n508), .B1(new_n498), .B2(new_n499), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n514), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT85), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n522), .A2(new_n519), .A3(new_n514), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n569), .A2(new_n501), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT94), .B1(new_n567), .B2(new_n575), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n566), .A2(new_n552), .A3(new_n553), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT94), .ZN(new_n578));
  INV_X1    g377(.A(new_n472), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT89), .B1(new_n466), .B2(new_n468), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n577), .A2(new_n525), .A3(new_n578), .A4(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n576), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n525), .A2(new_n559), .A3(new_n565), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT35), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n265), .B1(new_n562), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT104), .ZN(new_n589));
  AND2_X1   g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT103), .ZN(new_n593));
  NAND2_X1  g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  INV_X1    g393(.A(G85gat), .ZN(new_n595));
  INV_X1    g394(.A(G92gat), .ZN(new_n596));
  AOI22_X1  g395(.A1(KEYINPUT8), .A2(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G85gat), .A2(G92gat), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT7), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n597), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G99gat), .B(G106gat), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n600), .A2(new_n601), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n603), .B1(new_n606), .B2(new_n597), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n593), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n602), .A2(new_n604), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n606), .A2(new_n603), .A3(new_n597), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(KEYINPUT103), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n592), .B1(new_n612), .B2(new_n240), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n612), .B1(new_n233), .B2(new_n234), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n614), .B(new_n615), .C1(KEYINPUT104), .C2(new_n588), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n617));
  XNOR2_X1  g416(.A(G134gat), .B(G162gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n588), .A2(KEYINPUT104), .ZN(new_n620));
  INV_X1    g419(.A(new_n615), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n620), .B1(new_n621), .B2(new_n613), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n616), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n619), .B1(new_n616), .B2(new_n622), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(G71gat), .A2(G78gat), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G71gat), .A2(G78gat), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(KEYINPUT99), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT9), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(G57gat), .ZN(new_n635));
  INV_X1    g434(.A(G64gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G57gat), .A2(G64gat), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n634), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n640));
  INV_X1    g439(.A(new_n631), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n640), .B1(new_n641), .B2(new_n629), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n632), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n630), .A2(new_n631), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT100), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n636), .B1(new_n645), .B2(new_n635), .ZN(new_n646));
  NAND3_X1  g445(.A1(KEYINPUT100), .A2(G57gat), .A3(G64gat), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n644), .A2(new_n646), .A3(new_n634), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n649), .B1(new_n605), .B2(new_n607), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT10), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n609), .A2(new_n610), .A3(new_n643), .A4(new_n648), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n649), .A2(new_n651), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n654), .A2(new_n608), .A3(new_n611), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n628), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n650), .A2(new_n652), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n656), .B1(new_n628), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G120gat), .B(G148gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT105), .ZN(new_n660));
  XNOR2_X1  g459(.A(G176gat), .B(G204gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n658), .A2(new_n662), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(G183gat), .B(G211gat), .Z(new_n667));
  INV_X1    g466(.A(KEYINPUT21), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n649), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(KEYINPUT101), .Z(new_n670));
  INV_X1    g469(.A(KEYINPUT102), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n670), .B(KEYINPUT102), .ZN(new_n675));
  INV_X1    g474(.A(new_n673), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n667), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n213), .B1(new_n668), .B2(new_n649), .ZN(new_n679));
  XNOR2_X1  g478(.A(G127gat), .B(G155gat), .ZN(new_n680));
  NAND2_X1  g479(.A1(G231gat), .A2(G233gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n679), .B(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n672), .A2(new_n673), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n675), .A2(new_n676), .ZN(new_n685));
  INV_X1    g484(.A(new_n667), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n678), .A2(new_n683), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n683), .B1(new_n678), .B2(new_n687), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n626), .B(new_n666), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n587), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n448), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g495(.A(KEYINPUT16), .B(G8gat), .Z(new_n697));
  NAND3_X1  g496(.A1(new_n693), .A2(new_n473), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G8gat), .B1(new_n692), .B2(new_n581), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  MUX2_X1   g499(.A(new_n698), .B(new_n700), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g500(.A(G15gat), .B1(new_n692), .B2(new_n558), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n554), .A2(G15gat), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n692), .B2(new_n703), .ZN(G1326gat));
  NOR2_X1   g503(.A1(new_n692), .A2(new_n561), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT43), .B(G22gat), .Z(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1327gat));
  NOR2_X1   g506(.A1(new_n688), .A2(new_n689), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(new_n626), .A3(new_n665), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n587), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n448), .A2(G29gat), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT45), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AND4_X1   g513(.A1(KEYINPUT45), .A2(new_n587), .A3(new_n710), .A4(new_n713), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI221_X4 g515(.A(KEYINPUT107), .B1(new_n584), .B2(KEYINPUT35), .C1(new_n576), .C2(new_n582), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n718), .B1(new_n583), .B2(new_n585), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n562), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(KEYINPUT44), .B1(new_n720), .B2(new_n625), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722));
  AOI211_X1 g521(.A(new_n722), .B(new_n626), .C1(new_n562), .C2(new_n586), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n709), .A2(new_n665), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n264), .A2(KEYINPUT106), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n259), .A2(KEYINPUT98), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n245), .A2(new_n262), .A3(new_n261), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n728), .A2(new_n729), .A3(new_n257), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n724), .A2(new_n731), .ZN(new_n732));
  NOR4_X1   g531(.A1(new_n721), .A2(new_n723), .A3(new_n448), .A4(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n716), .B1(new_n733), .B2(new_n221), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n716), .B(KEYINPUT108), .C1(new_n221), .C2(new_n733), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(G1328gat));
  NAND2_X1  g537(.A1(new_n473), .A2(new_n222), .ZN(new_n739));
  OAI21_X1  g538(.A(KEYINPUT46), .B1(new_n711), .B2(new_n739), .ZN(new_n740));
  OR3_X1    g539(.A1(new_n711), .A2(KEYINPUT46), .A3(new_n739), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n720), .A2(new_n625), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n722), .ZN(new_n743));
  INV_X1    g542(.A(new_n723), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n745), .A2(new_n581), .A3(new_n732), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n740), .B(new_n741), .C1(new_n746), .C2(new_n222), .ZN(G1329gat));
  INV_X1    g546(.A(new_n558), .ZN(new_n748));
  INV_X1    g547(.A(new_n732), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n743), .A2(new_n748), .A3(new_n744), .A4(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n721), .A2(new_n723), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n753), .A2(KEYINPUT110), .A3(new_n748), .A4(new_n749), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n752), .A2(G43gat), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT47), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n554), .A2(G43gat), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n756), .B1(new_n712), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n750), .A2(G43gat), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n712), .A2(KEYINPUT109), .A3(new_n757), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n762));
  INV_X1    g561(.A(new_n757), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n711), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n756), .B1(new_n760), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n759), .A2(new_n766), .ZN(G1330gat));
  INV_X1    g566(.A(KEYINPUT48), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n561), .A2(G50gat), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n768), .B1(new_n712), .B2(new_n769), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n745), .A2(new_n525), .A3(new_n732), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(new_n511), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n525), .B(KEYINPUT88), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n753), .A2(new_n773), .A3(new_n749), .ZN(new_n774));
  AOI22_X1  g573(.A1(new_n774), .A2(G50gat), .B1(new_n712), .B2(new_n769), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n772), .B1(new_n775), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g575(.A1(new_n708), .A2(new_n731), .A3(new_n625), .A4(new_n666), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n720), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n694), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g579(.A1(new_n581), .A2(KEYINPUT111), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n581), .A2(KEYINPUT111), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT49), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n778), .B(new_n783), .C1(new_n784), .C2(new_n636), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n636), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1333gat));
  NAND2_X1  g586(.A1(new_n778), .A2(new_n748), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n554), .A2(G71gat), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n788), .A2(G71gat), .B1(new_n778), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g590(.A1(new_n778), .A2(new_n773), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g592(.A1(new_n709), .A2(new_n731), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n665), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n745), .A2(new_n448), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n720), .A2(new_n625), .A3(new_n794), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n720), .A2(KEYINPUT51), .A3(new_n625), .A4(new_n794), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n694), .A2(new_n595), .A3(new_n665), .ZN(new_n803));
  OAI22_X1  g602(.A1(new_n796), .A2(new_n595), .B1(new_n802), .B2(new_n803), .ZN(G1336gat));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n805));
  INV_X1    g604(.A(new_n783), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(G92gat), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n801), .A2(new_n805), .A3(new_n665), .A4(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n795), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n743), .A2(new_n473), .A3(new_n744), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G92gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT52), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n666), .B1(new_n799), .B2(new_n800), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n814), .A2(new_n807), .B1(new_n805), .B2(KEYINPUT52), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n743), .A2(new_n744), .A3(new_n783), .A4(new_n809), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n816), .A2(new_n817), .A3(G92gat), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n813), .A2(new_n819), .ZN(G1337gat));
  INV_X1    g619(.A(G99gat), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n814), .A2(new_n821), .A3(new_n565), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n745), .A2(new_n558), .A3(new_n795), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(new_n821), .ZN(G1338gat));
  NOR2_X1   g623(.A1(new_n525), .A2(G106gat), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n814), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n743), .A2(new_n575), .A3(new_n744), .A4(new_n809), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(G106gat), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n826), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n743), .A2(new_n773), .A3(new_n744), .A4(new_n809), .ZN(new_n831));
  AOI22_X1  g630(.A1(new_n814), .A2(new_n825), .B1(new_n831), .B2(G106gat), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n830), .B1(new_n827), .B2(new_n832), .ZN(G1339gat));
  NAND2_X1  g632(.A1(new_n653), .A2(new_n655), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n627), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n653), .A2(new_n655), .A3(new_n628), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(KEYINPUT54), .A3(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n662), .B1(new_n656), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(KEYINPUT55), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n840), .A2(KEYINPUT113), .A3(new_n664), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n837), .A2(new_n839), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT113), .B1(new_n840), .B2(new_n664), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n725), .A2(new_n730), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n238), .B1(new_n235), .B2(new_n237), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n242), .A2(new_n243), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n253), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n728), .A2(new_n665), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n625), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n728), .A2(new_n854), .A3(new_n851), .ZN(new_n855));
  INV_X1    g654(.A(new_n846), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n856), .A2(new_n625), .A3(new_n841), .A4(new_n844), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n854), .B1(new_n728), .B2(new_n851), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n855), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n708), .B1(new_n853), .B2(new_n859), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n690), .A2(new_n731), .ZN(new_n861));
  AOI211_X1 g660(.A(new_n554), .B(new_n773), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n694), .A3(new_n806), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT115), .ZN(new_n864));
  OAI21_X1  g663(.A(G113gat), .B1(new_n864), .B2(new_n265), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n448), .B1(new_n860), .B2(new_n861), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n525), .A3(new_n565), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n867), .A2(new_n783), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n374), .A2(new_n375), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n869), .A3(new_n731), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n865), .A2(new_n870), .ZN(G1340gat));
  OAI21_X1  g670(.A(G120gat), .B1(new_n864), .B2(new_n666), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n665), .A2(new_n377), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT116), .Z(new_n874));
  NAND2_X1  g673(.A1(new_n868), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n872), .A2(new_n875), .ZN(G1341gat));
  OAI21_X1  g675(.A(G127gat), .B1(new_n864), .B2(new_n708), .ZN(new_n877));
  NOR4_X1   g676(.A1(new_n867), .A2(G127gat), .A3(new_n708), .A4(new_n783), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n877), .A2(KEYINPUT117), .A3(new_n879), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1342gat));
  OAI21_X1  g683(.A(G134gat), .B1(new_n864), .B2(new_n626), .ZN(new_n885));
  NOR4_X1   g684(.A1(new_n867), .A2(G134gat), .A3(new_n473), .A4(new_n626), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT56), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(G1343gat));
  AND3_X1   g687(.A1(new_n866), .A2(new_n575), .A3(new_n558), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n806), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n890), .A2(G141gat), .A3(new_n265), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(KEYINPUT58), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n748), .A2(new_n448), .A3(new_n783), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n561), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n840), .A2(new_n664), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n844), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n852), .B1(new_n265), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n626), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT119), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n859), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n899), .A2(KEYINPUT119), .A3(new_n626), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n709), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n861), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n895), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n860), .A2(new_n861), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT57), .B1(new_n907), .B2(new_n575), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n906), .B1(new_n908), .B2(KEYINPUT118), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT118), .ZN(new_n910));
  AOI211_X1 g709(.A(new_n910), .B(KEYINPUT57), .C1(new_n907), .C2(new_n575), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n893), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(G141gat), .B1(new_n912), .B2(new_n265), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n892), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n731), .B(new_n893), .C1(new_n909), .C2(new_n911), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n915), .A2(new_n916), .A3(G141gat), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n915), .B2(G141gat), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n917), .A2(new_n918), .A3(new_n891), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT58), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n914), .B1(new_n919), .B2(new_n920), .ZN(G1344gat));
  NOR2_X1   g720(.A1(new_n912), .A2(new_n666), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n922), .A2(KEYINPUT59), .A3(new_n391), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT59), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n575), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT57), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n859), .B1(new_n626), .B2(new_n899), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n927), .A2(new_n709), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n690), .A2(new_n264), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n894), .B(new_n773), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n926), .A2(new_n665), .A3(new_n893), .A4(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n924), .B1(new_n931), .B2(G148gat), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n665), .A2(new_n391), .ZN(new_n933));
  OAI22_X1  g732(.A1(new_n923), .A2(new_n932), .B1(new_n890), .B2(new_n933), .ZN(G1345gat));
  NAND2_X1  g733(.A1(new_n709), .A2(G155gat), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT121), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n912), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n397), .B1(new_n890), .B2(new_n708), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT122), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n937), .A2(KEYINPUT122), .A3(new_n938), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1346gat));
  OAI21_X1  g742(.A(G162gat), .B1(new_n912), .B2(new_n626), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n889), .A2(new_n398), .A3(new_n581), .A4(new_n625), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1347gat));
  AOI21_X1  g745(.A(new_n694), .B1(new_n860), .B2(new_n861), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n947), .A2(new_n525), .A3(new_n565), .A4(new_n783), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(G169gat), .B1(new_n949), .B2(new_n731), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n581), .A2(new_n694), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n862), .A2(new_n951), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n952), .A2(new_n290), .A3(new_n265), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n950), .A2(new_n953), .ZN(G1348gat));
  NAND3_X1  g753(.A1(new_n949), .A2(new_n291), .A3(new_n665), .ZN(new_n955));
  OAI21_X1  g754(.A(G176gat), .B1(new_n952), .B2(new_n666), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1349gat));
  AND3_X1   g756(.A1(new_n709), .A2(new_n301), .A3(new_n302), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n862), .A2(new_n709), .A3(new_n951), .ZN(new_n959));
  AOI22_X1  g758(.A1(new_n949), .A2(new_n958), .B1(new_n959), .B2(G183gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n960), .B1(KEYINPUT124), .B2(KEYINPUT60), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT60), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n962), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n964));
  AOI22_X1  g763(.A1(new_n961), .A2(new_n963), .B1(new_n960), .B2(new_n964), .ZN(G1350gat));
  OAI21_X1  g764(.A(G190gat), .B1(new_n952), .B2(new_n626), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT61), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n949), .A2(new_n295), .A3(new_n625), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(G1351gat));
  NOR3_X1   g768(.A1(new_n748), .A2(new_n806), .A3(new_n525), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n970), .A2(new_n947), .ZN(new_n971));
  INV_X1    g770(.A(G197gat), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n971), .A2(new_n972), .A3(new_n731), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n558), .A2(new_n951), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n926), .A2(new_n930), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g774(.A(KEYINPUT125), .B1(new_n975), .B2(new_n265), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(G197gat), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n975), .A2(KEYINPUT125), .A3(new_n265), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n973), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(KEYINPUT126), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n981));
  OAI211_X1 g780(.A(new_n981), .B(new_n973), .C1(new_n977), .C2(new_n978), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n980), .A2(new_n982), .ZN(G1352gat));
  INV_X1    g782(.A(new_n971), .ZN(new_n984));
  NOR3_X1   g783(.A1(new_n984), .A2(G204gat), .A3(new_n666), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT62), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n975), .A2(new_n987), .A3(new_n666), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n987), .B1(new_n975), .B2(new_n666), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(G204gat), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n986), .B1(new_n988), .B2(new_n990), .ZN(G1353gat));
  OAI21_X1  g790(.A(G211gat), .B1(new_n975), .B2(new_n708), .ZN(new_n992));
  XNOR2_X1  g791(.A(new_n992), .B(KEYINPUT63), .ZN(new_n993));
  NOR3_X1   g792(.A1(new_n984), .A2(G211gat), .A3(new_n708), .ZN(new_n994));
  OR2_X1    g793(.A1(new_n993), .A2(new_n994), .ZN(G1354gat));
  OAI21_X1  g794(.A(G218gat), .B1(new_n975), .B2(new_n626), .ZN(new_n996));
  OR2_X1    g795(.A1(new_n626), .A2(G218gat), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n996), .B1(new_n984), .B2(new_n997), .ZN(G1355gat));
endmodule


