//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n578, new_n579, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n634, new_n637, new_n639, new_n640,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1230, new_n1231, new_n1232,
    new_n1233;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT64), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT64), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(new_n464), .A3(G137), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n470), .A2(new_n472), .A3(G125), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n470), .A2(new_n472), .A3(KEYINPUT65), .A4(G125), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n463), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n469), .B1(new_n478), .B2(new_n479), .ZN(G160));
  NAND2_X1  g055(.A1(new_n470), .A2(new_n472), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n463), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OAI221_X1 g058(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n463), .C2(G112), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n481), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND2_X1  g063(.A1(G114), .A2(G2104), .ZN(new_n489));
  INV_X1    g064(.A(G126), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n489), .B1(new_n481), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n463), .A2(new_n464), .A3(G138), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n467), .A2(G102), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT4), .A4(G138), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n492), .A2(new_n495), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n500));
  OR2_X1    g075(.A1(KEYINPUT66), .A2(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT66), .A2(G651), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(G50), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT67), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NOR3_X1   g089(.A1(new_n503), .A2(new_n514), .A3(new_n505), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G88), .ZN(new_n516));
  INV_X1    g091(.A(G75), .ZN(new_n517));
  OR3_X1    g092(.A1(new_n517), .A2(new_n510), .A3(KEYINPUT68), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT68), .B1(new_n517), .B2(new_n510), .ZN(new_n519));
  INV_X1    g094(.A(G62), .ZN(new_n520));
  OAI211_X1 g095(.A(new_n518), .B(new_n519), .C1(new_n520), .C2(new_n514), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT66), .B(G651), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT67), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n506), .A2(new_n525), .A3(new_n507), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n509), .A2(new_n516), .A3(new_n524), .A4(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  INV_X1    g103(.A(G63), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n514), .A2(KEYINPUT69), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT69), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n511), .A2(new_n513), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n529), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(G76), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT7), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g111(.A(G651), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n515), .A2(G89), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n522), .A2(KEYINPUT6), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT70), .ZN(new_n541));
  INV_X1    g116(.A(new_n505), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g118(.A(KEYINPUT70), .B1(new_n503), .B2(new_n505), .ZN(new_n544));
  XNOR2_X1  g119(.A(KEYINPUT71), .B(G51), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n543), .A2(new_n544), .A3(G543), .A4(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n537), .A2(new_n539), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g124(.A1(new_n537), .A2(new_n539), .A3(new_n546), .A4(KEYINPUT72), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(G168));
  NAND2_X1  g126(.A1(new_n530), .A2(new_n532), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n552), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n522), .ZN(new_n554));
  AND3_X1   g129(.A1(new_n543), .A2(new_n544), .A3(G543), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G52), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n515), .A2(G90), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(G301));
  INV_X1    g133(.A(G301), .ZN(G171));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n560));
  NAND2_X1  g135(.A1(G68), .A2(G543), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n530), .A2(new_n532), .ZN(new_n562));
  INV_X1    g137(.A(G56), .ZN(new_n563));
  OAI211_X1 g138(.A(new_n560), .B(new_n561), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n563), .B1(new_n530), .B2(new_n532), .ZN(new_n565));
  INV_X1    g140(.A(new_n561), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT73), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AND3_X1   g142(.A1(new_n564), .A2(new_n567), .A3(new_n523), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n515), .A2(G81), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n543), .A2(new_n544), .A3(G543), .ZN(new_n570));
  INV_X1    g145(.A(G43), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G860), .ZN(G153));
  AND3_X1   g149(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G36), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT74), .ZN(G176));
  NAND2_X1  g152(.A1(G1), .A2(G3), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT8), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n575), .A2(new_n579), .ZN(G188));
  NAND2_X1  g155(.A1(G78), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G65), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n514), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G651), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n583), .A2(KEYINPUT75), .A3(G651), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n586), .A2(new_n587), .B1(new_n515), .B2(G91), .ZN(new_n588));
  INV_X1    g163(.A(G53), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT9), .B1(new_n570), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  NOR3_X1   g166(.A1(new_n570), .A2(KEYINPUT9), .A3(new_n589), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n588), .B1(new_n591), .B2(new_n592), .ZN(G299));
  INV_X1    g168(.A(G168), .ZN(G286));
  NAND2_X1  g169(.A1(new_n555), .A2(G49), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n552), .B2(G74), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n515), .A2(G87), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G288));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G61), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n514), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(new_n523), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(KEYINPUT76), .ZN(new_n603));
  NAND2_X1  g178(.A1(G48), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G86), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n514), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n506), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT76), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n601), .A2(new_n608), .A3(new_n523), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n603), .A2(new_n607), .A3(new_n609), .ZN(G305));
  NAND2_X1  g185(.A1(G72), .A2(G543), .ZN(new_n611));
  INV_X1    g186(.A(G60), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n562), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(new_n523), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n555), .A2(G47), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n515), .A2(G85), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(G290));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  OR3_X1    g193(.A1(G171), .A2(KEYINPUT77), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(KEYINPUT77), .B1(G171), .B2(new_n618), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT78), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n570), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g197(.A1(new_n543), .A2(new_n544), .A3(KEYINPUT78), .A4(G543), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n622), .A2(G54), .A3(new_n623), .ZN(new_n624));
  AND2_X1   g199(.A1(new_n511), .A2(new_n513), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n506), .A2(G92), .A3(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT10), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n625), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(new_n504), .ZN(new_n630));
  AND3_X1   g205(.A1(new_n624), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n619), .B(new_n620), .C1(G868), .C2(new_n631), .ZN(G284));
  OAI211_X1 g207(.A(new_n619), .B(new_n620), .C1(G868), .C2(new_n631), .ZN(G321));
  NAND2_X1  g208(.A1(G299), .A2(new_n618), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n618), .B2(G168), .ZN(G297));
  OAI21_X1  g210(.A(new_n634), .B1(new_n618), .B2(G168), .ZN(G280));
  INV_X1    g211(.A(G559), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n631), .B1(new_n637), .B2(G860), .ZN(G148));
  NAND2_X1  g213(.A1(new_n631), .A2(new_n637), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G868), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(G868), .B2(new_n573), .ZN(G323));
  XNOR2_X1  g216(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g217(.A1(G123), .A2(new_n482), .B1(new_n485), .B2(G135), .ZN(new_n643));
  OAI221_X1 g218(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n463), .C2(G111), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT80), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2096), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n464), .A2(new_n467), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT12), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2100), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n650), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n647), .A2(new_n653), .A3(new_n654), .ZN(G156));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT15), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n660), .A2(G2435), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(G2435), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(KEYINPUT14), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2443), .B(G2446), .Z(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2451), .B(G2454), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n663), .A2(new_n664), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n665), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n668), .B1(new_n665), .B2(new_n669), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n657), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n672), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n674), .A2(new_n670), .A3(new_n656), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n673), .A2(new_n675), .A3(G14), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G401));
  XOR2_X1   g252(.A(G2072), .B(G2078), .Z(new_n678));
  XOR2_X1   g253(.A(G2067), .B(G2678), .Z(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G2084), .B(G2090), .Z(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n678), .B1(new_n682), .B2(KEYINPUT18), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G2096), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G2100), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n682), .A2(KEYINPUT17), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n680), .A2(new_n681), .ZN(new_n687));
  AOI21_X1  g262(.A(KEYINPUT18), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n685), .B(new_n688), .Z(G227));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1971), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT19), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n690), .A2(new_n691), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT20), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n693), .A2(new_n695), .A3(new_n697), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n700), .B(new_n701), .C1(new_n699), .C2(new_n698), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1991), .B(G1996), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1981), .ZN(new_n706));
  INV_X1    g281(.A(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n704), .B(new_n708), .ZN(G229));
  INV_X1    g284(.A(KEYINPUT99), .ZN(new_n710));
  INV_X1    g285(.A(G2072), .ZN(new_n711));
  NOR2_X1   g286(.A1(G29), .A2(G33), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT90), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT25), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT91), .Z(new_n718));
  AOI22_X1  g293(.A1(new_n718), .A2(new_n479), .B1(G139), .B2(new_n485), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT92), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n716), .A2(new_n719), .A3(KEYINPUT92), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n711), .B(new_n713), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n725), .B1(new_n722), .B2(new_n723), .ZN(new_n727));
  OAI21_X1  g302(.A(G2072), .B1(new_n727), .B2(new_n712), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n730), .A2(G5), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G301), .B2(G16), .ZN(new_n732));
  INV_X1    g307(.A(G1961), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT30), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n725), .B1(new_n735), .B2(G28), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT96), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n735), .B2(G28), .ZN(new_n738));
  AOI22_X1  g313(.A1(G129), .A2(new_n482), .B1(new_n485), .B2(G141), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n467), .A2(G105), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT26), .Z(new_n742));
  NAND3_X1  g317(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G29), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G29), .B2(G32), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT27), .B(G1996), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n738), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AND2_X1   g323(.A1(KEYINPUT82), .A2(G29), .ZN(new_n749));
  NOR2_X1   g324(.A1(KEYINPUT82), .A2(G29), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT24), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(G34), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(KEYINPUT93), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(G34), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT93), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n751), .B(new_n756), .C1(new_n752), .C2(G34), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(KEYINPUT94), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(KEYINPUT94), .ZN(new_n760));
  NAND2_X1  g335(.A1(G160), .A2(G29), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G2084), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n748), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT31), .B(G11), .Z(new_n767));
  NOR3_X1   g342(.A1(new_n734), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(G168), .A2(G16), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G16), .B2(G21), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(KEYINPUT95), .ZN(new_n771));
  INV_X1    g346(.A(G1966), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT95), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n769), .B(new_n773), .C1(G16), .C2(G21), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n771), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  AND3_X1   g350(.A1(new_n729), .A2(new_n768), .A3(new_n775), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n746), .A2(new_n747), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n751), .A2(G27), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G164), .B2(new_n751), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT97), .B(G2078), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT98), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n779), .B(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n772), .B1(new_n771), .B2(new_n774), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n776), .A2(new_n777), .A3(new_n782), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n646), .A2(new_n751), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n710), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n729), .A2(new_n775), .A3(new_n768), .ZN(new_n788));
  INV_X1    g363(.A(new_n782), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n788), .A2(new_n789), .A3(new_n783), .ZN(new_n790));
  INV_X1    g365(.A(new_n786), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n790), .A2(KEYINPUT99), .A3(new_n791), .A4(new_n777), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  OR2_X1    g368(.A1(G16), .A2(G22), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G303), .B2(new_n730), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1971), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n730), .A2(G6), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G305), .B2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT32), .B(G1981), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT33), .B(G1976), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n730), .A2(G23), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G288), .B2(G16), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(KEYINPUT84), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT84), .ZN(new_n808));
  AOI211_X1 g383(.A(new_n808), .B(new_n805), .C1(G288), .C2(G16), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n804), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n806), .A2(KEYINPUT84), .ZN(new_n812));
  NOR3_X1   g387(.A1(new_n812), .A2(new_n809), .A3(new_n803), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n802), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n814), .A2(KEYINPUT85), .A3(KEYINPUT34), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT85), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n807), .A2(new_n810), .A3(new_n804), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n803), .B1(new_n812), .B2(new_n809), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n801), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT34), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n816), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n815), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n751), .A2(G25), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n482), .A2(G119), .ZN(new_n824));
  OAI221_X1 g399(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n463), .C2(G107), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n485), .A2(G131), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n823), .B1(new_n828), .B2(new_n751), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT83), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT35), .B(G1991), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n830), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT86), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n819), .B2(new_n820), .ZN(new_n835));
  NOR2_X1   g410(.A1(G16), .A2(G24), .ZN(new_n836));
  INV_X1    g411(.A(G290), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n836), .B1(new_n837), .B2(G16), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n707), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n822), .A2(new_n833), .A3(new_n835), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT36), .ZN(new_n841));
  OAI21_X1  g416(.A(KEYINPUT86), .B1(new_n814), .B2(KEYINPUT34), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(new_n821), .B2(new_n815), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT36), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n843), .A2(new_n844), .A3(new_n833), .A4(new_n839), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n751), .A2(G26), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  OAI221_X1 g424(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n463), .C2(G116), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT88), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n482), .A2(G128), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n485), .A2(G140), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT87), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n849), .B1(new_n857), .B2(G29), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(G2067), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n751), .A2(G35), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(G162), .B2(new_n751), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT29), .B(G2090), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(KEYINPUT100), .B(G1956), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n730), .A2(KEYINPUT23), .A3(G20), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT23), .ZN(new_n866));
  INV_X1    g441(.A(G20), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n867), .B2(G16), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n586), .A2(new_n587), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n515), .A2(G91), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OR3_X1    g446(.A1(new_n570), .A2(KEYINPUT9), .A3(new_n589), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n871), .B1(new_n872), .B2(new_n590), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n865), .B(new_n868), .C1(new_n873), .C2(new_n730), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n859), .B(new_n863), .C1(new_n864), .C2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n573), .A2(G16), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(G16), .B2(G19), .ZN(new_n878));
  INV_X1    g453(.A(G1341), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n730), .A2(G4), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(new_n631), .B2(new_n730), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n882), .A2(G1348), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n882), .A2(G1348), .B1(new_n874), .B2(new_n864), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n876), .A2(new_n880), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(new_n879), .B2(new_n878), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n793), .A2(new_n846), .A3(new_n886), .ZN(G311));
  NAND3_X1  g462(.A1(new_n793), .A2(new_n846), .A3(new_n886), .ZN(G150));
  INV_X1    g463(.A(G67), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n889), .B1(new_n530), .B2(new_n532), .ZN(new_n890));
  AND2_X1   g465(.A1(G80), .A2(G543), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n523), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n543), .A2(new_n544), .A3(G55), .A4(G543), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n515), .A2(G93), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(G860), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT102), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT37), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n631), .A2(G559), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT38), .ZN(new_n900));
  INV_X1    g475(.A(new_n572), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n564), .A2(new_n567), .A3(new_n523), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n902), .A3(new_n895), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n895), .B1(new_n901), .B2(new_n902), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n900), .B(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT39), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n909), .B(KEYINPUT101), .Z(new_n910));
  INV_X1    g485(.A(G860), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(new_n907), .B2(new_n908), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n898), .B1(new_n910), .B2(new_n912), .ZN(G145));
  XNOR2_X1  g488(.A(new_n646), .B(G160), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(new_n487), .ZN(new_n915));
  AOI22_X1  g490(.A1(G130), .A2(new_n482), .B1(new_n485), .B2(G142), .ZN(new_n916));
  OAI221_X1 g491(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n463), .C2(G118), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n828), .B(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT103), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n918), .B(new_n827), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(new_n650), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n854), .A2(new_n498), .A3(new_n856), .ZN(new_n926));
  INV_X1    g501(.A(new_n856), .ZN(new_n927));
  OAI21_X1  g502(.A(G164), .B1(new_n853), .B2(new_n927), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n926), .A2(new_n744), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n744), .B1(new_n926), .B2(new_n928), .ZN(new_n930));
  OR3_X1    g505(.A1(new_n929), .A2(new_n930), .A3(new_n720), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n724), .B1(new_n929), .B2(new_n930), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n925), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n915), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n924), .B(new_n649), .ZN(new_n936));
  INV_X1    g511(.A(new_n932), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n929), .A2(new_n930), .A3(new_n720), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n931), .A2(new_n925), .A3(new_n932), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(KEYINPUT104), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(G37), .B1(new_n935), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n939), .A2(new_n940), .A3(new_n915), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g520(.A(G303), .B(G305), .Z(new_n946));
  AND3_X1   g521(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(G290), .ZN(new_n948));
  NAND4_X1  g523(.A1(G288), .A2(new_n615), .A3(new_n614), .A4(new_n616), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n950), .B1(new_n948), .B2(new_n949), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n946), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OR2_X1    g528(.A1(new_n952), .A2(new_n946), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n955), .B1(new_n956), .B2(KEYINPUT42), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n906), .B(new_n639), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT41), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n631), .A2(G299), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n624), .A2(new_n628), .A3(new_n630), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n873), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n960), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n631), .A2(G299), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n873), .A2(new_n962), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(KEYINPUT41), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n959), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT105), .B1(new_n965), .B2(new_n966), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n965), .A2(KEYINPUT105), .A3(new_n966), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n959), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n958), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n956), .A2(KEYINPUT42), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n957), .A2(new_n969), .A3(new_n972), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n975), .B1(new_n974), .B2(new_n976), .ZN(new_n978));
  OAI21_X1  g553(.A(G868), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n895), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n979), .B1(G868), .B2(new_n980), .ZN(G295));
  OAI21_X1  g556(.A(new_n979), .B1(G868), .B2(new_n980), .ZN(G331));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n980), .B1(new_n568), .B2(new_n572), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n984), .A2(G168), .A3(new_n903), .ZN(new_n985));
  AOI21_X1  g560(.A(G168), .B1(new_n984), .B2(new_n903), .ZN(new_n986));
  OAI21_X1  g561(.A(G301), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(G286), .B1(new_n904), .B2(new_n905), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n984), .A2(G168), .A3(new_n903), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(G171), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n971), .A2(new_n970), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n983), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n968), .A2(new_n990), .A3(new_n987), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n991), .A2(new_n983), .A3(new_n992), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n955), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n965), .A2(new_n966), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n985), .A2(new_n986), .A3(G301), .ZN(new_n1002));
  AOI21_X1  g577(.A(G171), .B1(new_n988), .B2(new_n989), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(new_n994), .A3(new_n955), .ZN(new_n1005));
  INV_X1    g580(.A(G37), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n999), .A2(new_n1000), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n955), .B1(new_n1004), .B2(new_n994), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(KEYINPUT43), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT44), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n997), .A2(new_n993), .A3(new_n995), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1013), .B(new_n1000), .C1(new_n1014), .C2(new_n955), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT43), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT44), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1012), .A2(new_n1019), .ZN(G397));
  XNOR2_X1  g595(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT109), .B(G1384), .Z(new_n1022));
  AOI21_X1  g597(.A(new_n1021), .B1(new_n498), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G40), .ZN(new_n1024));
  AOI211_X1 g599(.A(new_n1024), .B(new_n469), .C1(new_n479), .C2(new_n478), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G2067), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n857), .B(new_n1027), .ZN(new_n1028));
  XOR2_X1   g603(.A(new_n743), .B(G1996), .Z(new_n1029));
  AND2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1030), .A2(new_n832), .A3(new_n828), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n854), .A2(new_n1027), .A3(new_n856), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1026), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1026), .A2(G1996), .ZN(new_n1034));
  OR2_X1    g609(.A1(new_n1034), .A2(KEYINPUT46), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(KEYINPUT46), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1028), .A2(new_n744), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1026), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n1040), .B(KEYINPUT47), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1030), .B1(new_n831), .B2(new_n827), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n828), .A2(new_n832), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1039), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n837), .A2(new_n707), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1045), .A2(new_n1026), .ZN(new_n1046));
  XOR2_X1   g621(.A(new_n1046), .B(KEYINPUT48), .Z(new_n1047));
  AOI211_X1 g622(.A(new_n1033), .B(new_n1041), .C1(new_n1044), .C2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1384), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n495), .A2(new_n497), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n464), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n496), .B1(new_n1051), .B2(new_n459), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1049), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT50), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT50), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n498), .A2(new_n1055), .A3(new_n1049), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1054), .A2(new_n763), .A3(new_n1025), .A4(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT119), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT45), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1053), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n498), .A2(new_n1049), .A3(new_n1021), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1025), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n772), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n478), .A2(new_n479), .ZN(new_n1064));
  INV_X1    g639(.A(new_n469), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(G40), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(KEYINPUT50), .B2(new_n1053), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(new_n763), .A4(new_n1056), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1058), .A2(new_n1063), .A3(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT113), .B(G8), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n549), .A2(new_n550), .A3(new_n1071), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n1073), .A2(KEYINPUT51), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1073), .B1(new_n1070), .B2(G8), .ZN(new_n1075));
  XOR2_X1   g650(.A(KEYINPUT126), .B(KEYINPUT51), .Z(new_n1076));
  OAI22_X1  g651(.A1(new_n1072), .A2(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1072), .A2(G286), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1971), .ZN(new_n1080));
  OAI211_X1 g655(.A(KEYINPUT45), .B(new_n1022), .C1(new_n1050), .C2(new_n1052), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1025), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1021), .B1(new_n498), .B2(new_n1049), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1080), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1054), .A2(KEYINPUT118), .A3(new_n1025), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1055), .B1(new_n498), .B2(new_n1049), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(new_n1087), .B2(new_n1066), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(new_n1088), .A3(new_n1056), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1084), .B1(new_n1089), .B2(G2090), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n1071), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT111), .B(KEYINPUT55), .Z(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1093), .B1(G303), .B2(G8), .ZN(new_n1094));
  AND2_X1   g669(.A1(G303), .A2(G8), .ZN(new_n1095));
  NOR2_X1   g670(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1091), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1100), .B1(new_n1102), .B2(G2078), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1067), .A2(new_n1056), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n733), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(G301), .B(KEYINPUT54), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1023), .ZN(new_n1109));
  INV_X1    g684(.A(G2078), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1110), .A2(KEYINPUT127), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(KEYINPUT127), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1100), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1109), .A2(new_n1025), .A3(new_n1081), .A4(new_n1113), .ZN(new_n1114));
  OR3_X1    g689(.A1(new_n1062), .A2(new_n1100), .A3(G2078), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1103), .A2(new_n1115), .A3(new_n1105), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1108), .A2(new_n1114), .B1(new_n1116), .B2(new_n1107), .ZN(new_n1117));
  OR2_X1    g692(.A1(G305), .A2(G1981), .ZN(new_n1118));
  NAND2_X1  g693(.A1(G305), .A2(G1981), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT114), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(KEYINPUT49), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1053), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n1025), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1125), .A2(new_n1071), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1118), .B(new_n1119), .C1(new_n1121), .C2(KEYINPUT49), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1123), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(G1976), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1125), .B(new_n1071), .C1(G288), .C2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT52), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n947), .A2(G1976), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT52), .B1(G288), .B2(new_n1129), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1126), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1128), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(G2090), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1054), .A2(new_n1136), .A3(new_n1025), .A4(new_n1056), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1084), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1138), .A2(G8), .A3(new_n1097), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT112), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT112), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1138), .A2(new_n1097), .A3(new_n1141), .A4(G8), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1135), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1079), .A2(new_n1099), .A3(new_n1117), .A4(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1124), .A2(new_n1145), .A3(new_n1025), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT122), .B1(new_n1053), .B2(new_n1066), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1146), .A2(new_n1027), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(G1348), .B1(new_n1067), .B2(new_n1056), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n962), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(G1348), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1104), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1146), .A2(new_n1027), .A3(new_n1147), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1152), .A2(new_n631), .A3(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1150), .A2(KEYINPUT60), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1152), .A2(new_n1156), .A3(new_n631), .A4(new_n1153), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT125), .ZN(new_n1159));
  INV_X1    g734(.A(G1956), .ZN(new_n1160));
  XNOR2_X1  g735(.A(KEYINPUT56), .B(G2072), .ZN(new_n1161));
  AOI22_X1  g736(.A1(new_n1089), .A2(new_n1160), .B1(new_n1101), .B2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(G299), .A2(new_n1164), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n588), .B(new_n1163), .C1(new_n591), .C2(new_n592), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1159), .B1(new_n1162), .B2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1162), .A2(new_n1167), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1089), .A2(new_n1160), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1101), .A2(new_n1161), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1171), .A2(new_n1167), .A3(new_n1159), .A4(new_n1172), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n1173), .A2(KEYINPUT61), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1158), .B1(new_n1170), .B2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g750(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n1176));
  AND2_X1   g751(.A1(new_n1162), .A2(new_n1167), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1176), .B1(new_n1177), .B2(new_n1169), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT124), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1180), .B(new_n1176), .C1(new_n1177), .C2(new_n1169), .ZN(new_n1181));
  XNOR2_X1  g756(.A(KEYINPUT58), .B(G1341), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1182), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n1082), .A2(G1996), .A3(new_n1083), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n573), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT59), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1175), .A2(new_n1179), .A3(new_n1181), .A4(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1177), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n962), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1188), .B1(new_n1169), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1144), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1135), .ZN(new_n1193));
  AND3_X1   g768(.A1(new_n1070), .A2(G168), .A3(new_n1071), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1192), .A2(new_n1099), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT63), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1138), .A2(G8), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1196), .B1(new_n1198), .B2(new_n1098), .ZN(new_n1199));
  NAND4_X1  g774(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .A4(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT120), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1143), .A2(KEYINPUT120), .A3(new_n1194), .A4(new_n1199), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1197), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1192), .A2(new_n1135), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1128), .A2(new_n1129), .A3(new_n947), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT117), .ZN(new_n1207));
  XOR2_X1   g782(.A(new_n1118), .B(KEYINPUT116), .Z(new_n1208));
  AND3_X1   g783(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1207), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  XOR2_X1   g786(.A(new_n1126), .B(KEYINPUT115), .Z(new_n1212));
  AOI21_X1  g787(.A(new_n1205), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1204), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1070), .A2(G8), .ZN(new_n1216));
  INV_X1    g791(.A(new_n1073), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1076), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1074), .B1(new_n1071), .B2(new_n1070), .ZN(new_n1219));
  OAI211_X1 g794(.A(new_n1078), .B(new_n1215), .C1(new_n1218), .C2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1220), .A2(G171), .A3(new_n1116), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1143), .A2(new_n1099), .ZN(new_n1222));
  AOI21_X1  g797(.A(new_n1215), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1223));
  NOR3_X1   g798(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  NOR3_X1   g799(.A1(new_n1191), .A2(new_n1214), .A3(new_n1224), .ZN(new_n1225));
  AOI211_X1 g800(.A(new_n1043), .B(new_n1042), .C1(G1986), .C2(G290), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1026), .B1(new_n1226), .B2(new_n1045), .ZN(new_n1227));
  OAI21_X1  g802(.A(new_n1048), .B1(new_n1225), .B2(new_n1227), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g803(.A(G229), .ZN(new_n1230));
  INV_X1    g804(.A(G227), .ZN(new_n1231));
  NAND2_X1  g805(.A1(new_n676), .A2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g806(.A(new_n1232), .B1(new_n942), .B2(new_n943), .ZN(new_n1233));
  AND4_X1   g807(.A1(G319), .A2(new_n1017), .A3(new_n1230), .A4(new_n1233), .ZN(G308));
  NAND4_X1  g808(.A1(new_n1017), .A2(new_n1233), .A3(G319), .A4(new_n1230), .ZN(G225));
endmodule


