

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X2 U549 ( .A1(n829), .A2(n831), .ZN(n740) );
  NAND2_X2 U550 ( .A1(n535), .A2(n532), .ZN(n897) );
  XNOR2_X1 U551 ( .A(n745), .B(n523), .ZN(n748) );
  INV_X1 U552 ( .A(KEYINPUT95), .ZN(n523) );
  XNOR2_X1 U553 ( .A(n522), .B(n746), .ZN(n521) );
  INV_X1 U554 ( .A(KEYINPUT97), .ZN(n746) );
  NOR2_X1 U555 ( .A1(n748), .A2(G299), .ZN(n522) );
  XNOR2_X1 U556 ( .A(KEYINPUT29), .B(KEYINPUT98), .ZN(n753) );
  NOR2_X1 U557 ( .A1(n723), .A2(G1966), .ZN(n770) );
  NOR2_X1 U558 ( .A1(G2104), .A2(KEYINPUT17), .ZN(n536) );
  NAND2_X1 U559 ( .A1(G2105), .A2(KEYINPUT17), .ZN(n533) );
  INV_X1 U560 ( .A(KEYINPUT104), .ZN(n782) );
  NAND2_X1 U561 ( .A1(n515), .A2(n531), .ZN(n530) );
  INV_X1 U562 ( .A(n978), .ZN(n531) );
  NOR2_X1 U563 ( .A1(n740), .A2(n954), .ZN(n742) );
  NOR2_X1 U564 ( .A1(n752), .A2(n751), .ZN(n754) );
  NOR2_X1 U565 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U566 ( .A(n538), .B(n537), .ZN(n829) );
  INV_X1 U567 ( .A(KEYINPUT64), .ZN(n537) );
  NOR2_X1 U568 ( .A1(G164), .A2(G1384), .ZN(n538) );
  XNOR2_X1 U569 ( .A(n526), .B(KEYINPUT103), .ZN(n525) );
  INV_X1 U570 ( .A(KEYINPUT33), .ZN(n524) );
  AND2_X1 U571 ( .A1(n534), .A2(n533), .ZN(n532) );
  NAND2_X1 U572 ( .A1(n536), .A2(n580), .ZN(n535) );
  NAND2_X1 U573 ( .A1(G2104), .A2(KEYINPUT17), .ZN(n534) );
  XNOR2_X1 U574 ( .A(KEYINPUT65), .B(KEYINPUT23), .ZN(n587) );
  NAND2_X1 U575 ( .A1(n518), .A2(n515), .ZN(n527) );
  OR2_X1 U576 ( .A1(n529), .A2(n530), .ZN(n528) );
  OR2_X1 U577 ( .A1(n841), .A2(n840), .ZN(n515) );
  XOR2_X1 U578 ( .A(KEYINPUT75), .B(n559), .Z(n516) );
  XNOR2_X1 U579 ( .A(KEYINPUT87), .B(n584), .ZN(n517) );
  OR2_X1 U580 ( .A1(n834), .A2(n540), .ZN(n518) );
  NOR2_X1 U581 ( .A1(n770), .A2(n769), .ZN(n519) );
  AND2_X1 U582 ( .A1(n585), .A2(n539), .ZN(G164) );
  AND2_X1 U583 ( .A1(n790), .A2(n524), .ZN(n520) );
  NOR2_X1 U584 ( .A1(n747), .A2(n521), .ZN(n752) );
  NAND2_X1 U585 ( .A1(n525), .A2(n520), .ZN(n781) );
  NAND2_X1 U586 ( .A1(n778), .A2(n986), .ZN(n526) );
  NAND2_X1 U587 ( .A1(n528), .A2(n527), .ZN(n842) );
  XNOR2_X1 U588 ( .A(n783), .B(n782), .ZN(n529) );
  NAND2_X1 U589 ( .A1(n897), .A2(G138), .ZN(n583) );
  NOR2_X1 U590 ( .A1(n586), .A2(n517), .ZN(n539) );
  AND2_X2 U591 ( .A1(G2105), .A2(G2104), .ZN(n894) );
  AND2_X2 U592 ( .A1(n580), .A2(G2104), .ZN(n898) );
  NAND2_X1 U593 ( .A1(n833), .A2(n835), .ZN(n540) );
  XNOR2_X1 U594 ( .A(n774), .B(KEYINPUT102), .ZN(n784) );
  INV_X1 U595 ( .A(G8), .ZN(n711) );
  OR2_X1 U596 ( .A1(n768), .A2(n711), .ZN(n712) );
  INV_X1 U597 ( .A(KEYINPUT30), .ZN(n713) );
  XNOR2_X1 U598 ( .A(n714), .B(n713), .ZN(n715) );
  INV_X1 U599 ( .A(KEYINPUT32), .ZN(n764) );
  NOR2_X1 U600 ( .A1(G543), .A2(n544), .ZN(n541) );
  NOR2_X1 U601 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U602 ( .A(n588), .B(n587), .ZN(n591) );
  NOR2_X1 U603 ( .A1(G651), .A2(n649), .ZN(n670) );
  INV_X1 U604 ( .A(KEYINPUT8), .ZN(n560) );
  NOR2_X1 U605 ( .A1(G651), .A2(G543), .ZN(n669) );
  NAND2_X1 U606 ( .A1(n669), .A2(G91), .ZN(n543) );
  XOR2_X1 U607 ( .A(G651), .B(KEYINPUT68), .Z(n544) );
  XOR2_X2 U608 ( .A(KEYINPUT1), .B(n541), .Z(n677) );
  NAND2_X1 U609 ( .A1(G65), .A2(n677), .ZN(n542) );
  NAND2_X1 U610 ( .A1(n543), .A2(n542), .ZN(n548) );
  XOR2_X1 U611 ( .A(G543), .B(KEYINPUT0), .Z(n649) );
  NAND2_X1 U612 ( .A1(n670), .A2(G53), .ZN(n546) );
  NOR2_X1 U613 ( .A1(n649), .A2(n544), .ZN(n673) );
  NAND2_X1 U614 ( .A1(G78), .A2(n673), .ZN(n545) );
  NAND2_X1 U615 ( .A1(n546), .A2(n545), .ZN(n547) );
  OR2_X1 U616 ( .A1(n548), .A2(n547), .ZN(G299) );
  NAND2_X1 U617 ( .A1(G63), .A2(n677), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n549), .B(KEYINPUT74), .ZN(n551) );
  NAND2_X1 U619 ( .A1(G51), .A2(n670), .ZN(n550) );
  NAND2_X1 U620 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U621 ( .A(KEYINPUT6), .B(n552), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n669), .A2(G89), .ZN(n553) );
  XNOR2_X1 U623 ( .A(n553), .B(KEYINPUT4), .ZN(n555) );
  NAND2_X1 U624 ( .A1(G76), .A2(n673), .ZN(n554) );
  NAND2_X1 U625 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U626 ( .A(n556), .B(KEYINPUT5), .Z(n557) );
  XOR2_X1 U627 ( .A(KEYINPUT7), .B(n516), .Z(G168) );
  XNOR2_X1 U628 ( .A(G168), .B(n560), .ZN(G286) );
  XNOR2_X1 U629 ( .A(G2454), .B(G2443), .ZN(n570) );
  XOR2_X1 U630 ( .A(KEYINPUT108), .B(G2430), .Z(n562) );
  XNOR2_X1 U631 ( .A(G2446), .B(KEYINPUT109), .ZN(n561) );
  XNOR2_X1 U632 ( .A(n562), .B(n561), .ZN(n566) );
  XOR2_X1 U633 ( .A(G2451), .B(G2427), .Z(n564) );
  XNOR2_X1 U634 ( .A(G1341), .B(G1348), .ZN(n563) );
  XNOR2_X1 U635 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U636 ( .A(n566), .B(n565), .Z(n568) );
  XNOR2_X1 U637 ( .A(G2435), .B(G2438), .ZN(n567) );
  XNOR2_X1 U638 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U639 ( .A(n570), .B(n569), .ZN(n571) );
  AND2_X1 U640 ( .A1(n571), .A2(G14), .ZN(G401) );
  NAND2_X1 U641 ( .A1(n670), .A2(G52), .ZN(n573) );
  NAND2_X1 U642 ( .A1(G64), .A2(n677), .ZN(n572) );
  NAND2_X1 U643 ( .A1(n573), .A2(n572), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n669), .A2(G90), .ZN(n574) );
  XOR2_X1 U645 ( .A(KEYINPUT69), .B(n574), .Z(n576) );
  NAND2_X1 U646 ( .A1(G77), .A2(n673), .ZN(n575) );
  NAND2_X1 U647 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U648 ( .A(KEYINPUT9), .B(n577), .Z(n578) );
  NOR2_X1 U649 ( .A1(n579), .A2(n578), .ZN(G171) );
  AND2_X1 U650 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U651 ( .A(G2105), .ZN(n580) );
  NOR2_X2 U652 ( .A1(G2104), .A2(n580), .ZN(n893) );
  NAND2_X1 U653 ( .A1(G126), .A2(n893), .ZN(n582) );
  NAND2_X1 U654 ( .A1(G102), .A2(n898), .ZN(n581) );
  NAND2_X1 U655 ( .A1(n582), .A2(n581), .ZN(n586) );
  XNOR2_X1 U656 ( .A(n583), .B(KEYINPUT88), .ZN(n585) );
  NAND2_X1 U657 ( .A1(G114), .A2(n894), .ZN(n584) );
  NAND2_X1 U658 ( .A1(G101), .A2(n898), .ZN(n588) );
  NAND2_X1 U659 ( .A1(G113), .A2(n894), .ZN(n589) );
  XNOR2_X1 U660 ( .A(n589), .B(KEYINPUT66), .ZN(n590) );
  NAND2_X1 U661 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U662 ( .A1(G125), .A2(n893), .ZN(n593) );
  NAND2_X1 U663 ( .A1(G137), .A2(n897), .ZN(n592) );
  NAND2_X1 U664 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U665 ( .A1(n595), .A2(n594), .ZN(G160) );
  INV_X1 U666 ( .A(G57), .ZN(G237) );
  NAND2_X1 U667 ( .A1(G7), .A2(G661), .ZN(n596) );
  XNOR2_X1 U668 ( .A(n596), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U669 ( .A(G223), .ZN(n843) );
  NAND2_X1 U670 ( .A1(n843), .A2(G567), .ZN(n597) );
  XOR2_X1 U671 ( .A(KEYINPUT11), .B(n597), .Z(G234) );
  NAND2_X1 U672 ( .A1(G56), .A2(n677), .ZN(n598) );
  XNOR2_X1 U673 ( .A(KEYINPUT14), .B(n598), .ZN(n605) );
  NAND2_X1 U674 ( .A1(G68), .A2(n673), .ZN(n599) );
  XNOR2_X1 U675 ( .A(KEYINPUT70), .B(n599), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n669), .A2(G81), .ZN(n600) );
  XNOR2_X1 U677 ( .A(KEYINPUT12), .B(n600), .ZN(n601) );
  NAND2_X1 U678 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U679 ( .A(KEYINPUT13), .B(n603), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U681 ( .A(n606), .B(KEYINPUT71), .ZN(n608) );
  NAND2_X1 U682 ( .A1(G43), .A2(n670), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n994) );
  INV_X1 U684 ( .A(G860), .ZN(n623) );
  OR2_X1 U685 ( .A1(n994), .A2(n623), .ZN(G153) );
  XOR2_X1 U686 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  NAND2_X1 U687 ( .A1(G868), .A2(G301), .ZN(n618) );
  NAND2_X1 U688 ( .A1(n670), .A2(G54), .ZN(n615) );
  NAND2_X1 U689 ( .A1(G66), .A2(n677), .ZN(n610) );
  NAND2_X1 U690 ( .A1(G79), .A2(n673), .ZN(n609) );
  NAND2_X1 U691 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U692 ( .A1(G92), .A2(n669), .ZN(n611) );
  XNOR2_X1 U693 ( .A(KEYINPUT73), .B(n611), .ZN(n612) );
  NOR2_X1 U694 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U696 ( .A(KEYINPUT15), .B(n616), .Z(n980) );
  INV_X1 U697 ( .A(G868), .ZN(n619) );
  NAND2_X1 U698 ( .A1(n980), .A2(n619), .ZN(n617) );
  NAND2_X1 U699 ( .A1(n618), .A2(n617), .ZN(G284) );
  NOR2_X1 U700 ( .A1(G286), .A2(n619), .ZN(n621) );
  NOR2_X1 U701 ( .A1(G868), .A2(G299), .ZN(n620) );
  NOR2_X1 U702 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U703 ( .A(KEYINPUT76), .B(n622), .ZN(G297) );
  NAND2_X1 U704 ( .A1(n623), .A2(G559), .ZN(n624) );
  INV_X1 U705 ( .A(n980), .ZN(n913) );
  NAND2_X1 U706 ( .A1(n624), .A2(n913), .ZN(n625) );
  XNOR2_X1 U707 ( .A(n625), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U708 ( .A1(G868), .A2(n994), .ZN(n628) );
  NAND2_X1 U709 ( .A1(G868), .A2(n913), .ZN(n626) );
  NOR2_X1 U710 ( .A1(G559), .A2(n626), .ZN(n627) );
  NOR2_X1 U711 ( .A1(n628), .A2(n627), .ZN(G282) );
  NAND2_X1 U712 ( .A1(n893), .A2(G123), .ZN(n629) );
  XNOR2_X1 U713 ( .A(n629), .B(KEYINPUT18), .ZN(n631) );
  NAND2_X1 U714 ( .A1(G135), .A2(n897), .ZN(n630) );
  NAND2_X1 U715 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U716 ( .A(n632), .B(KEYINPUT77), .ZN(n634) );
  NAND2_X1 U717 ( .A1(G111), .A2(n894), .ZN(n633) );
  NAND2_X1 U718 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n898), .A2(G99), .ZN(n635) );
  XOR2_X1 U720 ( .A(KEYINPUT78), .B(n635), .Z(n636) );
  NOR2_X1 U721 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U722 ( .A(KEYINPUT79), .B(n638), .Z(n936) );
  XNOR2_X1 U723 ( .A(n936), .B(G2096), .ZN(n640) );
  INV_X1 U724 ( .A(G2100), .ZN(n639) );
  NAND2_X1 U725 ( .A1(n640), .A2(n639), .ZN(G156) );
  NAND2_X1 U726 ( .A1(G559), .A2(n913), .ZN(n641) );
  XNOR2_X1 U727 ( .A(n994), .B(n641), .ZN(n688) );
  NOR2_X1 U728 ( .A1(n688), .A2(G860), .ZN(n648) );
  NAND2_X1 U729 ( .A1(n670), .A2(G55), .ZN(n643) );
  NAND2_X1 U730 ( .A1(G67), .A2(n677), .ZN(n642) );
  NAND2_X1 U731 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U732 ( .A1(G93), .A2(n669), .ZN(n645) );
  NAND2_X1 U733 ( .A1(G80), .A2(n673), .ZN(n644) );
  NAND2_X1 U734 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U735 ( .A1(n647), .A2(n646), .ZN(n683) );
  XNOR2_X1 U736 ( .A(n648), .B(n683), .ZN(G145) );
  NAND2_X1 U737 ( .A1(G87), .A2(n649), .ZN(n651) );
  NAND2_X1 U738 ( .A1(G74), .A2(G651), .ZN(n650) );
  NAND2_X1 U739 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U740 ( .A1(n677), .A2(n652), .ZN(n654) );
  NAND2_X1 U741 ( .A1(n670), .A2(G49), .ZN(n653) );
  NAND2_X1 U742 ( .A1(n654), .A2(n653), .ZN(G288) );
  NAND2_X1 U743 ( .A1(G60), .A2(n677), .ZN(n656) );
  NAND2_X1 U744 ( .A1(G72), .A2(n673), .ZN(n655) );
  NAND2_X1 U745 ( .A1(n656), .A2(n655), .ZN(n659) );
  NAND2_X1 U746 ( .A1(G85), .A2(n669), .ZN(n657) );
  XNOR2_X1 U747 ( .A(KEYINPUT67), .B(n657), .ZN(n658) );
  NOR2_X1 U748 ( .A1(n659), .A2(n658), .ZN(n661) );
  NAND2_X1 U749 ( .A1(n670), .A2(G47), .ZN(n660) );
  NAND2_X1 U750 ( .A1(n661), .A2(n660), .ZN(G290) );
  NAND2_X1 U751 ( .A1(G88), .A2(n669), .ZN(n663) );
  NAND2_X1 U752 ( .A1(G75), .A2(n673), .ZN(n662) );
  NAND2_X1 U753 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U754 ( .A(KEYINPUT80), .B(n664), .Z(n668) );
  NAND2_X1 U755 ( .A1(n677), .A2(G62), .ZN(n666) );
  NAND2_X1 U756 ( .A1(n670), .A2(G50), .ZN(n665) );
  AND2_X1 U757 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U758 ( .A1(n668), .A2(n667), .ZN(G303) );
  NAND2_X1 U759 ( .A1(G86), .A2(n669), .ZN(n672) );
  NAND2_X1 U760 ( .A1(G48), .A2(n670), .ZN(n671) );
  NAND2_X1 U761 ( .A1(n672), .A2(n671), .ZN(n676) );
  NAND2_X1 U762 ( .A1(n673), .A2(G73), .ZN(n674) );
  XOR2_X1 U763 ( .A(KEYINPUT2), .B(n674), .Z(n675) );
  NOR2_X1 U764 ( .A1(n676), .A2(n675), .ZN(n679) );
  NAND2_X1 U765 ( .A1(G61), .A2(n677), .ZN(n678) );
  NAND2_X1 U766 ( .A1(n679), .A2(n678), .ZN(G305) );
  NOR2_X1 U767 ( .A1(n683), .A2(G868), .ZN(n680) );
  XNOR2_X1 U768 ( .A(KEYINPUT83), .B(n680), .ZN(n692) );
  XNOR2_X1 U769 ( .A(KEYINPUT81), .B(G299), .ZN(n681) );
  XNOR2_X1 U770 ( .A(n681), .B(G288), .ZN(n682) );
  XNOR2_X1 U771 ( .A(KEYINPUT19), .B(n682), .ZN(n685) );
  XNOR2_X1 U772 ( .A(G290), .B(n683), .ZN(n684) );
  XNOR2_X1 U773 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U774 ( .A(n686), .B(G303), .ZN(n687) );
  XNOR2_X1 U775 ( .A(n687), .B(G305), .ZN(n916) );
  XOR2_X1 U776 ( .A(n916), .B(n688), .Z(n689) );
  NAND2_X1 U777 ( .A1(n689), .A2(G868), .ZN(n690) );
  XNOR2_X1 U778 ( .A(KEYINPUT82), .B(n690), .ZN(n691) );
  NAND2_X1 U779 ( .A1(n692), .A2(n691), .ZN(G295) );
  NAND2_X1 U780 ( .A1(G2084), .A2(G2078), .ZN(n693) );
  XOR2_X1 U781 ( .A(KEYINPUT20), .B(n693), .Z(n694) );
  NAND2_X1 U782 ( .A1(G2090), .A2(n694), .ZN(n695) );
  XNOR2_X1 U783 ( .A(KEYINPUT21), .B(n695), .ZN(n696) );
  NAND2_X1 U784 ( .A1(n696), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U785 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U786 ( .A1(G120), .A2(G69), .ZN(n697) );
  NOR2_X1 U787 ( .A1(G237), .A2(n697), .ZN(n698) );
  XNOR2_X1 U788 ( .A(KEYINPUT86), .B(n698), .ZN(n699) );
  NAND2_X1 U789 ( .A1(n699), .A2(G108), .ZN(n847) );
  NAND2_X1 U790 ( .A1(n847), .A2(G567), .ZN(n706) );
  NAND2_X1 U791 ( .A1(G132), .A2(G82), .ZN(n700) );
  XNOR2_X1 U792 ( .A(n700), .B(KEYINPUT22), .ZN(n701) );
  XNOR2_X1 U793 ( .A(n701), .B(KEYINPUT84), .ZN(n702) );
  NOR2_X1 U794 ( .A1(G218), .A2(n702), .ZN(n703) );
  XOR2_X1 U795 ( .A(KEYINPUT85), .B(n703), .Z(n704) );
  NAND2_X1 U796 ( .A1(G96), .A2(n704), .ZN(n848) );
  NAND2_X1 U797 ( .A1(n848), .A2(G2106), .ZN(n705) );
  NAND2_X1 U798 ( .A1(n706), .A2(n705), .ZN(n849) );
  NAND2_X1 U799 ( .A1(G661), .A2(G483), .ZN(n707) );
  NOR2_X1 U800 ( .A1(n849), .A2(n707), .ZN(n846) );
  NAND2_X1 U801 ( .A1(n846), .A2(G36), .ZN(G176) );
  INV_X1 U802 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U803 ( .A(G1981), .B(G305), .ZN(n978) );
  NAND2_X1 U804 ( .A1(G160), .A2(G40), .ZN(n831) );
  NAND2_X1 U805 ( .A1(n740), .A2(G8), .ZN(n710) );
  XOR2_X2 U806 ( .A(KEYINPUT92), .B(n710), .Z(n790) );
  INV_X1 U807 ( .A(n790), .ZN(n723) );
  NOR2_X1 U808 ( .A1(G2084), .A2(n740), .ZN(n768) );
  NOR2_X1 U809 ( .A1(n770), .A2(n712), .ZN(n714) );
  NOR2_X1 U810 ( .A1(G168), .A2(n715), .ZN(n719) );
  XNOR2_X1 U811 ( .A(G1961), .B(KEYINPUT93), .ZN(n1001) );
  NAND2_X1 U812 ( .A1(n740), .A2(n1001), .ZN(n717) );
  INV_X1 U813 ( .A(n740), .ZN(n728) );
  XNOR2_X1 U814 ( .A(G2078), .B(KEYINPUT25), .ZN(n964) );
  NAND2_X1 U815 ( .A1(n728), .A2(n964), .ZN(n716) );
  NAND2_X1 U816 ( .A1(n717), .A2(n716), .ZN(n755) );
  NOR2_X1 U817 ( .A1(G171), .A2(n755), .ZN(n718) );
  NOR2_X1 U818 ( .A1(n719), .A2(n718), .ZN(n722) );
  XNOR2_X1 U819 ( .A(KEYINPUT31), .B(KEYINPUT99), .ZN(n720) );
  XNOR2_X1 U820 ( .A(n720), .B(KEYINPUT100), .ZN(n721) );
  XNOR2_X1 U821 ( .A(n722), .B(n721), .ZN(n766) );
  NOR2_X1 U822 ( .A1(n723), .A2(G1971), .ZN(n724) );
  XNOR2_X1 U823 ( .A(KEYINPUT101), .B(n724), .ZN(n727) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n740), .ZN(n725) );
  NOR2_X1 U825 ( .A1(G166), .A2(n725), .ZN(n726) );
  NAND2_X1 U826 ( .A1(n727), .A2(n726), .ZN(n759) );
  AND2_X1 U827 ( .A1(n766), .A2(n759), .ZN(n758) );
  NAND2_X1 U828 ( .A1(G1348), .A2(n740), .ZN(n730) );
  NAND2_X1 U829 ( .A1(G2067), .A2(n728), .ZN(n729) );
  NAND2_X1 U830 ( .A1(n730), .A2(n729), .ZN(n737) );
  NOR2_X1 U831 ( .A1(n980), .A2(n737), .ZN(n736) );
  INV_X1 U832 ( .A(G1996), .ZN(n955) );
  NOR2_X1 U833 ( .A1(n740), .A2(n955), .ZN(n731) );
  XOR2_X1 U834 ( .A(n731), .B(KEYINPUT26), .Z(n733) );
  NAND2_X1 U835 ( .A1(n740), .A2(G1341), .ZN(n732) );
  NAND2_X1 U836 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U837 ( .A1(n734), .A2(n994), .ZN(n735) );
  NOR2_X1 U838 ( .A1(n736), .A2(n735), .ZN(n739) );
  AND2_X1 U839 ( .A1(n980), .A2(n737), .ZN(n738) );
  NOR2_X1 U840 ( .A1(n739), .A2(n738), .ZN(n747) );
  INV_X1 U841 ( .A(G2072), .ZN(n954) );
  XNOR2_X1 U842 ( .A(KEYINPUT27), .B(KEYINPUT94), .ZN(n741) );
  XNOR2_X1 U843 ( .A(n742), .B(n741), .ZN(n744) );
  NAND2_X1 U844 ( .A1(n740), .A2(G1956), .ZN(n743) );
  NAND2_X1 U845 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U846 ( .A(KEYINPUT28), .B(KEYINPUT96), .Z(n750) );
  NAND2_X1 U847 ( .A1(n748), .A2(G299), .ZN(n749) );
  XNOR2_X1 U848 ( .A(n750), .B(n749), .ZN(n751) );
  XNOR2_X1 U849 ( .A(n754), .B(n753), .ZN(n757) );
  NAND2_X1 U850 ( .A1(G171), .A2(n755), .ZN(n756) );
  NAND2_X1 U851 ( .A1(n757), .A2(n756), .ZN(n767) );
  NAND2_X1 U852 ( .A1(n758), .A2(n767), .ZN(n763) );
  INV_X1 U853 ( .A(n759), .ZN(n760) );
  OR2_X1 U854 ( .A1(G286), .A2(n760), .ZN(n761) );
  AND2_X1 U855 ( .A1(n761), .A2(G8), .ZN(n762) );
  NAND2_X1 U856 ( .A1(n763), .A2(n762), .ZN(n765) );
  XNOR2_X1 U857 ( .A(n765), .B(n764), .ZN(n773) );
  NAND2_X1 U858 ( .A1(n766), .A2(n767), .ZN(n771) );
  AND2_X1 U859 ( .A1(G8), .A2(n768), .ZN(n769) );
  AND2_X1 U860 ( .A1(n771), .A2(n519), .ZN(n772) );
  INV_X1 U861 ( .A(n784), .ZN(n777) );
  NOR2_X1 U862 ( .A1(G1971), .A2(G303), .ZN(n775) );
  NOR2_X1 U863 ( .A1(G1976), .A2(G288), .ZN(n983) );
  NOR2_X1 U864 ( .A1(n775), .A2(n983), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U866 ( .A1(G1976), .A2(G288), .ZN(n986) );
  NAND2_X1 U867 ( .A1(n983), .A2(n790), .ZN(n779) );
  NAND2_X1 U868 ( .A1(n779), .A2(KEYINPUT33), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G166), .A2(G8), .ZN(n785) );
  NOR2_X1 U871 ( .A1(G2090), .A2(n785), .ZN(n786) );
  NOR2_X1 U872 ( .A1(n784), .A2(n786), .ZN(n787) );
  XOR2_X1 U873 ( .A(KEYINPUT105), .B(n787), .Z(n788) );
  NOR2_X1 U874 ( .A1(n790), .A2(n788), .ZN(n834) );
  NOR2_X1 U875 ( .A1(G1981), .A2(G305), .ZN(n789) );
  XNOR2_X1 U876 ( .A(n789), .B(KEYINPUT24), .ZN(n791) );
  NAND2_X1 U877 ( .A1(n791), .A2(n790), .ZN(n833) );
  NAND2_X1 U878 ( .A1(G140), .A2(n897), .ZN(n793) );
  NAND2_X1 U879 ( .A1(G104), .A2(n898), .ZN(n792) );
  NAND2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U881 ( .A(KEYINPUT34), .B(n794), .ZN(n799) );
  NAND2_X1 U882 ( .A1(G128), .A2(n893), .ZN(n796) );
  NAND2_X1 U883 ( .A1(G116), .A2(n894), .ZN(n795) );
  NAND2_X1 U884 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U885 ( .A(KEYINPUT35), .B(n797), .Z(n798) );
  NOR2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U887 ( .A(KEYINPUT36), .B(n800), .ZN(n910) );
  XOR2_X1 U888 ( .A(G2067), .B(KEYINPUT37), .Z(n801) );
  XNOR2_X1 U889 ( .A(KEYINPUT89), .B(n801), .ZN(n825) );
  NAND2_X1 U890 ( .A1(n910), .A2(n825), .ZN(n947) );
  XOR2_X1 U891 ( .A(KEYINPUT38), .B(KEYINPUT90), .Z(n803) );
  NAND2_X1 U892 ( .A1(G105), .A2(n898), .ZN(n802) );
  XNOR2_X1 U893 ( .A(n803), .B(n802), .ZN(n807) );
  NAND2_X1 U894 ( .A1(G129), .A2(n893), .ZN(n805) );
  NAND2_X1 U895 ( .A1(G141), .A2(n897), .ZN(n804) );
  NAND2_X1 U896 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n809) );
  NAND2_X1 U898 ( .A1(n894), .A2(G117), .ZN(n808) );
  NAND2_X1 U899 ( .A1(n809), .A2(n808), .ZN(n904) );
  NOR2_X1 U900 ( .A1(G1996), .A2(n904), .ZN(n929) );
  NAND2_X1 U901 ( .A1(G1996), .A2(n904), .ZN(n810) );
  XOR2_X1 U902 ( .A(KEYINPUT91), .B(n810), .Z(n818) );
  NAND2_X1 U903 ( .A1(G119), .A2(n893), .ZN(n812) );
  NAND2_X1 U904 ( .A1(G131), .A2(n897), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n816) );
  NAND2_X1 U906 ( .A1(G107), .A2(n894), .ZN(n814) );
  NAND2_X1 U907 ( .A1(G95), .A2(n898), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n815) );
  OR2_X1 U909 ( .A1(n816), .A2(n815), .ZN(n879) );
  NAND2_X1 U910 ( .A1(G1991), .A2(n879), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n818), .A2(n817), .ZN(n836) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n879), .ZN(n932) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n819) );
  XNOR2_X1 U914 ( .A(KEYINPUT106), .B(n819), .ZN(n820) );
  NOR2_X1 U915 ( .A1(n932), .A2(n820), .ZN(n821) );
  XOR2_X1 U916 ( .A(KEYINPUT107), .B(n821), .Z(n822) );
  NOR2_X1 U917 ( .A1(n836), .A2(n822), .ZN(n823) );
  NOR2_X1 U918 ( .A1(n929), .A2(n823), .ZN(n824) );
  XNOR2_X1 U919 ( .A(n824), .B(KEYINPUT39), .ZN(n827) );
  NOR2_X1 U920 ( .A1(n910), .A2(n825), .ZN(n837) );
  INV_X1 U921 ( .A(n837), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U923 ( .A1(n947), .A2(n828), .ZN(n832) );
  INV_X1 U924 ( .A(n829), .ZN(n830) );
  NOR2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n838) );
  NAND2_X1 U926 ( .A1(n832), .A2(n838), .ZN(n835) );
  INV_X1 U927 ( .A(n835), .ZN(n841) );
  NOR2_X1 U928 ( .A1(n837), .A2(n836), .ZN(n934) );
  XOR2_X1 U929 ( .A(G1986), .B(G290), .Z(n988) );
  NAND2_X1 U930 ( .A1(n934), .A2(n988), .ZN(n839) );
  NAND2_X1 U931 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U932 ( .A(n842), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U933 ( .A1(G2106), .A2(n843), .ZN(G217) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n844) );
  NAND2_X1 U935 ( .A1(G661), .A2(n844), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n845) );
  NAND2_X1 U937 ( .A1(n846), .A2(n845), .ZN(G188) );
  INV_X1 U939 ( .A(G132), .ZN(G219) );
  INV_X1 U940 ( .A(G120), .ZN(G236) );
  INV_X1 U941 ( .A(G108), .ZN(G238) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  INV_X1 U943 ( .A(G82), .ZN(G220) );
  INV_X1 U944 ( .A(G69), .ZN(G235) );
  NOR2_X1 U945 ( .A1(n848), .A2(n847), .ZN(G325) );
  INV_X1 U946 ( .A(G325), .ZN(G261) );
  INV_X1 U947 ( .A(n849), .ZN(G319) );
  XOR2_X1 U948 ( .A(G2474), .B(G1971), .Z(n851) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1981), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U951 ( .A(n852), .B(KEYINPUT112), .Z(n854) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1991), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U954 ( .A(G1976), .B(G1956), .Z(n856) );
  XNOR2_X1 U955 ( .A(G1966), .B(G1961), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U957 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U958 ( .A(KEYINPUT41), .B(KEYINPUT113), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(G229) );
  XOR2_X1 U960 ( .A(G2100), .B(KEYINPUT111), .Z(n862) );
  XNOR2_X1 U961 ( .A(G2678), .B(KEYINPUT43), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U963 ( .A(KEYINPUT42), .B(G2090), .Z(n864) );
  XNOR2_X1 U964 ( .A(G2067), .B(G2072), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U966 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U967 ( .A(KEYINPUT110), .B(G2096), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n868), .B(n867), .ZN(n870) );
  XOR2_X1 U969 ( .A(G2084), .B(G2078), .Z(n869) );
  XNOR2_X1 U970 ( .A(n870), .B(n869), .ZN(G227) );
  NAND2_X1 U971 ( .A1(G112), .A2(n894), .ZN(n871) );
  XNOR2_X1 U972 ( .A(n871), .B(KEYINPUT114), .ZN(n874) );
  NAND2_X1 U973 ( .A1(G124), .A2(n893), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n872), .B(KEYINPUT44), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n878) );
  NAND2_X1 U976 ( .A1(G136), .A2(n897), .ZN(n876) );
  NAND2_X1 U977 ( .A1(G100), .A2(n898), .ZN(n875) );
  NAND2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U979 ( .A1(n878), .A2(n877), .ZN(G162) );
  XNOR2_X1 U980 ( .A(KEYINPUT48), .B(KEYINPUT116), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n879), .B(KEYINPUT46), .ZN(n880) );
  XNOR2_X1 U982 ( .A(n881), .B(n880), .ZN(n890) );
  NAND2_X1 U983 ( .A1(G127), .A2(n893), .ZN(n883) );
  NAND2_X1 U984 ( .A1(G115), .A2(n894), .ZN(n882) );
  NAND2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n884), .B(KEYINPUT47), .ZN(n886) );
  NAND2_X1 U987 ( .A1(G139), .A2(n897), .ZN(n885) );
  NAND2_X1 U988 ( .A1(n886), .A2(n885), .ZN(n889) );
  NAND2_X1 U989 ( .A1(G103), .A2(n898), .ZN(n887) );
  XNOR2_X1 U990 ( .A(KEYINPUT115), .B(n887), .ZN(n888) );
  NOR2_X1 U991 ( .A1(n889), .A2(n888), .ZN(n940) );
  XOR2_X1 U992 ( .A(n890), .B(n940), .Z(n892) );
  XNOR2_X1 U993 ( .A(G160), .B(G164), .ZN(n891) );
  XNOR2_X1 U994 ( .A(n892), .B(n891), .ZN(n907) );
  NAND2_X1 U995 ( .A1(G130), .A2(n893), .ZN(n896) );
  NAND2_X1 U996 ( .A1(G118), .A2(n894), .ZN(n895) );
  NAND2_X1 U997 ( .A1(n896), .A2(n895), .ZN(n903) );
  NAND2_X1 U998 ( .A1(G142), .A2(n897), .ZN(n900) );
  NAND2_X1 U999 ( .A1(G106), .A2(n898), .ZN(n899) );
  NAND2_X1 U1000 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U1001 ( .A(n901), .B(KEYINPUT45), .Z(n902) );
  NOR2_X1 U1002 ( .A1(n903), .A2(n902), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1004 ( .A(n907), .B(n906), .Z(n909) );
  XNOR2_X1 U1005 ( .A(G162), .B(n936), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n912), .ZN(G395) );
  XOR2_X1 U1009 ( .A(KEYINPUT117), .B(G286), .Z(n915) );
  XNOR2_X1 U1010 ( .A(G171), .B(n913), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n915), .B(n914), .ZN(n918) );
  XNOR2_X1 U1012 ( .A(n994), .B(n916), .ZN(n917) );
  XNOR2_X1 U1013 ( .A(n918), .B(n917), .ZN(n919) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n919), .ZN(G397) );
  NOR2_X1 U1015 ( .A1(G229), .A2(G227), .ZN(n921) );
  XNOR2_X1 U1016 ( .A(KEYINPUT49), .B(KEYINPUT118), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(n921), .B(n920), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(G401), .A2(n922), .ZN(n923) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n923), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(KEYINPUT119), .B(n924), .ZN(n926) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(KEYINPUT120), .B(n927), .ZN(G225) );
  XNOR2_X1 U1024 ( .A(KEYINPUT121), .B(G225), .ZN(G308) );
  XOR2_X1 U1025 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1027 ( .A(KEYINPUT51), .B(n930), .Z(n939) );
  XOR2_X1 U1028 ( .A(G160), .B(G2084), .Z(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(n937), .B(KEYINPUT122), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n945) );
  XOR2_X1 U1034 ( .A(G164), .B(G2078), .Z(n942) );
  XNOR2_X1 U1035 ( .A(n954), .B(n940), .ZN(n941) );
  NOR2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1037 ( .A(KEYINPUT50), .B(n943), .Z(n944) );
  NOR2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(n948), .B(KEYINPUT52), .ZN(n949) );
  XNOR2_X1 U1041 ( .A(KEYINPUT123), .B(n949), .ZN(n950) );
  INV_X1 U1042 ( .A(KEYINPUT55), .ZN(n973) );
  NAND2_X1 U1043 ( .A1(n950), .A2(n973), .ZN(n951) );
  NAND2_X1 U1044 ( .A1(n951), .A2(G29), .ZN(n1030) );
  XNOR2_X1 U1045 ( .A(KEYINPUT54), .B(G34), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(n952), .B(KEYINPUT125), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(G2084), .B(n953), .ZN(n971) );
  XNOR2_X1 U1048 ( .A(G2090), .B(G35), .ZN(n969) );
  XNOR2_X1 U1049 ( .A(G33), .B(n954), .ZN(n963) );
  XOR2_X1 U1050 ( .A(G2067), .B(G26), .Z(n957) );
  XNOR2_X1 U1051 ( .A(n955), .B(G32), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n961) );
  XOR2_X1 U1053 ( .A(G1991), .B(G25), .Z(n958) );
  NAND2_X1 U1054 ( .A1(n958), .A2(G28), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(KEYINPUT124), .B(n959), .ZN(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n966) );
  XOR2_X1 U1058 ( .A(G27), .B(n964), .Z(n965) );
  NOR2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(KEYINPUT53), .B(n967), .ZN(n968) );
  NOR2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1063 ( .A(n973), .B(n972), .ZN(n975) );
  INV_X1 U1064 ( .A(G29), .ZN(n974) );
  NAND2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1066 ( .A1(G11), .A2(n976), .ZN(n1028) );
  XNOR2_X1 U1067 ( .A(G16), .B(KEYINPUT56), .ZN(n1000) );
  XOR2_X1 U1068 ( .A(G168), .B(G1966), .Z(n977) );
  NOR2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1070 ( .A(KEYINPUT57), .B(n979), .Z(n998) );
  XOR2_X1 U1071 ( .A(G171), .B(G1961), .Z(n982) );
  XNOR2_X1 U1072 ( .A(n980), .B(G1348), .ZN(n981) );
  NOR2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n993) );
  XNOR2_X1 U1074 ( .A(G299), .B(G1956), .ZN(n985) );
  XNOR2_X1 U1075 ( .A(n983), .B(KEYINPUT126), .ZN(n984) );
  NOR2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n991) );
  XNOR2_X1 U1078 ( .A(G166), .B(G1971), .ZN(n989) );
  NAND2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n996) );
  XNOR2_X1 U1082 ( .A(G1341), .B(n994), .ZN(n995) );
  NOR2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1085 ( .A1(n1000), .A2(n999), .ZN(n1026) );
  INV_X1 U1086 ( .A(G16), .ZN(n1024) );
  XNOR2_X1 U1087 ( .A(G5), .B(n1001), .ZN(n1014) );
  XNOR2_X1 U1088 ( .A(G1348), .B(KEYINPUT59), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(n1002), .B(G4), .ZN(n1006) );
  XNOR2_X1 U1090 ( .A(G1956), .B(G20), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G19), .B(G1341), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XOR2_X1 U1094 ( .A(KEYINPUT127), .B(G1981), .Z(n1007) );
  XNOR2_X1 U1095 ( .A(G6), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1097 ( .A(KEYINPUT60), .B(n1010), .Z(n1012) );
  XNOR2_X1 U1098 ( .A(G1966), .B(G21), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1021) );
  XNOR2_X1 U1101 ( .A(G1971), .B(G22), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(G23), .B(G1976), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XOR2_X1 U1104 ( .A(G1986), .B(G24), .Z(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(KEYINPUT58), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(KEYINPUT61), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1112 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

