//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202));
  INV_X1    g001(.A(G183gat), .ZN(new_n203));
  INV_X1    g002(.A(G190gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT26), .ZN(new_n208));
  NOR2_X1   g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n205), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT27), .B(G183gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT69), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(new_n204), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT28), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT70), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT27), .ZN(new_n219));
  AOI211_X1 g018(.A(KEYINPUT28), .B(G190gat), .C1(new_n219), .C2(KEYINPUT68), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(KEYINPUT68), .B2(new_n213), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n217), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n218), .B1(new_n217), .B2(new_n221), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n212), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n209), .B1(KEYINPUT23), .B2(new_n206), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n225), .B1(KEYINPUT23), .B2(new_n209), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n205), .A2(KEYINPUT66), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n205), .A2(KEYINPUT66), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n233));
  MUX2_X1   g032(.A(G183gat), .B(new_n233), .S(G190gat), .Z(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n230), .A2(new_n231), .ZN(new_n236));
  OAI211_X1 g035(.A(KEYINPUT25), .B(new_n226), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n234), .B1(KEYINPUT24), .B2(new_n205), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n239));
  OR2_X1    g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n239), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n240), .A2(new_n226), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n237), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n224), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G113gat), .B(G120gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n246), .A2(KEYINPUT1), .ZN(new_n247));
  XNOR2_X1  g046(.A(G127gat), .B(G134gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n202), .B1(new_n245), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G227gat), .A2(G233gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n245), .A2(new_n249), .ZN(new_n252));
  INV_X1    g051(.A(new_n249), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n224), .A2(new_n244), .A3(KEYINPUT71), .A4(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n250), .A2(new_n251), .A3(new_n252), .A4(new_n254), .ZN(new_n255));
  OR2_X1    g054(.A1(new_n255), .A2(KEYINPUT34), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(KEYINPUT34), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n250), .A2(new_n252), .A3(new_n254), .ZN(new_n259));
  INV_X1    g058(.A(new_n251), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT33), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G15gat), .B(G43gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(G71gat), .B(G99gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n256), .B(new_n257), .C1(new_n261), .C2(new_n264), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n259), .A2(new_n260), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT32), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G78gat), .B(G106gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT31), .B(G50gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT29), .ZN(new_n275));
  INV_X1    g074(.A(G141gat), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n276), .A2(G148gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT75), .B(G148gat), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n277), .B1(new_n278), .B2(G141gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(G155gat), .B(G162gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT2), .ZN(new_n281));
  NAND2_X1  g080(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n280), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT77), .ZN(new_n285));
  OR3_X1    g084(.A1(new_n279), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n285), .B1(new_n279), .B2(new_n284), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G141gat), .B(G148gat), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(KEYINPUT74), .B(KEYINPUT2), .Z(new_n291));
  AOI21_X1  g090(.A(new_n280), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n275), .B1(new_n294), .B2(KEYINPUT3), .ZN(new_n295));
  XNOR2_X1  g094(.A(G197gat), .B(G204gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT22), .ZN(new_n297));
  INV_X1    g096(.A(G211gat), .ZN(new_n298));
  INV_X1    g097(.A(G218gat), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G211gat), .B(G218gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n295), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n305), .B1(new_n303), .B2(KEYINPUT29), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n294), .A2(new_n306), .ZN(new_n307));
  AND4_X1   g106(.A1(G228gat), .A2(new_n304), .A3(G233gat), .A4(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n303), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(KEYINPUT84), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n302), .A2(new_n296), .A3(new_n300), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT84), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n275), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n305), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(new_n294), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n304), .A2(new_n315), .B1(G228gat), .B2(G233gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n308), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G22gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n274), .B1(new_n319), .B2(KEYINPUT85), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n317), .B(new_n318), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n270), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n266), .A2(new_n323), .A3(new_n267), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n271), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G226gat), .A2(G233gat), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n326), .B1(new_n224), .B2(new_n244), .ZN(new_n327));
  XOR2_X1   g126(.A(new_n327), .B(KEYINPUT73), .Z(new_n328));
  INV_X1    g127(.A(KEYINPUT72), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n245), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n224), .A2(new_n244), .A3(KEYINPUT72), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n326), .B1(new_n332), .B2(KEYINPUT29), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n303), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n332), .A2(G226gat), .A3(G233gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n245), .A2(new_n275), .A3(new_n326), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n303), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G8gat), .B(G36gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(G64gat), .B(G92gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n340), .B(new_n341), .Z(new_n342));
  NAND4_X1  g141(.A1(new_n335), .A2(new_n339), .A3(KEYINPUT30), .A4(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n342), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n309), .B1(new_n328), .B2(new_n333), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n344), .B1(new_n345), .B2(new_n338), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n345), .A2(new_n338), .A3(new_n344), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n348), .A2(KEYINPUT30), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NOR3_X1   g149(.A1(new_n325), .A2(new_n350), .A3(KEYINPUT35), .ZN(new_n351));
  XNOR2_X1  g150(.A(G1gat), .B(G29gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT0), .ZN(new_n353));
  XNOR2_X1  g152(.A(G57gat), .B(G85gat), .ZN(new_n354));
  XOR2_X1   g153(.A(new_n353), .B(new_n354), .Z(new_n355));
  XOR2_X1   g154(.A(new_n355), .B(KEYINPUT86), .Z(new_n356));
  AOI21_X1  g155(.A(new_n253), .B1(new_n294), .B2(KEYINPUT3), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n357), .B1(KEYINPUT3), .B2(new_n294), .ZN(new_n358));
  NAND2_X1  g157(.A1(G225gat), .A2(G233gat), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n359), .B(KEYINPUT78), .Z(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT79), .B1(new_n294), .B2(new_n249), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n288), .A2(new_n364), .A3(new_n253), .A4(new_n293), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT4), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT80), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n294), .A2(new_n249), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT4), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n371), .B1(new_n366), .B2(new_n367), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n362), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  OR2_X1    g172(.A1(new_n373), .A2(KEYINPUT81), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(KEYINPUT81), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n294), .A2(new_n249), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n363), .A2(new_n365), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n360), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT5), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n374), .A2(new_n375), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n363), .A2(new_n365), .ZN(new_n383));
  OR3_X1    g182(.A1(new_n383), .A2(KEYINPUT83), .A3(new_n370), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n370), .ZN(new_n385));
  OAI211_X1 g184(.A(KEYINPUT83), .B(new_n385), .C1(new_n383), .C2(new_n370), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  OR3_X1    g186(.A1(new_n387), .A2(KEYINPUT5), .A3(new_n362), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n382), .A2(KEYINPUT89), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT89), .B1(new_n382), .B2(new_n388), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n356), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n382), .A2(new_n355), .A3(new_n388), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT6), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n355), .B1(new_n382), .B2(new_n388), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT6), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n351), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n350), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n398), .B1(new_n394), .B2(new_n397), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n324), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n323), .B1(new_n266), .B2(new_n267), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n406), .A2(KEYINPUT90), .A3(new_n322), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT90), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n325), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n403), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT35), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n400), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT36), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(new_n404), .B2(new_n405), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n271), .A2(KEYINPUT36), .A3(new_n324), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n345), .A2(new_n338), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT37), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n342), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n420), .B1(new_n419), .B2(new_n418), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT38), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n336), .A2(new_n337), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n419), .B1(new_n423), .B2(new_n303), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n334), .A2(new_n309), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT38), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n348), .B1(new_n420), .B2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n396), .A2(new_n398), .A3(new_n422), .A4(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n322), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT88), .ZN(new_n430));
  INV_X1    g229(.A(new_n356), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n384), .A2(new_n358), .A3(new_n386), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n360), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n431), .B1(new_n433), .B2(KEYINPUT39), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n363), .A2(new_n361), .A3(new_n365), .A4(new_n376), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n435), .A2(KEYINPUT87), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT39), .B1(new_n435), .B2(KEYINPUT87), .ZN(new_n437));
  AOI211_X1 g236(.A(new_n436), .B(new_n437), .C1(new_n432), .C2(new_n360), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n430), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT40), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n430), .B(KEYINPUT40), .C1(new_n434), .C2(new_n438), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n347), .A2(new_n349), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n429), .B1(new_n443), .B2(new_n391), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n417), .B1(new_n428), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n403), .A2(new_n429), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n412), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G134gat), .B(G162gat), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT15), .ZN(new_n453));
  XOR2_X1   g252(.A(G43gat), .B(G50gat), .Z(new_n454));
  NOR2_X1   g253(.A1(G29gat), .A2(G36gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT14), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT14), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n457), .B1(G29gat), .B2(G36gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n459), .A2(KEYINPUT91), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT92), .B(G29gat), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n459), .A2(KEYINPUT91), .B1(G36gat), .B2(new_n461), .ZN(new_n462));
  AOI211_X1 g261(.A(new_n453), .B(new_n454), .C1(new_n460), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n454), .A2(new_n453), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n461), .A2(G36gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n454), .A2(new_n453), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n466), .A2(new_n467), .A3(new_n459), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  OR2_X1    g268(.A1(new_n469), .A2(KEYINPUT17), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(KEYINPUT17), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT99), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n472), .A2(G85gat), .A3(G92gat), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT100), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n474), .A2(KEYINPUT7), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT7), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n476), .A2(KEYINPUT100), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n473), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G85gat), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n479), .A2(KEYINPUT99), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n476), .A2(KEYINPUT100), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n474), .A2(KEYINPUT7), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n480), .A2(new_n481), .A3(new_n482), .A4(G92gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  AND2_X1   g283(.A1(G99gat), .A2(G106gat), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT8), .ZN(new_n486));
  OAI22_X1  g285(.A1(new_n485), .A2(new_n486), .B1(G85gat), .B2(G92gat), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  OR2_X1    g288(.A1(G99gat), .A2(G106gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(KEYINPUT101), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT101), .ZN(new_n493));
  NOR2_X1   g292(.A1(G99gat), .A2(G106gat), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n493), .B1(new_n485), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n489), .A2(new_n497), .ZN(new_n498));
  AND4_X1   g297(.A1(KEYINPUT102), .A2(new_n484), .A3(new_n496), .A4(new_n488), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n487), .B1(new_n478), .B2(new_n483), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT102), .B1(new_n500), .B2(new_n496), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n498), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n470), .A2(new_n471), .A3(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G190gat), .B(G218gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(KEYINPUT103), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  AND3_X1   g305(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n507));
  INV_X1    g306(.A(new_n469), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n484), .A2(new_n496), .A3(new_n488), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT102), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n500), .A2(KEYINPUT102), .A3(new_n496), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n511), .A2(new_n512), .B1(new_n497), .B2(new_n489), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n507), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n503), .A2(new_n506), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n506), .B1(new_n503), .B2(new_n514), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n452), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n517), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n519), .A2(new_n451), .A3(new_n515), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT93), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT16), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n525), .B1(new_n526), .B2(G1gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n523), .B(KEYINPUT93), .ZN(new_n528));
  INV_X1    g327(.A(G1gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G8gat), .ZN(new_n532));
  INV_X1    g331(.A(G8gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n527), .A2(new_n533), .A3(new_n530), .ZN(new_n534));
  AND2_X1   g333(.A1(G71gat), .A2(G78gat), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n535), .A2(KEYINPUT96), .ZN(new_n536));
  NOR2_X1   g335(.A1(G71gat), .A2(G78gat), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT96), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n535), .A2(KEYINPUT9), .ZN(new_n539));
  XNOR2_X1  g338(.A(G57gat), .B(G64gat), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n536), .B(new_n538), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G57gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(G64gat), .ZN(new_n543));
  INV_X1    g342(.A(G64gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(G57gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT9), .ZN(new_n546));
  NAND2_X1  g345(.A1(G71gat), .A2(G78gat), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n543), .A2(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n537), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT97), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(new_n550), .A3(new_n547), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT97), .B1(new_n535), .B2(new_n537), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n548), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n541), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT21), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n532), .A2(new_n534), .A3(new_n556), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n557), .A2(KEYINPUT98), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(KEYINPUT98), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n561));
  INV_X1    g360(.A(G155gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n563), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n558), .A2(new_n559), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT21), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n554), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G127gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(G183gat), .B(G211gat), .Z(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n571), .B(G127gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n574), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n567), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n564), .A2(new_n575), .A3(new_n578), .A4(new_n566), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR3_X1   g381(.A1(new_n522), .A2(new_n582), .A3(KEYINPUT104), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n511), .A2(new_n512), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT105), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n484), .A2(new_n488), .B1(new_n496), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n492), .A2(new_n495), .A3(KEYINPUT105), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n554), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n502), .A2(new_n554), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G230gat), .A2(G233gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G120gat), .B(G148gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(G176gat), .B(G204gat), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n592), .B(new_n593), .Z(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n496), .A2(new_n585), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n489), .A2(new_n587), .A3(new_n597), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n555), .B(new_n598), .C1(new_n499), .C2(new_n501), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT10), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n599), .B(new_n600), .C1(new_n513), .C2(new_n555), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT106), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n502), .A2(new_n554), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT106), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n603), .A2(new_n604), .A3(new_n600), .A4(new_n599), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n554), .A2(new_n600), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n513), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT107), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n513), .A2(KEYINPUT107), .A3(new_n606), .ZN(new_n610));
  AOI22_X1  g409(.A1(new_n602), .A2(new_n605), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT108), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n590), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n602), .A2(new_n605), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n609), .A2(new_n610), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n614), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n596), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT109), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT109), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n619), .B(new_n596), .C1(new_n613), .C2(new_n616), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n594), .B(KEYINPUT110), .Z(new_n622));
  INV_X1    g421(.A(new_n590), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n611), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n622), .B1(new_n624), .B2(new_n591), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT104), .ZN(new_n627));
  INV_X1    g426(.A(new_n582), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n627), .B1(new_n628), .B2(new_n521), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n532), .A2(new_n534), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT94), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT94), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n532), .A2(new_n632), .A3(new_n534), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n631), .A2(new_n470), .A3(new_n471), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G229gat), .A2(G233gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n630), .A2(new_n508), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT18), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT95), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n469), .A2(new_n532), .A3(new_n534), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n636), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n635), .B(KEYINPUT13), .Z(new_n643));
  NAND3_X1  g442(.A1(new_n630), .A2(new_n508), .A3(KEYINPUT95), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n634), .A2(KEYINPUT18), .A3(new_n635), .A4(new_n636), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n639), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G113gat), .B(G141gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G197gat), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT11), .B(G169gat), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(KEYINPUT12), .Z(new_n652));
  NAND2_X1  g451(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n652), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n639), .A2(new_n654), .A3(new_n645), .A4(new_n646), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NOR4_X1   g456(.A1(new_n583), .A2(new_n626), .A3(new_n629), .A4(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n448), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n659), .A2(new_n402), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(new_n529), .ZN(G1324gat));
  AND2_X1   g460(.A1(new_n448), .A2(new_n658), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n350), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT42), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n526), .A2(new_n533), .ZN(new_n665));
  NOR2_X1   g464(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OR3_X1    g466(.A1(new_n663), .A2(new_n664), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n664), .B1(new_n663), .B2(new_n667), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n663), .A2(G8gat), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(G1325gat));
  AOI21_X1  g470(.A(G15gat), .B1(new_n662), .B2(new_n406), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n417), .A2(G15gat), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n673), .B(KEYINPUT111), .Z(new_n674));
  AOI21_X1  g473(.A(new_n672), .B1(new_n662), .B2(new_n674), .ZN(G1326gat));
  INV_X1    g474(.A(KEYINPUT112), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n676), .B1(new_n662), .B2(new_n429), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n659), .A2(KEYINPUT112), .A3(new_n322), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  AOI21_X1  g480(.A(new_n521), .B1(new_n412), .B2(new_n447), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n626), .A2(new_n657), .A3(new_n628), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n684), .A2(new_n402), .A3(new_n461), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n685), .A2(KEYINPUT45), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n402), .A2(new_n349), .A3(new_n347), .ZN(new_n687));
  INV_X1    g486(.A(new_n409), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n325), .A2(new_n408), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT35), .ZN(new_n691));
  AOI22_X1  g490(.A1(new_n691), .A2(new_n400), .B1(new_n445), .B2(new_n446), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT44), .B1(new_n692), .B2(new_n521), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT113), .B1(new_n687), .B2(new_n322), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n428), .A2(new_n444), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT113), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n403), .A2(new_n696), .A3(new_n429), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n694), .A2(new_n695), .A3(new_n416), .A4(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n412), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT114), .B(KEYINPUT44), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(new_n522), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n693), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n402), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(new_n703), .A3(new_n683), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n461), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n685), .A2(KEYINPUT45), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n686), .A2(new_n705), .A3(new_n706), .ZN(G1328gat));
  NOR3_X1   g506(.A1(new_n684), .A2(G36gat), .A3(new_n401), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT46), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n702), .A2(new_n350), .A3(new_n683), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(G36gat), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(G1329gat));
  NAND4_X1  g511(.A1(new_n702), .A2(G43gat), .A3(new_n417), .A4(new_n683), .ZN(new_n713));
  INV_X1    g512(.A(G43gat), .ZN(new_n714));
  INV_X1    g513(.A(new_n406), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n684), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT47), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT47), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n713), .A2(new_n719), .A3(new_n716), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(G1330gat));
  NAND4_X1  g520(.A1(new_n702), .A2(G50gat), .A3(new_n429), .A4(new_n683), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT115), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n723), .A2(KEYINPUT48), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n682), .A2(new_n429), .A3(new_n683), .ZN(new_n725));
  INV_X1    g524(.A(G50gat), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n725), .A2(new_n726), .B1(new_n723), .B2(KEYINPUT48), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n722), .A2(new_n724), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n724), .B1(new_n722), .B2(new_n727), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(G1331gat));
  INV_X1    g529(.A(new_n626), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(new_n656), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n629), .A2(new_n583), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n699), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n402), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(new_n542), .ZN(G1332gat));
  NOR2_X1   g536(.A1(new_n735), .A2(new_n401), .ZN(new_n738));
  NOR2_X1   g537(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n739));
  AND2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n738), .B2(new_n739), .ZN(G1333gat));
  OAI21_X1  g541(.A(G71gat), .B1(new_n735), .B2(new_n416), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n715), .A2(G71gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n735), .B2(new_n744), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g545(.A1(new_n735), .A2(new_n322), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n582), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n702), .A2(new_n703), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT116), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n749), .B1(new_n693), .B2(new_n701), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT116), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n753), .A2(new_n754), .A3(new_n703), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n752), .A2(G85gat), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n521), .B1(new_n698), .B2(new_n412), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n656), .A2(new_n628), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT51), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n757), .A2(KEYINPUT51), .A3(new_n758), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n762), .A2(new_n479), .A3(new_n703), .A4(new_n626), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n756), .A2(new_n763), .ZN(G1336gat));
  INV_X1    g563(.A(G92gat), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(new_n753), .B2(new_n350), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n401), .A2(G92gat), .A3(new_n731), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n768), .B1(new_n760), .B2(new_n761), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT52), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n682), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n700), .ZN(new_n773));
  AOI211_X1 g572(.A(new_n521), .B(new_n773), .C1(new_n698), .C2(new_n412), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n350), .B(new_n750), .C1(new_n772), .C2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G92gat), .ZN(new_n776));
  INV_X1    g575(.A(new_n761), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n767), .B1(new_n777), .B2(new_n759), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n770), .A2(new_n780), .ZN(G1337gat));
  NAND2_X1  g580(.A1(new_n753), .A2(new_n417), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G99gat), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n715), .A2(G99gat), .A3(new_n731), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n762), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1338gat));
  INV_X1    g585(.A(G106gat), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n787), .B1(new_n753), .B2(new_n429), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n322), .A2(new_n731), .A3(G106gat), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT117), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n791), .B1(new_n760), .B2(new_n761), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT53), .B1(new_n788), .B2(new_n792), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n429), .B(new_n750), .C1(new_n772), .C2(new_n774), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G106gat), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n790), .B1(new_n777), .B2(new_n759), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n793), .A2(new_n798), .ZN(G1339gat));
  NOR2_X1   g598(.A1(new_n657), .A2(G113gat), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n733), .A2(new_n731), .A3(new_n657), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n801), .B(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT120), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n805), .B1(new_n611), .B2(new_n623), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n613), .B2(new_n616), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n594), .B1(new_n624), .B2(new_n805), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n804), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AOI211_X1 g610(.A(KEYINPUT120), .B(KEYINPUT55), .C1(new_n807), .C2(new_n808), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n635), .B1(new_n634), .B2(new_n636), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n643), .B1(new_n642), .B2(new_n644), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n651), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n655), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n813), .A2(new_n522), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n807), .A2(KEYINPUT55), .A3(new_n808), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n820), .A2(KEYINPUT119), .B1(new_n618), .B2(new_n620), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n807), .A2(new_n808), .A3(new_n822), .A4(KEYINPUT55), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT121), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n813), .A2(new_n656), .A3(new_n823), .A4(new_n821), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n626), .A2(new_n818), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n809), .A2(new_n810), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT120), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n809), .A2(new_n804), .A3(new_n810), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n820), .A2(KEYINPUT119), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n835), .A2(new_n621), .A3(new_n656), .A4(new_n823), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n827), .B(new_n829), .C1(new_n834), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n521), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n826), .B1(new_n830), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n803), .B1(new_n839), .B2(new_n582), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n402), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n841), .B(new_n401), .C1(new_n688), .C2(new_n689), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n842), .A2(KEYINPUT122), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(KEYINPUT122), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n800), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n840), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n402), .A2(new_n350), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n846), .A2(new_n322), .A3(new_n406), .A4(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(G113gat), .B1(new_n848), .B2(new_n657), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n845), .A2(new_n849), .ZN(G1340gat));
  NOR2_X1   g649(.A1(new_n731), .A2(G120gat), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n851), .B1(new_n843), .B2(new_n844), .ZN(new_n852));
  OAI21_X1  g651(.A(G120gat), .B1(new_n848), .B2(new_n731), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(G1341gat));
  OAI21_X1  g653(.A(G127gat), .B1(new_n848), .B2(new_n582), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n628), .A2(new_n572), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n842), .B2(new_n856), .ZN(G1342gat));
  OR2_X1    g656(.A1(new_n521), .A2(G134gat), .ZN(new_n858));
  OR3_X1    g657(.A1(new_n842), .A2(KEYINPUT56), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(G134gat), .B1(new_n848), .B2(new_n521), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT56), .B1(new_n842), .B2(new_n858), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(G1343gat));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  INV_X1    g662(.A(new_n803), .ZN(new_n864));
  INV_X1    g663(.A(new_n605), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n604), .B1(new_n589), .B2(new_n600), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n615), .B(new_n623), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT54), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n615), .B1(new_n865), .B2(new_n866), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n623), .B1(new_n869), .B2(KEYINPUT108), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n611), .A2(new_n612), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n590), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n595), .B1(new_n873), .B2(KEYINPUT54), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT123), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n807), .A2(new_n876), .A3(new_n808), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n810), .A3(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n875), .A2(KEYINPUT124), .A3(new_n810), .A4(new_n877), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n829), .B1(new_n882), .B2(new_n836), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n522), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI211_X1 g684(.A(KEYINPUT125), .B(new_n829), .C1(new_n882), .C2(new_n836), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n825), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n864), .B1(new_n887), .B2(new_n628), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n863), .B1(new_n888), .B2(new_n429), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n840), .A2(KEYINPUT57), .A3(new_n322), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n847), .A2(new_n416), .ZN(new_n891));
  NOR4_X1   g690(.A1(new_n889), .A2(new_n657), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT126), .B1(new_n892), .B2(new_n276), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n841), .A2(new_n401), .A3(new_n429), .A4(new_n416), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n276), .A3(new_n656), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n896), .B1(new_n892), .B2(new_n276), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n893), .A2(new_n897), .A3(KEYINPUT58), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT58), .ZN(new_n899));
  OAI221_X1 g698(.A(new_n896), .B1(KEYINPUT126), .B2(new_n899), .C1(new_n892), .C2(new_n276), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(G1344gat));
  NAND3_X1  g700(.A1(new_n895), .A2(new_n278), .A3(new_n626), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n903));
  AOI211_X1 g702(.A(KEYINPUT59), .B(new_n278), .C1(new_n903), .C2(new_n626), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n846), .A2(new_n429), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n801), .B1(new_n887), .B2(new_n628), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n322), .A2(KEYINPUT57), .ZN(new_n908));
  AOI22_X1  g707(.A1(new_n906), .A2(KEYINPUT57), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n909), .A2(new_n416), .A3(new_n626), .A4(new_n847), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n905), .B1(new_n910), .B2(G148gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n902), .B1(new_n904), .B2(new_n911), .ZN(G1345gat));
  NAND3_X1  g711(.A1(new_n895), .A2(new_n562), .A3(new_n628), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n903), .A2(new_n628), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n562), .ZN(G1346gat));
  NOR2_X1   g714(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n283), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n895), .A2(new_n522), .A3(new_n917), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n903), .A2(new_n522), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n917), .ZN(G1347gat));
  NOR2_X1   g719(.A1(new_n840), .A2(new_n703), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n401), .B1(new_n407), .B2(new_n409), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n923), .A2(G169gat), .A3(new_n657), .ZN(new_n924));
  XOR2_X1   g723(.A(new_n924), .B(KEYINPUT127), .Z(new_n925));
  NAND2_X1  g724(.A1(new_n402), .A2(new_n350), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n926), .A2(new_n715), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n846), .A2(new_n322), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G169gat), .B1(new_n928), .B2(new_n657), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n925), .A2(new_n929), .ZN(G1348gat));
  INV_X1    g729(.A(G176gat), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n928), .A2(new_n931), .A3(new_n731), .ZN(new_n932));
  INV_X1    g731(.A(new_n923), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(new_n626), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n932), .B1(new_n934), .B2(new_n931), .ZN(G1349gat));
  OAI21_X1  g734(.A(G183gat), .B1(new_n928), .B2(new_n582), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n628), .A2(new_n215), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n923), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g738(.A1(new_n933), .A2(new_n204), .A3(new_n522), .ZN(new_n940));
  OAI21_X1  g739(.A(G190gat), .B1(new_n928), .B2(new_n521), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n941), .A2(KEYINPUT61), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n941), .A2(KEYINPUT61), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(G1351gat));
  NOR3_X1   g744(.A1(new_n417), .A2(new_n401), .A3(new_n322), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n921), .A2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(G197gat), .B1(new_n948), .B2(new_n656), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n417), .A2(new_n926), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n909), .A2(new_n950), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n656), .A2(G197gat), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(G1352gat));
  NAND3_X1  g752(.A1(new_n909), .A2(new_n626), .A3(new_n950), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(G204gat), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n731), .A2(G204gat), .ZN(new_n956));
  OAI21_X1  g755(.A(KEYINPUT62), .B1(new_n947), .B2(new_n956), .ZN(new_n957));
  OR3_X1    g756(.A1(new_n947), .A2(KEYINPUT62), .A3(new_n956), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n955), .A2(new_n957), .A3(new_n958), .ZN(G1353gat));
  NAND3_X1  g758(.A1(new_n948), .A2(new_n298), .A3(new_n628), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n909), .A2(new_n628), .A3(new_n950), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n961), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT63), .B1(new_n961), .B2(G211gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(G1354gat));
  NAND3_X1  g763(.A1(new_n948), .A2(new_n299), .A3(new_n522), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n951), .A2(new_n522), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n965), .B1(new_n966), .B2(new_n299), .ZN(G1355gat));
endmodule


