//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966;
  INV_X1    g000(.A(KEYINPUT14), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT91), .ZN(new_n208));
  XOR2_X1   g007(.A(G43gat), .B(G50gat), .Z(new_n209));
  INV_X1    g008(.A(KEYINPUT15), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n210), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n208), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n203), .A2(new_n204), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT90), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n206), .B1(new_n205), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n218), .B1(new_n217), .B2(new_n205), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n211), .B1(new_n219), .B2(new_n215), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G15gat), .B(G22gat), .ZN(new_n222));
  INV_X1    g021(.A(G1gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(KEYINPUT16), .A3(new_n223), .ZN(new_n224));
  OAI221_X1 g023(.A(new_n224), .B1(KEYINPUT92), .B2(G8gat), .C1(new_n223), .C2(new_n222), .ZN(new_n225));
  NAND2_X1  g024(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n226));
  XOR2_X1   g025(.A(new_n225), .B(new_n226), .Z(new_n227));
  NOR2_X1   g026(.A1(new_n221), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT17), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n216), .A2(new_n230), .A3(new_n220), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n230), .B1(new_n216), .B2(new_n220), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n227), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n229), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT18), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n216), .A2(new_n220), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT17), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n231), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n228), .B1(new_n241), .B2(new_n227), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(KEYINPUT18), .A3(new_n235), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n221), .B(new_n227), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n235), .B(KEYINPUT13), .Z(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n238), .A2(new_n243), .A3(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(G169gat), .B(G197gat), .Z(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G113gat), .B(G141gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(new_n252), .B(KEYINPUT12), .Z(new_n253));
  NAND2_X1  g052(.A1(new_n247), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n253), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n238), .A2(new_n243), .A3(new_n255), .A4(new_n246), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n254), .A2(KEYINPUT93), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT93), .B1(new_n254), .B2(new_n256), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G228gat), .A2(G233gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT29), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT80), .B(G141gat), .ZN(new_n263));
  INV_X1    g062(.A(G148gat), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT81), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(G141gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT81), .ZN(new_n267));
  INV_X1    g066(.A(G141gat), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n268), .A2(KEYINPUT80), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(KEYINPUT80), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n267), .B(G148gat), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n265), .A2(new_n266), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G155gat), .ZN(new_n273));
  INV_X1    g072(.A(G162gat), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT2), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G155gat), .B(G162gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n272), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT79), .B(KEYINPUT2), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n268), .A2(G148gat), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n278), .B1(new_n266), .B2(new_n279), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n280), .A2(new_n276), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n262), .B1(new_n282), .B2(KEYINPUT3), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n283), .A2(KEYINPUT85), .ZN(new_n284));
  XNOR2_X1  g083(.A(G197gat), .B(G204gat), .ZN(new_n285));
  INV_X1    g084(.A(G211gat), .ZN(new_n286));
  INV_X1    g085(.A(G218gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n285), .B1(KEYINPUT22), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G211gat), .B(G218gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n283), .A2(KEYINPUT85), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n284), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n291), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT3), .B1(new_n294), .B2(new_n262), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT82), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n277), .A2(KEYINPUT82), .A3(new_n281), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n296), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n261), .B1(new_n293), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G22gat), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n283), .A2(new_n291), .B1(G228gat), .B2(G233gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n296), .A2(new_n282), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n302), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n306), .ZN(new_n308));
  OAI21_X1  g107(.A(G22gat), .B1(new_n301), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G78gat), .B(G106gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(KEYINPUT84), .ZN(new_n311));
  XOR2_X1   g110(.A(KEYINPUT31), .B(G50gat), .Z(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n307), .A2(new_n309), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n313), .B1(new_n307), .B2(new_n309), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G1gat), .B(G29gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(G85gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT0), .B(G57gat), .ZN(new_n320));
  XOR2_X1   g119(.A(new_n319), .B(new_n320), .Z(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n298), .A2(KEYINPUT3), .A3(new_n299), .ZN(new_n323));
  INV_X1    g122(.A(G120gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G113gat), .ZN(new_n325));
  INV_X1    g124(.A(G113gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G120gat), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT1), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G127gat), .B(G134gat), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT69), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AND2_X1   g129(.A1(G127gat), .A2(G134gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(G127gat), .A2(G134gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT69), .ZN(new_n334));
  XNOR2_X1  g133(.A(G113gat), .B(G120gat), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n333), .B(new_n334), .C1(new_n335), .C2(KEYINPUT1), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n333), .A2(KEYINPUT1), .ZN(new_n337));
  OR3_X1    g136(.A1(new_n326), .A2(KEYINPUT70), .A3(G120gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n325), .A2(KEYINPUT70), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n339), .A3(new_n327), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n330), .A2(new_n336), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n282), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n323), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n277), .A2(new_n281), .A3(new_n341), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT83), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT83), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n277), .A2(new_n341), .A3(new_n350), .A4(new_n281), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n347), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n349), .A2(new_n347), .A3(new_n351), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n346), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT86), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT86), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n354), .A2(new_n359), .A3(new_n356), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT39), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n322), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n298), .A2(new_n342), .A3(new_n299), .ZN(new_n364));
  INV_X1    g163(.A(new_n348), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n365), .A2(new_n356), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n362), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT87), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n358), .A2(new_n360), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT40), .B1(new_n363), .B2(new_n370), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n354), .A2(new_n359), .A3(new_n356), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n359), .B1(new_n354), .B2(new_n356), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n362), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n374), .A2(new_n370), .A3(KEYINPUT40), .A4(new_n321), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n364), .A2(new_n348), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n366), .A2(new_n347), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n348), .A2(new_n347), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n346), .A2(new_n378), .ZN(new_n379));
  OAI221_X1 g178(.A(KEYINPUT5), .B1(new_n376), .B2(new_n355), .C1(new_n377), .C2(new_n379), .ZN(new_n380));
  OR3_X1    g179(.A1(new_n354), .A2(KEYINPUT5), .A3(new_n356), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n322), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n375), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n371), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT27), .ZN(new_n386));
  INV_X1    g185(.A(G183gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n389));
  AOI21_X1  g188(.A(G190gat), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g189(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n391));
  NOR2_X1   g190(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT67), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n390), .A2(KEYINPUT28), .ZN(new_n395));
  INV_X1    g194(.A(G190gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n389), .ZN(new_n397));
  NOR2_X1   g196(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT67), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n394), .A2(new_n395), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT68), .ZN(new_n404));
  NAND2_X1  g203(.A1(G169gat), .A2(G176gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(G169gat), .ZN(new_n407));
  INV_X1    g206(.A(G176gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n406), .B1(KEYINPUT26), .B2(new_n409), .ZN(new_n410));
  OR2_X1    g209(.A1(new_n409), .A2(KEYINPUT26), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n410), .A2(new_n411), .B1(G183gat), .B2(G190gat), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT68), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n394), .A2(new_n402), .A3(new_n413), .A4(new_n395), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n404), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n407), .A2(new_n408), .A3(KEYINPUT23), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT23), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n417), .B1(G169gat), .B2(G176gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n418), .A3(new_n405), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n387), .B2(new_n396), .ZN(new_n421));
  NAND3_X1  g220(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n422));
  AOI211_X1 g221(.A(KEYINPUT25), .B(new_n419), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n420), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(KEYINPUT64), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n387), .A2(new_n396), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT64), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n427), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n424), .A2(new_n425), .A3(new_n426), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT65), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT65), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n421), .A2(new_n431), .A3(new_n425), .A4(new_n428), .ZN(new_n432));
  INV_X1    g231(.A(new_n419), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n423), .B1(KEYINPUT25), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n415), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(G226gat), .ZN(new_n437));
  INV_X1    g236(.A(G233gat), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n436), .A2(new_n262), .ZN(new_n442));
  INV_X1    g241(.A(new_n439), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(KEYINPUT74), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT74), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT29), .B1(new_n415), .B2(new_n435), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n445), .B1(new_n446), .B2(new_n439), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n441), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT75), .B1(new_n448), .B2(new_n294), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT74), .B1(new_n442), .B2(new_n443), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n446), .A2(new_n445), .A3(new_n439), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n440), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT75), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(new_n453), .A3(new_n291), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n294), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n449), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G64gat), .B(G92gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(new_n204), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT76), .B(G8gat), .ZN(new_n460));
  XOR2_X1   g259(.A(new_n459), .B(new_n460), .Z(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n449), .A2(new_n454), .A3(new_n456), .A4(new_n461), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT30), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XOR2_X1   g265(.A(KEYINPUT77), .B(KEYINPUT30), .Z(new_n467));
  AND3_X1   g266(.A1(new_n464), .A2(KEYINPUT78), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT78), .B1(new_n464), .B2(new_n467), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n463), .B(new_n466), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n385), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT37), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n449), .A2(new_n454), .A3(new_n472), .A4(new_n456), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n455), .A2(new_n291), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n474), .B(KEYINPUT37), .C1(new_n291), .C2(new_n448), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n473), .A2(new_n462), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT38), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n457), .A2(KEYINPUT37), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n462), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT88), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n477), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n473), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n461), .B1(new_n457), .B2(KEYINPUT37), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n483), .B1(new_n484), .B2(KEYINPUT88), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n478), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n380), .A2(new_n381), .A3(new_n321), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT6), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n383), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n382), .A2(KEYINPUT6), .A3(new_n322), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n490), .A3(new_n464), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n317), .B(new_n471), .C1(new_n486), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n436), .A2(new_n342), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n415), .A2(new_n435), .A3(new_n341), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(G227gat), .A2(G233gat), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT32), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT33), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(G15gat), .B(G43gat), .Z(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(KEYINPUT71), .ZN(new_n503));
  XOR2_X1   g302(.A(G71gat), .B(G99gat), .Z(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n499), .A2(new_n501), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n505), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n498), .B(KEYINPUT32), .C1(new_n500), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT34), .B1(new_n497), .B2(KEYINPUT72), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n511), .B1(new_n495), .B2(new_n497), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT73), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n493), .A2(new_n496), .A3(new_n494), .A4(new_n510), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n509), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n515), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n513), .B1(new_n512), .B2(new_n514), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n508), .B(new_n506), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT36), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n516), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n520), .B1(new_n516), .B2(new_n519), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n489), .A2(new_n490), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n316), .B1(new_n526), .B2(new_n470), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n492), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n516), .A2(new_n519), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n316), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n464), .A2(new_n465), .ZN(new_n531));
  INV_X1    g330(.A(new_n469), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n464), .A2(KEYINPUT78), .A3(new_n467), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n530), .A2(new_n534), .A3(new_n525), .A4(new_n463), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT35), .ZN(new_n536));
  INV_X1    g335(.A(new_n470), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT35), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n537), .A2(new_n538), .A3(new_n525), .A4(new_n530), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n260), .B1(new_n528), .B2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT21), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT94), .ZN(new_n546));
  XOR2_X1   g345(.A(G57gat), .B(G64gat), .Z(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(G71gat), .B(G78gat), .Z(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G64gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(G57gat), .ZN(new_n552));
  XOR2_X1   g351(.A(KEYINPUT95), .B(G57gat), .Z(new_n553));
  OAI21_X1  g352(.A(new_n552), .B1(new_n553), .B2(new_n551), .ZN(new_n554));
  INV_X1    g353(.A(new_n549), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(new_n555), .A3(new_n546), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n227), .B1(new_n544), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(new_n387), .ZN(new_n559));
  INV_X1    g358(.A(new_n557), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n559), .B1(KEYINPUT21), .B2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n558), .B(G183gat), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n562), .A2(new_n544), .A3(new_n557), .ZN(new_n563));
  AND4_X1   g362(.A1(G231gat), .A2(new_n561), .A3(new_n563), .A4(G233gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(G127gat), .B(G155gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(G211gat), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n561), .A2(new_n563), .B1(G231gat), .B2(G233gat), .ZN(new_n567));
  NOR3_X1   g366(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n566), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n561), .A2(new_n563), .ZN(new_n570));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n561), .A2(new_n563), .A3(G231gat), .A4(G233gat), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n569), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n543), .B1(new_n568), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n566), .B1(new_n564), .B2(new_n567), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n572), .A2(new_n569), .A3(new_n573), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(new_n542), .A3(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT98), .ZN(new_n580));
  NAND2_X1  g379(.A1(G85gat), .A2(G92gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT7), .ZN(new_n582));
  INV_X1    g381(.A(G99gat), .ZN(new_n583));
  INV_X1    g382(.A(G106gat), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT8), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n582), .B(new_n585), .C1(G85gat), .C2(G92gat), .ZN(new_n586));
  XOR2_X1   g385(.A(G99gat), .B(G106gat), .Z(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n586), .A2(new_n587), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n241), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n591), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n239), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n597), .B(KEYINPUT96), .Z(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n580), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n601), .A2(KEYINPUT98), .A3(new_n598), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n596), .A2(new_n599), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n600), .A2(new_n602), .A3(KEYINPUT97), .ZN(new_n605));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606));
  AOI21_X1  g405(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n606), .B(new_n607), .Z(new_n608));
  AND3_X1   g407(.A1(new_n604), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n604), .B1(new_n605), .B2(new_n608), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT103), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT10), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n586), .A2(new_n587), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT99), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n588), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT100), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n590), .A2(KEYINPUT99), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n616), .A2(new_n617), .A3(new_n560), .A4(new_n618), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n616), .A2(new_n560), .A3(new_n618), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT100), .B1(new_n591), .B2(new_n557), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n613), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n593), .A2(KEYINPUT10), .A3(new_n560), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT101), .ZN(new_n625));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT101), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n622), .A2(new_n627), .A3(new_n623), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G120gat), .B(G148gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(G176gat), .B(G204gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n620), .A2(new_n621), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n634), .B1(new_n617), .B2(new_n620), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n629), .B(new_n633), .C1(new_n626), .C2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n626), .B(KEYINPUT102), .Z(new_n637));
  AND2_X1   g436(.A1(new_n624), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n635), .A2(new_n626), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n632), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n579), .A2(new_n611), .A3(new_n612), .A4(new_n642), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n600), .A2(new_n602), .ZN(new_n644));
  INV_X1    g443(.A(new_n608), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n644), .B(new_n603), .C1(KEYINPUT97), .C2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n604), .A2(new_n605), .A3(new_n608), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n575), .A2(new_n646), .A3(new_n647), .A4(new_n578), .ZN(new_n648));
  OAI21_X1  g447(.A(KEYINPUT103), .B1(new_n648), .B2(new_n641), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n643), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n541), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n651), .A2(new_n525), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(new_n223), .ZN(G1324gat));
  INV_X1    g452(.A(new_n651), .ZN(new_n654));
  NAND2_X1  g453(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n655));
  OR2_X1    g454(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n654), .A2(new_n470), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT42), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(G8gat), .B1(new_n651), .B2(new_n537), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(G1325gat));
  INV_X1    g461(.A(new_n523), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n663), .A2(KEYINPUT105), .A3(new_n521), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n665), .B1(new_n522), .B2(new_n523), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n654), .A2(G15gat), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n529), .ZN(new_n669));
  AOI21_X1  g468(.A(G15gat), .B1(new_n654), .B2(new_n669), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n670), .A2(KEYINPUT104), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(KEYINPUT104), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n668), .B1(new_n671), .B2(new_n672), .ZN(G1326gat));
  NOR2_X1   g472(.A1(new_n651), .A2(new_n317), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G22gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  NAND2_X1  g476(.A1(new_n646), .A2(new_n647), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n528), .A2(new_n540), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n254), .A2(new_n256), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT93), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n257), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n579), .A2(new_n641), .ZN(new_n684));
  AND4_X1   g483(.A1(new_n678), .A2(new_n679), .A3(new_n683), .A4(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n685), .A2(new_n203), .A3(new_n526), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT45), .ZN(new_n687));
  INV_X1    g486(.A(new_n667), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n492), .A2(new_n527), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n540), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n678), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n679), .A2(KEYINPUT44), .A3(new_n678), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n693), .A2(new_n680), .A3(new_n684), .A4(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(G29gat), .B1(new_n695), .B2(new_n525), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n687), .A2(new_n696), .ZN(G1328gat));
  NAND3_X1  g496(.A1(new_n685), .A2(new_n204), .A3(new_n470), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n698), .A2(KEYINPUT46), .ZN(new_n699));
  OAI21_X1  g498(.A(G36gat), .B1(new_n695), .B2(new_n537), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(KEYINPUT46), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(G1329gat));
  OAI21_X1  g501(.A(G43gat), .B1(new_n695), .B2(new_n688), .ZN(new_n703));
  INV_X1    g502(.A(G43gat), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n685), .A2(new_n704), .A3(new_n669), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT47), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n709), .B1(new_n695), .B2(new_n688), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n611), .B1(new_n689), .B2(new_n540), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(KEYINPUT44), .ZN(new_n712));
  AOI211_X1 g511(.A(new_n692), .B(new_n611), .C1(new_n528), .C2(new_n540), .ZN(new_n713));
  INV_X1    g512(.A(new_n684), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n715), .A2(KEYINPUT107), .A3(new_n680), .A4(new_n667), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n710), .A2(new_n716), .A3(G43gat), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n705), .A2(KEYINPUT47), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n708), .B1(new_n717), .B2(new_n718), .ZN(G1330gat));
  OAI21_X1  g518(.A(G50gat), .B1(new_n695), .B2(new_n317), .ZN(new_n720));
  INV_X1    g519(.A(G50gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n685), .A2(new_n721), .A3(new_n316), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT48), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(KEYINPUT108), .B1(new_n695), .B2(new_n317), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n715), .A2(new_n727), .A3(new_n316), .A4(new_n680), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n726), .A2(new_n728), .A3(G50gat), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n722), .A2(KEYINPUT48), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n725), .B1(new_n729), .B2(new_n730), .ZN(G1331gat));
  INV_X1    g530(.A(new_n680), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n648), .A2(new_n642), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n690), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n526), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(new_n553), .ZN(G1332gat));
  XNOR2_X1  g537(.A(new_n734), .B(KEYINPUT109), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n537), .ZN(new_n740));
  NOR2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  AND2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(new_n740), .B2(new_n741), .ZN(G1333gat));
  NAND3_X1  g543(.A1(new_n736), .A2(G71gat), .A3(new_n667), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(G71gat), .B1(new_n736), .B2(new_n669), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT50), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n739), .A2(new_n529), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n749), .B(new_n745), .C1(new_n750), .C2(G71gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n751), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n316), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g553(.A1(new_n579), .A2(new_n642), .A3(new_n680), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n694), .B(new_n755), .C1(KEYINPUT44), .C2(new_n711), .ZN(new_n756));
  INV_X1    g555(.A(G85gat), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n756), .A2(new_n757), .A3(new_n525), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n579), .A2(new_n680), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT110), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n690), .A2(new_n678), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n760), .A2(KEYINPUT110), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n762), .B(new_n764), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n765), .A2(new_n641), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n526), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n758), .B1(new_n767), .B2(new_n757), .ZN(G1336gat));
  NOR2_X1   g567(.A1(new_n537), .A2(G92gat), .ZN(new_n769));
  INV_X1    g568(.A(new_n761), .ZN(new_n770));
  AOI211_X1 g569(.A(new_n611), .B(new_n770), .C1(new_n689), .C2(new_n540), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n763), .B1(new_n771), .B2(new_n759), .ZN(new_n772));
  AND4_X1   g571(.A1(new_n711), .A2(new_n763), .A3(new_n759), .A4(new_n761), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n641), .B(new_n769), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(G92gat), .B1(new_n756), .B2(new_n537), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(KEYINPUT111), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n774), .B(new_n775), .C1(KEYINPUT111), .C2(KEYINPUT52), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(G1337gat));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n583), .A3(new_n669), .ZN(new_n782));
  OAI21_X1  g581(.A(G99gat), .B1(new_n756), .B2(new_n688), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(G1338gat));
  OAI211_X1 g583(.A(KEYINPUT53), .B(G106gat), .C1(new_n756), .C2(new_n317), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n317), .A2(G106gat), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n641), .B(new_n786), .C1(new_n772), .C2(new_n773), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n785), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n712), .A2(new_n713), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n792), .A2(KEYINPUT113), .A3(new_n316), .A4(new_n755), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(new_n756), .B2(new_n317), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n793), .A2(new_n795), .A3(G106gat), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n765), .A2(new_n788), .A3(new_n641), .A4(new_n786), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n791), .B1(new_n798), .B2(new_n789), .ZN(G1339gat));
  NAND2_X1  g598(.A1(new_n575), .A2(new_n578), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n801));
  OR3_X1    g600(.A1(new_n624), .A2(new_n801), .A3(new_n637), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n624), .B2(new_n637), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n629), .A2(new_n802), .A3(KEYINPUT54), .A4(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n633), .B1(new_n638), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n804), .A2(KEYINPUT55), .A3(new_n806), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n809), .A2(new_n636), .A3(new_n680), .A4(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n242), .A2(new_n235), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n244), .A2(new_n245), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n252), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n256), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n641), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n678), .B1(new_n811), .B2(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n809), .A2(new_n636), .A3(new_n810), .A4(new_n815), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n611), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n800), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n579), .A2(new_n611), .A3(new_n642), .A4(new_n732), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n822), .A2(new_n530), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n470), .A2(new_n525), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n326), .A3(new_n680), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n825), .A2(new_n683), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n826), .B1(new_n827), .B2(new_n326), .ZN(G1340gat));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n641), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g629(.A1(new_n825), .A2(new_n579), .ZN(new_n831));
  INV_X1    g630(.A(G127gat), .ZN(new_n832));
  OR3_X1    g631(.A1(new_n831), .A2(KEYINPUT115), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT115), .B1(new_n831), .B2(new_n832), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(G1342gat));
  NOR2_X1   g635(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(G134gat), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n823), .A2(new_n839), .A3(new_n678), .A4(new_n824), .ZN(new_n840));
  AND2_X1   g639(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n840), .A2(new_n838), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n823), .A2(new_n678), .A3(new_n824), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(KEYINPUT117), .A3(G134gat), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT117), .B1(new_n844), .B2(G134gat), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n842), .B(new_n843), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT118), .ZN(new_n849));
  INV_X1    g648(.A(new_n847), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n845), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n851), .A2(new_n852), .A3(new_n842), .A4(new_n843), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n849), .A2(new_n853), .ZN(G1343gat));
  NAND3_X1  g653(.A1(new_n809), .A2(new_n636), .A3(new_n810), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n816), .B1(new_n260), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n611), .ZN(new_n857));
  INV_X1    g656(.A(new_n819), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n579), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n821), .ZN(new_n860));
  OAI211_X1 g659(.A(KEYINPUT57), .B(new_n316), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT119), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n683), .A2(new_n636), .A3(new_n809), .A4(new_n810), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n678), .B1(new_n864), .B2(new_n816), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n800), .B1(new_n865), .B2(new_n819), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n821), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n867), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n316), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n317), .B1(new_n820), .B2(new_n821), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n863), .A2(new_n868), .A3(new_n872), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n667), .A2(new_n525), .A3(new_n470), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n683), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n263), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n869), .A2(new_n526), .A3(new_n688), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT120), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n260), .A2(G141gat), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n869), .A2(new_n880), .A3(new_n526), .A4(new_n688), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n878), .A2(new_n537), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT58), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT121), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n876), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n883), .A2(KEYINPUT121), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n870), .A2(new_n667), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n888), .A2(new_n824), .A3(new_n879), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n873), .A2(new_n680), .A3(new_n874), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(new_n263), .ZN(new_n891));
  OAI22_X1  g690(.A1(new_n886), .A2(new_n887), .B1(new_n891), .B2(new_n883), .ZN(G1344gat));
  NOR2_X1   g691(.A1(new_n642), .A2(G148gat), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n878), .A2(new_n537), .A3(new_n881), .A4(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n870), .A2(KEYINPUT57), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n643), .A2(new_n649), .A3(new_n260), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n871), .B(new_n316), .C1(new_n897), .C2(new_n859), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n896), .A2(new_n898), .A3(new_n641), .A4(new_n874), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n899), .A2(KEYINPUT122), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n264), .B1(new_n899), .B2(KEYINPUT122), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n895), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n873), .A2(new_n641), .A3(new_n874), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n903), .A2(new_n895), .A3(G148gat), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n894), .B1(new_n902), .B2(new_n904), .ZN(G1345gat));
  AND2_X1   g704(.A1(new_n873), .A2(new_n874), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n800), .A2(new_n273), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n878), .A2(new_n579), .A3(new_n537), .A4(new_n881), .ZN(new_n908));
  AOI22_X1  g707(.A1(new_n906), .A2(new_n907), .B1(new_n273), .B2(new_n908), .ZN(G1346gat));
  NOR2_X1   g708(.A1(new_n611), .A2(new_n274), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n878), .A2(new_n678), .A3(new_n537), .A4(new_n881), .ZN(new_n911));
  AOI22_X1  g710(.A1(new_n906), .A2(new_n910), .B1(new_n274), .B2(new_n911), .ZN(G1347gat));
  NAND2_X1  g711(.A1(new_n470), .A2(new_n525), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n823), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n407), .A3(new_n680), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n915), .A2(new_n683), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(new_n407), .ZN(G1348gat));
  NAND2_X1  g717(.A1(new_n915), .A2(new_n641), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g719(.A1(new_n915), .A2(new_n579), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G183gat), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n388), .A2(new_n389), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n823), .A2(new_n579), .A3(new_n923), .A4(new_n914), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT123), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n924), .A2(KEYINPUT123), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n922), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT60), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n922), .A2(new_n929), .A3(new_n926), .A4(new_n925), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1350gat));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n678), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(G190gat), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT124), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n935), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n932), .A2(G190gat), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n936), .B(new_n939), .C1(G190gat), .C2(new_n932), .ZN(G1351gat));
  NAND2_X1  g739(.A1(new_n888), .A2(new_n914), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT125), .ZN(new_n942));
  INV_X1    g741(.A(G197gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(new_n943), .A3(new_n680), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n667), .A2(new_n913), .ZN(new_n945));
  XOR2_X1   g744(.A(new_n945), .B(KEYINPUT126), .Z(new_n946));
  NAND3_X1  g745(.A1(new_n896), .A2(new_n898), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n260), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n944), .A2(new_n948), .ZN(G1352gat));
  NOR3_X1   g748(.A1(new_n941), .A2(G204gat), .A3(new_n642), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n896), .A2(new_n898), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(new_n641), .A3(new_n946), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(G204gat), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n950), .A2(new_n951), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n952), .A2(new_n955), .A3(new_n956), .ZN(G1353gat));
  NAND3_X1  g756(.A1(new_n942), .A2(new_n286), .A3(new_n579), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n953), .A2(new_n579), .A3(new_n945), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n959), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT63), .B1(new_n959), .B2(G211gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(G1354gat));
  AOI21_X1  g761(.A(new_n611), .B1(new_n947), .B2(KEYINPUT127), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n963), .B1(KEYINPUT127), .B2(new_n947), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G218gat), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n942), .A2(new_n287), .A3(new_n678), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(G1355gat));
endmodule


