//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT26), .B(G101), .Z(new_n188));
  NOR2_X1   g002(.A1(G237), .A2(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G137), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT66), .B1(new_n197), .B2(G134), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT11), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n196), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT66), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n201), .B(new_n199), .C1(new_n195), .C2(G137), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(G131), .B1(new_n200), .B2(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n201), .B1(new_n195), .B2(G137), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT11), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n206), .A2(new_n207), .A3(new_n202), .A4(new_n196), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(G146), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT65), .A3(G143), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n212), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  OR2_X1    g031(.A1(new_n217), .A2(KEYINPUT64), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT0), .ZN(new_n219));
  INV_X1    g033(.A(G128), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT64), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n216), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(G143), .B(G146), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n223), .B1(new_n216), .B2(new_n218), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n209), .B(new_n222), .C1(new_n217), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT1), .B1(new_n211), .B2(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G128), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n216), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n223), .A2(new_n229), .A3(G128), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n196), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n195), .A2(G137), .ZN(new_n235));
  OAI21_X1  g049(.A(G131), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n208), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n228), .A2(KEYINPUT68), .A3(new_n230), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n233), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT67), .B(G119), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G116), .ZN(new_n241));
  INV_X1    g055(.A(G119), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n241), .B1(G116), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT2), .B(G113), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n244), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n241), .B(new_n246), .C1(G116), .C2(new_n242), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n225), .A2(new_n239), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT28), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(KEYINPUT71), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n231), .A2(new_n208), .A3(new_n236), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n204), .A2(new_n208), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n222), .B1(new_n224), .B2(new_n217), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n245), .A2(new_n247), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n250), .B1(new_n258), .B2(new_n249), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT71), .B1(new_n249), .B2(new_n250), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n252), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT29), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n194), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n225), .A2(new_n239), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n257), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n250), .B1(new_n265), .B2(new_n249), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n266), .A2(new_n252), .A3(new_n260), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n263), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n249), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT30), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n256), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n225), .A2(new_n239), .A3(KEYINPUT30), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(new_n257), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT69), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n271), .A2(new_n272), .A3(new_n275), .A4(new_n257), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n269), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n193), .A2(KEYINPUT29), .ZN(new_n278));
  AOI21_X1  g092(.A(G902), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n187), .B1(new_n268), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(G472), .A2(G902), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n274), .A2(new_n276), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n249), .A2(new_n193), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT31), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n283), .A2(KEYINPUT31), .A3(new_n285), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT72), .B1(new_n261), .B2(new_n193), .ZN(new_n291));
  INV_X1    g105(.A(new_n259), .ZN(new_n292));
  INV_X1    g106(.A(new_n260), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n293), .A3(new_n251), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n295), .A3(new_n194), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n282), .B1(new_n290), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n280), .B1(KEYINPUT32), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT73), .B1(new_n298), .B2(KEYINPUT32), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n261), .A2(KEYINPUT72), .A3(new_n193), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n295), .B1(new_n294), .B2(new_n194), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT31), .B1(new_n283), .B2(new_n285), .ZN(new_n303));
  AOI211_X1 g117(.A(new_n287), .B(new_n284), .C1(new_n274), .C2(new_n276), .ZN(new_n304));
  OAI22_X1  g118(.A1(new_n301), .A2(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n281), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT32), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n299), .A2(new_n300), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT74), .B(G217), .ZN(new_n311));
  INV_X1    g125(.A(G902), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n311), .B1(G234), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT25), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT23), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n240), .B2(G128), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n242), .A2(new_n220), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n318), .B1(new_n240), .B2(new_n220), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n317), .B1(new_n319), .B2(new_n316), .ZN(new_n320));
  XOR2_X1   g134(.A(KEYINPUT24), .B(G110), .Z(new_n321));
  OAI22_X1  g135(.A1(new_n320), .A2(G110), .B1(new_n321), .B2(new_n319), .ZN(new_n322));
  INV_X1    g136(.A(G140), .ZN(new_n323));
  OR2_X1    g137(.A1(KEYINPUT75), .A2(G125), .ZN(new_n324));
  NAND2_X1  g138(.A1(KEYINPUT75), .A2(G125), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(G125), .A2(G140), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT16), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT75), .B(G125), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT16), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(new_n323), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(G146), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT77), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n328), .A2(new_n334), .A3(G146), .A4(new_n331), .ZN(new_n335));
  XOR2_X1   g149(.A(G125), .B(G140), .Z(new_n336));
  OR2_X1    g150(.A1(new_n336), .A2(G146), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n322), .A2(new_n333), .A3(new_n335), .A4(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n327), .B1(new_n329), .B2(G140), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n331), .B1(new_n339), .B2(new_n330), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n214), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n332), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT76), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n320), .A2(G110), .B1(new_n321), .B2(new_n319), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n343), .B1(new_n342), .B2(new_n344), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n338), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT22), .B(G137), .ZN(new_n348));
  INV_X1    g162(.A(G953), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n349), .A2(G221), .A3(G234), .ZN(new_n350));
  XOR2_X1   g164(.A(new_n348), .B(new_n350), .Z(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n338), .B(new_n351), .C1(new_n345), .C2(new_n346), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n315), .B1(new_n355), .B2(G902), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n353), .A2(KEYINPUT25), .A3(new_n312), .A4(new_n354), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n314), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n355), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n313), .A2(G902), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n310), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G221), .ZN(new_n363));
  XNOR2_X1  g177(.A(KEYINPUT9), .B(G234), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n363), .B1(new_n365), .B2(new_n312), .ZN(new_n366));
  XOR2_X1   g180(.A(KEYINPUT83), .B(G469), .Z(new_n367));
  XNOR2_X1  g181(.A(G110), .B(G140), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n349), .A2(G227), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G107), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(G104), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(KEYINPUT3), .ZN(new_n374));
  INV_X1    g188(.A(G104), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(G107), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n372), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G101), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT78), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(KEYINPUT78), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n371), .A2(G104), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n377), .A2(new_n378), .A3(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(G101), .B1(new_n376), .B2(new_n372), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(new_n228), .A3(new_n230), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n226), .A2(G128), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n230), .B1(new_n223), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n384), .A3(new_n385), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n209), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT12), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(KEYINPUT12), .A3(new_n209), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n373), .A2(KEYINPUT3), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n374), .B1(new_n376), .B2(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n379), .A2(new_n371), .A3(KEYINPUT78), .A4(G104), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n375), .A2(G107), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n396), .B(G101), .C1(new_n398), .C2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT79), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n377), .A2(new_n383), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n405), .A2(KEYINPUT79), .A3(new_n396), .A4(G101), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n255), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n405), .A2(G101), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(KEYINPUT4), .A3(new_n384), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT10), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n386), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(new_n233), .A3(new_n238), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n390), .A2(new_n412), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT80), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n204), .A2(new_n416), .A3(new_n208), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n416), .B1(new_n204), .B2(new_n208), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n411), .A2(new_n414), .A3(new_n415), .A4(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT81), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n238), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT68), .B1(new_n228), .B2(new_n230), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n425), .A2(new_n413), .B1(new_n412), .B2(new_n390), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n426), .A2(KEYINPUT81), .A3(new_n411), .A4(new_n419), .ZN(new_n427));
  AOI221_X4 g241(.A(new_n370), .B1(new_n394), .B2(new_n395), .C1(new_n422), .C2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n370), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n422), .A2(new_n427), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n254), .B1(new_n426), .B2(new_n411), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n429), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n312), .B(new_n367), .C1(new_n428), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT84), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n430), .A2(new_n429), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n394), .A2(new_n395), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n431), .B1(new_n422), .B2(new_n427), .ZN(new_n439));
  OAI22_X1  g253(.A1(new_n436), .A2(new_n438), .B1(new_n439), .B2(new_n429), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT84), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n440), .A2(new_n441), .A3(new_n312), .A4(new_n367), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n435), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n429), .B1(new_n430), .B2(new_n437), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT82), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n431), .B1(new_n436), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n370), .B1(new_n422), .B2(new_n427), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT82), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n444), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(G469), .B1(new_n449), .B2(G902), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n366), .B1(new_n443), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G214), .B1(G237), .B2(G902), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n407), .A2(new_n257), .A3(new_n410), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT85), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT5), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n240), .A2(new_n455), .A3(G116), .ZN(new_n456));
  OAI211_X1 g270(.A(G113), .B(new_n456), .C1(new_n243), .C2(new_n455), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n247), .ZN(new_n458));
  OR2_X1    g272(.A1(new_n458), .A2(new_n386), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT85), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n407), .A2(new_n460), .A3(new_n257), .A4(new_n410), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n454), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(G110), .B(G122), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n454), .A2(new_n459), .A3(new_n463), .A4(new_n461), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(KEYINPUT6), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n462), .A2(new_n468), .A3(new_n464), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n231), .A2(new_n324), .A3(new_n325), .ZN(new_n470));
  INV_X1    g284(.A(new_n329), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n470), .B1(new_n255), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n349), .A2(G224), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT86), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n472), .B(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n467), .A2(new_n469), .A3(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n458), .B(new_n386), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n463), .B(KEYINPUT8), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n474), .A2(KEYINPUT7), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n472), .A2(new_n479), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n477), .A2(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(G902), .B1(new_n482), .B2(new_n466), .ZN(new_n483));
  OAI21_X1  g297(.A(G210), .B1(G237), .B2(G902), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n476), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n484), .B1(new_n476), .B2(new_n483), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n452), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT87), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n476), .A2(new_n483), .ZN(new_n489));
  INV_X1    g303(.A(new_n484), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n476), .A2(new_n483), .A3(new_n484), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT87), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n494), .A3(new_n452), .ZN(new_n495));
  NOR2_X1   g309(.A1(G475), .A2(G902), .ZN(new_n496));
  XNOR2_X1  g310(.A(G113), .B(G122), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(new_n375), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n339), .A2(KEYINPUT19), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n499), .B(new_n214), .C1(KEYINPUT19), .C2(new_n336), .ZN(new_n500));
  INV_X1    g314(.A(G237), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n349), .A3(G214), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n211), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n189), .A2(G143), .A3(G214), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G131), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n503), .A2(new_n207), .A3(new_n504), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n333), .A2(new_n500), .A3(new_n335), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n339), .A2(G146), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n337), .ZN(new_n511));
  NAND2_X1  g325(.A1(KEYINPUT18), .A2(G131), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n503), .A2(new_n504), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n505), .A2(KEYINPUT18), .A3(G131), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n511), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n498), .B1(new_n509), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n505), .A2(KEYINPUT17), .A3(G131), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n506), .A2(new_n518), .A3(new_n507), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n341), .A2(new_n332), .A3(new_n517), .A4(new_n519), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n520), .A2(new_n498), .A3(new_n515), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n496), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n525), .B1(KEYINPUT20), .B2(new_n522), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n498), .B1(new_n520), .B2(new_n515), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n312), .B1(new_n521), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(G475), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(G234), .A2(G237), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(G952), .A3(new_n349), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT21), .B(G898), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n531), .A2(G902), .A3(G953), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G116), .B(G122), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(new_n371), .ZN(new_n539));
  XNOR2_X1  g353(.A(G128), .B(G143), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n195), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n220), .A2(G143), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n542), .A2(KEYINPUT13), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(KEYINPUT13), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n211), .A2(G128), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n539), .B(new_n541), .C1(new_n546), .C2(new_n195), .ZN(new_n547));
  INV_X1    g361(.A(G122), .ZN(new_n548));
  OR3_X1    g362(.A1(new_n548), .A2(KEYINPUT14), .A3(G116), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT14), .B1(new_n548), .B2(G116), .ZN(new_n550));
  INV_X1    g364(.A(G116), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n549), .B(new_n550), .C1(new_n551), .C2(G122), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(G107), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n538), .A2(new_n371), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n540), .B(new_n195), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n547), .A2(new_n556), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n311), .A2(new_n364), .A3(G953), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n547), .A2(new_n556), .A3(new_n558), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n312), .ZN(new_n563));
  INV_X1    g377(.A(G478), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(KEYINPUT15), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n562), .B(new_n312), .C1(KEYINPUT15), .C2(new_n564), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n530), .A2(new_n537), .A3(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n451), .A2(new_n488), .A3(new_n495), .A4(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n362), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(new_n378), .ZN(G3));
  INV_X1    g386(.A(new_n451), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n288), .A2(new_n289), .B1(new_n291), .B2(new_n296), .ZN(new_n574));
  OAI21_X1  g388(.A(G472), .B1(new_n574), .B2(G902), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(new_n361), .A3(new_n306), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n487), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n563), .A2(new_n564), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT33), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n562), .A2(new_n580), .ZN(new_n581));
  OR2_X1    g395(.A1(new_n581), .A2(KEYINPUT89), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n561), .A2(KEYINPUT90), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n561), .A2(KEYINPUT90), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n583), .A2(KEYINPUT33), .A3(new_n560), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n581), .A2(KEYINPUT89), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n582), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n312), .A2(G478), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n579), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n530), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n578), .A2(new_n536), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n577), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT34), .B(G104), .Z(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(G6));
  OAI211_X1 g410(.A(new_n523), .B(new_n496), .C1(new_n516), .C2(new_n521), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n525), .A2(new_n597), .B1(new_n528), .B2(G475), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n536), .B(KEYINPUT91), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n598), .A2(new_n568), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n578), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n577), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT35), .B(G107), .Z(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G9));
  NAND3_X1  g419(.A1(new_n451), .A2(new_n488), .A3(new_n495), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n575), .A2(new_n306), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n356), .A2(new_n357), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n313), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n347), .B1(KEYINPUT36), .B2(new_n352), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n352), .A2(KEYINPUT36), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n338), .B(new_n611), .C1(new_n345), .C2(new_n346), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n610), .A2(new_n360), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT92), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n609), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n569), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n606), .A2(new_n607), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT37), .B(G110), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G12));
  AOI21_X1  g434(.A(new_n487), .B1(new_n609), .B2(new_n615), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n310), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n525), .A2(new_n597), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n532), .B(KEYINPUT93), .Z(new_n624));
  OAI21_X1  g438(.A(new_n624), .B1(G900), .B2(new_n535), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n623), .A2(new_n529), .A3(new_n568), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT94), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT94), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n598), .A2(new_n628), .A3(new_n568), .A4(new_n625), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  AOI211_X1 g444(.A(new_n366), .B(new_n630), .C1(new_n443), .C2(new_n450), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n622), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G128), .ZN(G30));
  XNOR2_X1  g447(.A(new_n625), .B(KEYINPUT39), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n451), .A2(new_n634), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n635), .A2(KEYINPUT40), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n493), .B(KEYINPUT38), .ZN(new_n637));
  INV_X1    g451(.A(new_n265), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n194), .B1(new_n638), .B2(new_n269), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n286), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n187), .B1(new_n640), .B2(new_n312), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n298), .B2(KEYINPUT32), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n300), .A2(new_n642), .A3(new_n309), .ZN(new_n643));
  INV_X1    g457(.A(new_n452), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n526), .A2(new_n529), .ZN(new_n645));
  INV_X1    g459(.A(new_n568), .ZN(new_n646));
  NOR4_X1   g460(.A1(new_n616), .A2(new_n644), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n637), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n635), .A2(KEYINPUT40), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n636), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT95), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n636), .A2(new_n648), .A3(KEYINPUT95), .A4(new_n649), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(new_n211), .ZN(G45));
  NAND3_X1  g469(.A1(new_n589), .A2(new_n530), .A3(new_n625), .ZN(new_n656));
  AOI211_X1 g470(.A(new_n366), .B(new_n656), .C1(new_n443), .C2(new_n450), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n622), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G146), .ZN(G48));
  NAND2_X1  g473(.A1(new_n359), .A2(new_n360), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n609), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n307), .B1(new_n306), .B2(new_n308), .ZN(new_n662));
  AOI211_X1 g476(.A(KEYINPUT73), .B(KEYINPUT32), .C1(new_n305), .C2(new_n281), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n661), .B1(new_n664), .B2(new_n299), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n430), .A2(new_n432), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n370), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n447), .A2(new_n437), .ZN(new_n668));
  AOI21_X1  g482(.A(G902), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(G469), .ZN(new_n670));
  OAI21_X1  g484(.A(KEYINPUT96), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n440), .A2(new_n312), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT96), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n672), .A2(new_n673), .A3(G469), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT97), .ZN(new_n676));
  INV_X1    g490(.A(new_n366), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n675), .A2(new_n676), .A3(new_n677), .A4(new_n443), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n675), .A2(new_n677), .A3(new_n443), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT97), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n665), .A2(new_n593), .A3(new_n678), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  NAND4_X1  g497(.A1(new_n665), .A2(new_n602), .A3(new_n678), .A4(new_n680), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G116), .ZN(G18));
  AOI21_X1  g499(.A(new_n617), .B1(new_n664), .B2(new_n299), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n686), .A2(new_n578), .A3(new_n678), .A4(new_n680), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G119), .ZN(G21));
  NOR2_X1   g502(.A1(new_n267), .A2(new_n193), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n288), .B2(new_n289), .ZN(new_n690));
  OAI21_X1  g504(.A(KEYINPUT98), .B1(new_n690), .B2(new_n282), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT98), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n303), .A2(new_n304), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n692), .B(new_n281), .C1(new_n693), .C2(new_n689), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n575), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n661), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n646), .B1(new_n526), .B2(new_n529), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n452), .B(new_n697), .C1(new_n485), .C2(new_n486), .ZN(new_n698));
  INV_X1    g512(.A(new_n599), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n680), .A2(new_n696), .A3(new_n678), .A4(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT99), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n548), .ZN(G24));
  NAND4_X1  g518(.A1(new_n575), .A2(new_n691), .A3(new_n616), .A4(new_n694), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n656), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n706), .A2(new_n680), .A3(new_n578), .A4(new_n678), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G125), .ZN(G27));
  NAND3_X1  g522(.A1(new_n491), .A2(new_n452), .A3(new_n492), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT101), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT101), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n491), .A2(new_n711), .A3(new_n452), .A4(new_n492), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT100), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n435), .A2(new_n442), .ZN(new_n715));
  INV_X1    g529(.A(new_n448), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n432), .B1(new_n447), .B2(KEYINPUT82), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n438), .B1(new_n422), .B2(new_n427), .ZN(new_n718));
  OAI22_X1  g532(.A1(new_n716), .A2(new_n717), .B1(new_n718), .B2(new_n429), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n670), .B1(new_n719), .B2(new_n312), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n714), .B1(new_n715), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n443), .A2(new_n450), .A3(KEYINPUT100), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n713), .A2(new_n677), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n306), .A2(new_n308), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n661), .B1(new_n299), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n656), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(KEYINPUT42), .B1(new_n723), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n710), .A2(new_n677), .A3(new_n712), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n443), .A2(new_n450), .A3(KEYINPUT100), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT100), .B1(new_n443), .B2(new_n450), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n656), .A2(KEYINPUT42), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(new_n665), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n728), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n207), .ZN(G33));
  INV_X1    g550(.A(new_n630), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n732), .A2(new_n665), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G134), .ZN(G36));
  INV_X1    g553(.A(KEYINPUT45), .ZN(new_n740));
  OR3_X1    g554(.A1(new_n719), .A2(KEYINPUT102), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(KEYINPUT102), .B1(new_n719), .B2(new_n740), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n670), .B1(new_n719), .B2(new_n740), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(G469), .A2(G902), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(KEYINPUT46), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT46), .B1(new_n744), .B2(new_n745), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT103), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n443), .B(new_n746), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n677), .B(new_n634), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n751), .A2(KEYINPUT104), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(KEYINPUT104), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n645), .A2(new_n589), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT43), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n755), .A2(KEYINPUT43), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n607), .A2(new_n616), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n759), .A2(KEYINPUT44), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(KEYINPUT44), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n713), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n754), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G137), .ZN(G39));
  OAI21_X1  g579(.A(new_n677), .B1(new_n749), .B2(new_n750), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT47), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g582(.A(KEYINPUT47), .B(new_n677), .C1(new_n749), .C2(new_n750), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n713), .ZN(new_n771));
  NOR4_X1   g585(.A1(new_n771), .A2(new_n310), .A3(new_n361), .A4(new_n656), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G140), .ZN(G42));
  AND2_X1   g588(.A1(new_n675), .A2(new_n443), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT49), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n637), .A2(new_n366), .A3(new_n644), .A4(new_n755), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n664), .A2(new_n361), .A3(new_n642), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT105), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n680), .A2(new_n678), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n771), .ZN(new_n783));
  INV_X1    g597(.A(new_n532), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n784), .A3(new_n779), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n785), .A2(new_n530), .A3(new_n589), .ZN(new_n786));
  INV_X1    g600(.A(new_n624), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n757), .A2(new_n787), .A3(new_n756), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT111), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n705), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(new_n783), .A3(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(new_n793), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n786), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n696), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n789), .A2(new_n637), .A3(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n680), .A2(KEYINPUT112), .A3(new_n644), .A4(new_n678), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n801), .B1(new_n782), .B2(new_n452), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT50), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  AND4_X1   g617(.A1(KEYINPUT50), .A2(new_n798), .A3(new_n802), .A4(new_n799), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n796), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n775), .A2(new_n366), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n768), .A2(new_n769), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n789), .A2(new_n797), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n807), .A2(new_n713), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT110), .B1(new_n805), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT51), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n790), .A2(new_n783), .A3(new_n725), .ZN(new_n812));
  NOR2_X1   g626(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n813));
  AND2_X1   g627(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n349), .A2(G952), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n680), .A2(new_n578), .A3(new_n678), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n816), .B1(new_n808), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(new_n590), .B2(new_n785), .ZN(new_n820));
  AOI211_X1 g634(.A(new_n815), .B(new_n820), .C1(new_n812), .C2(new_n813), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n811), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT108), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n609), .A2(new_n677), .A3(new_n615), .A4(new_n625), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n698), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n643), .A2(new_n721), .A3(new_n722), .A4(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT109), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n730), .A2(new_n731), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(KEYINPUT109), .A3(new_n643), .A4(new_n826), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n310), .B(new_n621), .C1(new_n631), .C2(new_n657), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n833), .A2(new_n707), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT52), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n829), .A2(new_n831), .A3(new_n833), .A4(new_n707), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n824), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n680), .A2(new_n310), .A3(new_n361), .A4(new_n678), .ZN(new_n841));
  INV_X1    g655(.A(new_n617), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n310), .A2(new_n842), .ZN(new_n843));
  OAI22_X1  g657(.A1(new_n841), .A2(new_n601), .B1(new_n817), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n841), .A2(new_n592), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n187), .B1(new_n305), .B2(new_n312), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n846), .A2(new_n661), .A3(new_n298), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n530), .A2(new_n646), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT106), .ZN(new_n849));
  AOI22_X1  g663(.A1(new_n848), .A2(new_n849), .B1(new_n530), .B2(new_n589), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT106), .B1(new_n530), .B2(new_n646), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n699), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n846), .A2(new_n298), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n847), .A2(new_n852), .B1(new_n842), .B2(new_n853), .ZN(new_n854));
  OAI22_X1  g668(.A1(new_n854), .A2(new_n606), .B1(new_n362), .B2(new_n570), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n844), .A2(new_n845), .A3(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n728), .A2(new_n734), .A3(new_n738), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n701), .B(KEYINPUT99), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n646), .A2(new_n625), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(KEYINPUT107), .A3(new_n598), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n613), .B(KEYINPUT92), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n860), .B1(new_n861), .B2(new_n358), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT107), .B1(new_n859), .B2(new_n598), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n451), .A2(new_n864), .A3(new_n712), .A4(new_n710), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n732), .A2(new_n706), .B1(new_n865), .B2(new_n310), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n856), .A2(new_n857), .A3(new_n858), .A4(new_n866), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n836), .B(KEYINPUT52), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n839), .B(new_n840), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n866), .A2(new_n728), .A3(new_n734), .A4(new_n738), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n451), .A2(new_n488), .A3(new_n495), .A4(new_n569), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n451), .A2(new_n488), .A3(new_n495), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n645), .A2(new_n849), .A3(new_n568), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(new_n590), .A3(new_n851), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n599), .ZN(new_n875));
  OAI22_X1  g689(.A1(new_n576), .A2(new_n875), .B1(new_n607), .B2(new_n617), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n665), .A2(new_n871), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n877), .A2(new_n681), .A3(new_n684), .A4(new_n687), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n870), .A2(new_n878), .A3(new_n703), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n832), .A2(new_n834), .A3(KEYINPUT52), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n836), .A2(new_n837), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n879), .B(new_n882), .C1(new_n824), .C2(KEYINPUT53), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n823), .B1(new_n869), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT53), .B1(new_n867), .B2(new_n868), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n879), .A2(new_n840), .A3(new_n882), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT54), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n810), .A2(KEYINPUT51), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n822), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(G952), .A2(G953), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n781), .B1(new_n890), .B2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n878), .A2(new_n703), .ZN(new_n893));
  INV_X1    g707(.A(new_n870), .ZN(new_n894));
  AND4_X1   g708(.A1(new_n840), .A2(new_n882), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n840), .B1(new_n879), .B2(new_n882), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(G210), .A3(G902), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n467), .A2(new_n469), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(new_n475), .Z(new_n901));
  XOR2_X1   g715(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n902));
  XNOR2_X1  g716(.A(new_n901), .B(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n898), .A2(new_n899), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n903), .B1(new_n898), .B2(new_n899), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n349), .A2(G952), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(G51));
  OAI21_X1  g721(.A(new_n823), .B1(new_n895), .B2(new_n896), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n885), .A2(KEYINPUT54), .A3(new_n886), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n745), .B(KEYINPUT57), .Z(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n440), .ZN(new_n913));
  OR4_X1    g727(.A1(new_n312), .A2(new_n895), .A3(new_n896), .A4(new_n744), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n906), .B1(new_n913), .B2(new_n914), .ZN(G54));
  NAND4_X1  g729(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n516), .A2(new_n521), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n916), .A2(new_n918), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n919), .A2(new_n920), .A3(new_n906), .ZN(G60));
  XNOR2_X1  g735(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n564), .A2(new_n312), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n922), .B(new_n923), .Z(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n884), .B2(new_n887), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n587), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n587), .A2(new_n924), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n906), .B1(new_n910), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT117), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT117), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n927), .A2(new_n929), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(G63));
  XOR2_X1   g748(.A(KEYINPUT118), .B(KEYINPUT60), .Z(new_n935));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n935), .B(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n885), .A2(new_n886), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n355), .ZN(new_n939));
  INV_X1    g753(.A(new_n906), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n610), .A2(new_n612), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n885), .A2(new_n942), .A3(new_n886), .A4(new_n937), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n939), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT120), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT119), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n938), .A2(new_n948), .A3(new_n355), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n938), .B2(new_n355), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n943), .A2(KEYINPUT61), .A3(new_n940), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n947), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n939), .A2(KEYINPUT119), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n938), .A2(new_n948), .A3(new_n355), .ZN(new_n955));
  AND4_X1   g769(.A1(new_n947), .A2(new_n952), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n946), .B1(new_n953), .B2(new_n956), .ZN(G66));
  NAND3_X1  g771(.A1(new_n534), .A2(G224), .A3(G953), .ZN(new_n958));
  INV_X1    g772(.A(new_n893), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(G953), .ZN(new_n960));
  INV_X1    g774(.A(G898), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n900), .B1(new_n961), .B2(G953), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n960), .B(new_n962), .ZN(G69));
  AOI22_X1  g777(.A1(new_n754), .A2(new_n763), .B1(new_n770), .B2(new_n772), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n652), .A2(new_n653), .A3(new_n834), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT62), .Z(new_n966));
  INV_X1    g780(.A(new_n635), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n665), .A2(new_n967), .A3(new_n713), .A4(new_n874), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n964), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n349), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n271), .A2(new_n272), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT121), .Z(new_n972));
  OAI21_X1  g786(.A(new_n499), .B1(KEYINPUT19), .B2(new_n336), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n972), .B(new_n973), .Z(new_n974));
  NAND2_X1  g788(.A1(new_n970), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n974), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n857), .A2(new_n834), .ZN(new_n977));
  AOI211_X1 g791(.A(new_n661), .B(new_n698), .C1(new_n299), .C2(new_n724), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n977), .B1(new_n754), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(G953), .B1(new_n964), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n349), .A2(G900), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT123), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n976), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n349), .B1(G227), .B2(G900), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT122), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n975), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n985), .B1(new_n975), .B2(new_n983), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n986), .A2(new_n987), .ZN(G72));
  NAND2_X1  g802(.A1(G472), .A2(G902), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT63), .Z(new_n990));
  OAI21_X1  g804(.A(new_n990), .B1(new_n969), .B2(new_n959), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n277), .B(KEYINPUT124), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n991), .A2(new_n193), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n964), .A2(new_n979), .A3(new_n893), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n990), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n992), .A2(new_n193), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT125), .Z(new_n997));
  NAND2_X1  g811(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n869), .A2(new_n883), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n286), .B1(new_n193), .B2(new_n277), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n990), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT126), .Z(new_n1002));
  AOI21_X1  g816(.A(new_n906), .B1(new_n999), .B2(new_n1002), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n993), .A2(new_n998), .A3(new_n1003), .ZN(G57));
endmodule


