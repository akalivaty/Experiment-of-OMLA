//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G104), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(G104), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G101), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(KEYINPUT78), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT78), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G107), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n197), .A3(G104), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT77), .B(KEYINPUT3), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n193), .B(new_n194), .C1(new_n198), .C2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT80), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n189), .A2(KEYINPUT77), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT77), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT3), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT78), .B(G107), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G104), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n208), .A2(KEYINPUT80), .A3(new_n194), .A4(new_n193), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n202), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(G128), .ZN(new_n217));
  INV_X1    g031(.A(G128), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n212), .B(new_n214), .C1(KEYINPUT1), .C2(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n195), .A2(new_n197), .ZN(new_n221));
  INV_X1    g035(.A(G104), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT81), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(G104), .B2(new_n190), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n194), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n221), .A2(new_n224), .A3(new_n222), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n210), .A2(KEYINPUT10), .A3(new_n220), .A4(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT82), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n202), .A2(new_n209), .B1(new_n226), .B2(new_n227), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT82), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n231), .A2(new_n232), .A3(KEYINPUT10), .A4(new_n220), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n193), .B1(new_n198), .B2(new_n199), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G101), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT79), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(KEYINPUT79), .A3(G101), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n210), .A2(new_n238), .A3(KEYINPUT4), .A4(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n236), .A2(KEYINPUT4), .ZN(new_n241));
  XNOR2_X1  g055(.A(G143), .B(G146), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT0), .B(G128), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT64), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AND2_X1   g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT64), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n215), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n244), .A2(new_n246), .A3(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n241), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n210), .A2(new_n220), .A3(new_n228), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT10), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n240), .A2(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT11), .ZN(new_n256));
  INV_X1    g070(.A(G134), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n256), .B1(new_n257), .B2(G137), .ZN(new_n258));
  INV_X1    g072(.A(G137), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT11), .A3(G134), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n257), .A2(G137), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G131), .ZN(new_n263));
  INV_X1    g077(.A(G131), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n258), .A2(new_n260), .A3(new_n264), .A4(new_n261), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n234), .A2(new_n255), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(G110), .B(G140), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n268), .B(KEYINPUT76), .ZN(new_n269));
  INV_X1    g083(.A(G953), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n270), .A2(G227), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n269), .B(new_n271), .Z(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n263), .A2(new_n265), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n210), .A2(new_n220), .A3(new_n228), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n220), .B1(new_n210), .B2(new_n228), .ZN(new_n277));
  OAI211_X1 g091(.A(KEYINPUT12), .B(new_n275), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT83), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT12), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n231), .B(new_n220), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT83), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT12), .A4(new_n275), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n274), .B1(new_n283), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n234), .A2(new_n255), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n275), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n273), .B1(new_n289), .B2(new_n267), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n187), .B(new_n188), .C1(new_n287), .C2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n187), .A2(new_n188), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n286), .A2(new_n279), .A3(new_n282), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n267), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n272), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n267), .A2(new_n273), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n289), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n291), .B(new_n293), .C1(new_n187), .C2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT9), .B(G234), .ZN(new_n301));
  OAI21_X1  g115(.A(G221), .B1(new_n301), .B2(G902), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G214), .B1(G237), .B2(G902), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(G116), .B(G119), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT2), .B(G113), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n308), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n306), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n241), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n240), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G116), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(G119), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT5), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g133(.A(G113), .B(new_n319), .C1(new_n307), .C2(new_n318), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n311), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n231), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n315), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT6), .ZN(new_n325));
  XNOR2_X1  g139(.A(G110), .B(G122), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n315), .A2(new_n323), .A3(new_n326), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT6), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n326), .B1(new_n315), .B2(new_n323), .ZN(new_n331));
  OAI211_X1 g145(.A(KEYINPUT84), .B(new_n328), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n331), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT84), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT6), .A4(new_n329), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n251), .A2(G125), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n337), .B1(G125), .B2(new_n220), .ZN(new_n338));
  INV_X1    g152(.A(G224), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(G953), .ZN(new_n340));
  XOR2_X1   g154(.A(new_n338), .B(new_n340), .Z(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n336), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(G210), .B1(G237), .B2(G902), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT7), .B1(new_n339), .B2(G953), .ZN(new_n345));
  XOR2_X1   g159(.A(new_n338), .B(new_n345), .Z(new_n346));
  AND2_X1   g160(.A1(new_n346), .A2(new_n329), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT85), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n231), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n322), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n231), .A2(new_n348), .A3(new_n321), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n326), .B(KEYINPUT8), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(G902), .B1(new_n347), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n343), .A2(new_n344), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n344), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n341), .B1(new_n332), .B2(new_n335), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n347), .A2(new_n353), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n188), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n356), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n305), .B1(new_n355), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n303), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT91), .ZN(new_n363));
  INV_X1    g177(.A(G237), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(new_n270), .A3(G214), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n213), .ZN(new_n366));
  NOR2_X1   g180(.A1(G237), .A2(G953), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(G143), .A3(G214), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n366), .A2(new_n264), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT87), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT17), .ZN(new_n371));
  INV_X1    g185(.A(new_n368), .ZN(new_n372));
  AOI21_X1  g186(.A(G143), .B1(new_n367), .B2(G214), .ZN(new_n373));
  OAI21_X1  g187(.A(G131), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT87), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n366), .A2(new_n375), .A3(new_n264), .A4(new_n368), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n370), .A2(new_n371), .A3(new_n374), .A4(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G140), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G125), .ZN(new_n379));
  INV_X1    g193(.A(G125), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G140), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT72), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n379), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n378), .A2(KEYINPUT72), .A3(G125), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(KEYINPUT16), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT16), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n379), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n211), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n385), .A2(new_n387), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G146), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n366), .A2(new_n368), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(KEYINPUT17), .A3(G131), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n377), .A2(new_n388), .A3(new_n390), .A4(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G113), .B(G122), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n394), .B(new_n222), .ZN(new_n395));
  NAND2_X1  g209(.A1(KEYINPUT18), .A2(G131), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n366), .A2(new_n368), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n383), .A2(G146), .A3(new_n384), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n379), .A2(new_n381), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n211), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n396), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT86), .B1(new_n391), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT86), .ZN(new_n404));
  AOI211_X1 g218(.A(new_n404), .B(new_n396), .C1(new_n366), .C2(new_n368), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n397), .B(new_n401), .C1(new_n403), .C2(new_n405), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n393), .A2(new_n395), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n370), .A2(new_n374), .A3(new_n376), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT19), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n409), .B1(new_n383), .B2(new_n384), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n399), .A2(KEYINPUT19), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n211), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n408), .A2(new_n390), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n395), .B1(new_n413), .B2(new_n406), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT88), .B1(new_n407), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(G475), .A2(G902), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n413), .A2(new_n406), .ZN(new_n417));
  INV_X1    g231(.A(new_n395), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT88), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n393), .A2(new_n395), .A3(new_n406), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n415), .A2(new_n416), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT89), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT20), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n424), .B1(new_n423), .B2(KEYINPUT20), .ZN(new_n426));
  INV_X1    g240(.A(new_n416), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(KEYINPUT20), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n419), .B2(new_n421), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n425), .A2(new_n426), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n395), .B1(new_n393), .B2(new_n406), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n188), .B1(new_n407), .B2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT90), .B(G475), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n363), .B1(new_n431), .B2(new_n436), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n420), .B1(new_n419), .B2(new_n421), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n438), .A2(new_n439), .A3(new_n427), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT89), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT20), .ZN(new_n443));
  INV_X1    g257(.A(new_n430), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(KEYINPUT91), .A3(new_n435), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n218), .A2(G143), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT13), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT93), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n213), .A2(G128), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n448), .A2(new_n450), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT13), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT93), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n451), .B(G134), .C1(new_n452), .C2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n450), .A2(new_n447), .A3(new_n257), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n316), .A2(G122), .ZN(new_n457));
  INV_X1    g271(.A(G122), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G116), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(new_n459), .A3(KEYINPUT92), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT92), .B1(new_n457), .B2(new_n459), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n461), .A2(new_n462), .A3(new_n207), .ZN(new_n463));
  INV_X1    g277(.A(new_n462), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n221), .B1(new_n464), .B2(new_n460), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n455), .B(new_n456), .C1(new_n463), .C2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT94), .ZN(new_n467));
  INV_X1    g281(.A(new_n456), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n257), .B1(new_n450), .B2(new_n447), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT14), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n457), .A2(new_n459), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(G107), .B1(new_n457), .B2(new_n470), .ZN(new_n472));
  OAI22_X1  g286(.A1(new_n468), .A2(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n467), .B1(new_n465), .B2(new_n473), .ZN(new_n474));
  OR2_X1    g288(.A1(new_n468), .A2(new_n469), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n471), .A2(new_n472), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n207), .B1(new_n461), .B2(new_n462), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n475), .A2(new_n476), .A3(new_n477), .A4(KEYINPUT94), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n466), .A2(new_n474), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G217), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n301), .A2(new_n480), .A3(G953), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n466), .A2(new_n474), .A3(new_n478), .A4(new_n481), .ZN(new_n484));
  AOI21_X1  g298(.A(G902), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G478), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n486), .A2(KEYINPUT15), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n485), .B(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n270), .A2(G952), .ZN(new_n490));
  NAND2_X1  g304(.A1(G234), .A2(G237), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(G902), .A3(G953), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(KEYINPUT95), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT21), .B(G898), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n489), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n437), .A2(new_n446), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT96), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n445), .A2(KEYINPUT91), .A3(new_n435), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT91), .B1(new_n445), .B2(new_n435), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n505), .A2(KEYINPUT96), .A3(new_n499), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n362), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n218), .A2(G119), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n508), .A2(KEYINPUT71), .A3(KEYINPUT23), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT71), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n218), .A2(G119), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT23), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n509), .B1(new_n513), .B2(new_n508), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(KEYINPUT70), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT70), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n516), .B1(new_n218), .B2(G119), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n515), .A2(new_n517), .B1(G119), .B2(new_n218), .ZN(new_n518));
  XOR2_X1   g332(.A(KEYINPUT24), .B(G110), .Z(new_n519));
  AOI22_X1  g333(.A1(new_n514), .A2(G110), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n388), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n211), .B1(new_n385), .B2(new_n387), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT73), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n520), .B(KEYINPUT73), .C1(new_n521), .C2(new_n522), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI22_X1  g341(.A1(new_n514), .A2(G110), .B1(new_n518), .B2(new_n519), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n390), .A3(new_n400), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT22), .B(G137), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n270), .A2(G221), .A3(G234), .ZN(new_n532));
  XOR2_X1   g346(.A(new_n531), .B(new_n532), .Z(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n527), .A2(new_n529), .A3(new_n533), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n188), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT25), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT25), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n535), .A2(new_n536), .A3(new_n539), .A4(new_n188), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n480), .B1(G234), .B2(new_n188), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n541), .A2(G902), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n535), .A2(new_n536), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT74), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n545), .B(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT75), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n545), .B(KEYINPUT74), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT75), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n550), .A3(new_n542), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n367), .A2(G210), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(KEYINPUT27), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT26), .B(G101), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n261), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n257), .A2(G137), .ZN(new_n559));
  OAI21_X1  g373(.A(G131), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n217), .A2(new_n560), .A3(new_n265), .A4(new_n219), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(new_n266), .B2(new_n251), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT65), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT30), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n275), .A2(new_n244), .A3(new_n246), .A4(new_n250), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT30), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT65), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n566), .A2(KEYINPUT65), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n565), .A2(new_n561), .A3(new_n567), .A4(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n312), .B1(new_n564), .B2(new_n570), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n312), .B(new_n561), .C1(new_n266), .C2(new_n251), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n557), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n312), .B1(new_n565), .B2(new_n561), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT28), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT28), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n572), .A2(KEYINPUT66), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n572), .A2(new_n577), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT66), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n576), .A2(new_n556), .A3(new_n578), .A4(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT29), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n574), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT68), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n582), .ZN(new_n587));
  AOI21_X1  g401(.A(G902), .B1(new_n587), .B2(KEYINPUT29), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n574), .A2(new_n582), .A3(KEYINPUT68), .A4(new_n583), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(G472), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT69), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT69), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n590), .A2(new_n593), .A3(G472), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT32), .ZN(new_n596));
  NOR4_X1   g410(.A1(new_n571), .A2(KEYINPUT31), .A3(new_n557), .A4(new_n573), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT31), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n562), .A2(new_n313), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n577), .B1(new_n599), .B2(new_n572), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n572), .A2(KEYINPUT66), .A3(new_n577), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT66), .B1(new_n572), .B2(new_n577), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n598), .B1(new_n603), .B2(new_n556), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n571), .A2(new_n557), .A3(new_n573), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n597), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(G472), .A2(G902), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n596), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n605), .A2(new_n598), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n576), .A2(new_n578), .A3(new_n581), .ZN(new_n612));
  AOI21_X1  g426(.A(KEYINPUT31), .B1(new_n612), .B2(new_n557), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n611), .B1(new_n613), .B2(new_n605), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(KEYINPUT32), .A3(new_n608), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n610), .A2(KEYINPUT67), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n608), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT67), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n617), .A2(new_n618), .A3(new_n596), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n552), .B1(new_n595), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n507), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G101), .ZN(G3));
  AND2_X1   g437(.A1(new_n548), .A2(new_n551), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT97), .ZN(new_n625));
  OAI21_X1  g439(.A(G472), .B1(new_n607), .B2(G902), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n626), .A2(new_n617), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n303), .A2(new_n624), .A3(new_n625), .A4(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n548), .A2(new_n627), .A3(new_n551), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n300), .A2(new_n302), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT97), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n483), .A2(new_n484), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT98), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT33), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n633), .A2(new_n634), .A3(KEYINPUT33), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n637), .A2(G478), .A3(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT99), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n486), .A2(new_n188), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n485), .B2(new_n486), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n640), .B1(new_n639), .B2(new_n642), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n646), .B1(new_n503), .B2(new_n504), .ZN(new_n647));
  INV_X1    g461(.A(new_n498), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n361), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n632), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT100), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT34), .B(G104), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G6));
  NOR2_X1   g468(.A1(new_n425), .A2(new_n426), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n438), .A2(new_n439), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n428), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n435), .A3(new_n489), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n649), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n632), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT35), .B(G107), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G9));
  NOR2_X1   g477(.A1(new_n534), .A2(KEYINPUT36), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n530), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n544), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n542), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n627), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n507), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  NAND2_X1  g486(.A1(new_n355), .A2(new_n360), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n304), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n630), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n667), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n676), .B1(new_n620), .B2(new_n595), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n658), .ZN(new_n679));
  INV_X1    g493(.A(new_n489), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n492), .B(KEYINPUT101), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(G900), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n682), .B1(new_n683), .B2(new_n496), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n435), .A2(new_n685), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n679), .A2(new_n680), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n678), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  XOR2_X1   g503(.A(KEYINPUT104), .B(KEYINPUT39), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n684), .B(new_n690), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n303), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT40), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n303), .A2(new_n691), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT40), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT105), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n693), .A2(new_n699), .A3(new_n696), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n557), .B1(new_n573), .B2(new_n575), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT102), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n188), .B1(new_n703), .B2(new_n605), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G472), .ZN(new_n705));
  AOI21_X1  g519(.A(KEYINPUT103), .B1(new_n620), .B2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT103), .ZN(new_n707));
  INV_X1    g521(.A(new_n705), .ZN(new_n708));
  AOI211_X1 g522(.A(new_n707), .B(new_n708), .C1(new_n616), .C2(new_n619), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n676), .B1(new_n706), .B2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n673), .B(KEYINPUT38), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n680), .B1(new_n437), .B2(new_n446), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n712), .A2(new_n304), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n698), .A2(new_n700), .A3(new_n711), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G143), .ZN(G45));
  AOI211_X1 g530(.A(new_n684), .B(new_n645), .C1(new_n437), .C2(new_n446), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n678), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT106), .B(G146), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G48));
  NAND2_X1  g534(.A1(new_n289), .A2(new_n267), .ZN(new_n721));
  AOI22_X1  g535(.A1(new_n272), .A2(new_n721), .B1(new_n297), .B2(new_n294), .ZN(new_n722));
  OAI21_X1  g536(.A(G469), .B1(new_n722), .B2(G902), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n302), .A3(new_n291), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT107), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n723), .A2(new_n726), .A3(new_n302), .A4(new_n291), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n650), .A2(new_n621), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT41), .B(G113), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G15));
  NAND3_X1  g545(.A1(new_n621), .A2(new_n660), .A3(new_n728), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G116), .ZN(G18));
  AND3_X1   g547(.A1(new_n725), .A2(new_n361), .A3(new_n727), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT96), .B1(new_n505), .B2(new_n499), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n500), .A2(new_n501), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n734), .B(new_n677), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G119), .ZN(G21));
  INV_X1    g552(.A(new_n649), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n549), .A2(new_n542), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n627), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n728), .A2(new_n739), .A3(new_n713), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  OAI211_X1 g558(.A(new_n646), .B(new_n685), .C1(new_n503), .C2(new_n504), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n668), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n734), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G125), .ZN(G27));
  AOI21_X1  g562(.A(KEYINPUT32), .B1(new_n614), .B2(new_n608), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n615), .B1(new_n749), .B2(KEYINPUT109), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n614), .A2(new_n751), .A3(KEYINPUT32), .A4(new_n608), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n740), .B1(new_n753), .B2(new_n595), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n266), .B1(new_n234), .B2(new_n255), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT108), .B1(new_n274), .B2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n289), .A2(new_n757), .A3(new_n267), .A4(new_n273), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(G469), .A3(new_n296), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n291), .A3(new_n293), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n302), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n355), .A2(new_n304), .A3(new_n360), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT42), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n754), .A2(new_n765), .A3(new_n717), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n620), .A2(new_n595), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n761), .A2(new_n302), .ZN(new_n770));
  INV_X1    g584(.A(new_n763), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n769), .A2(new_n624), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n764), .B1(new_n772), .B2(new_n745), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n754), .A2(new_n765), .A3(new_n717), .A4(KEYINPUT110), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n768), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G131), .ZN(G33));
  NOR2_X1   g590(.A1(new_n762), .A2(new_n763), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n621), .A2(new_n687), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n621), .A2(KEYINPUT111), .A3(new_n687), .A4(new_n777), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G134), .ZN(G36));
  NAND2_X1  g597(.A1(new_n505), .A2(new_n646), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT43), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT112), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n646), .B1(new_n786), .B2(KEYINPUT43), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n787), .B(new_n505), .C1(new_n786), .C2(new_n646), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n627), .A2(new_n676), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n785), .A2(new_n788), .A3(KEYINPUT44), .A4(new_n789), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n790), .A2(KEYINPUT113), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(KEYINPUT113), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n771), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT114), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n791), .A2(new_n795), .A3(new_n771), .A4(new_n792), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n785), .A2(new_n788), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT44), .B1(new_n797), .B2(new_n789), .ZN(new_n798));
  INV_X1    g612(.A(new_n302), .ZN(new_n799));
  INV_X1    g613(.A(new_n291), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT45), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n187), .B1(new_n299), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n759), .A2(KEYINPUT45), .A3(new_n296), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n292), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT46), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n800), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n804), .A2(KEYINPUT46), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n799), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n691), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n798), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n794), .A2(new_n796), .A3(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(KEYINPUT115), .B(G137), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n812), .B(new_n813), .ZN(G39));
  NOR4_X1   g628(.A1(new_n745), .A2(new_n769), .A3(new_n624), .A4(new_n763), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n809), .A2(KEYINPUT47), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n809), .A2(KEYINPUT47), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G140), .ZN(G42));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n797), .A2(new_n682), .A3(new_n742), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(KEYINPUT50), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n728), .A2(new_n305), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n825), .A2(KEYINPUT117), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n712), .B1(new_n825), .B2(KEYINPUT117), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n822), .A2(new_n824), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n728), .A2(new_n771), .ZN(new_n829));
  XOR2_X1   g643(.A(new_n829), .B(KEYINPUT119), .Z(new_n830));
  AOI21_X1  g644(.A(new_n708), .B1(new_n616), .B2(new_n619), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT103), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n832), .A2(new_n552), .A3(new_n492), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n830), .A2(new_n505), .A3(new_n645), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n826), .A2(new_n827), .ZN(new_n835));
  OAI22_X1  g649(.A1(new_n835), .A2(new_n821), .B1(new_n823), .B2(KEYINPUT50), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n797), .A2(new_n682), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n830), .A2(new_n669), .A3(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n828), .A2(new_n834), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n816), .A2(new_n817), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n723), .A2(new_n799), .A3(new_n291), .ZN(new_n841));
  AOI211_X1 g655(.A(new_n763), .B(new_n821), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n820), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n830), .A2(new_n833), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n490), .B1(new_n844), .B2(new_n647), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n734), .B2(new_n822), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n830), .A2(new_n754), .A3(new_n837), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(KEYINPUT48), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n847), .A2(KEYINPUT48), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n843), .B(new_n846), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n675), .B(new_n677), .C1(new_n717), .C2(new_n687), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n747), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n713), .A2(new_n770), .A3(new_n361), .A4(new_n685), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n710), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT52), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n361), .B(new_n489), .C1(new_n504), .C2(new_n503), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n761), .A2(new_n302), .A3(new_n685), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n832), .A2(new_n858), .A3(new_n676), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT52), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n859), .A2(new_n860), .A3(new_n747), .A4(new_n851), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n489), .A2(new_n686), .ZN(new_n863));
  NOR4_X1   g677(.A1(new_n630), .A2(new_n763), .A3(new_n679), .A4(new_n863), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n864), .A2(new_n677), .B1(new_n746), .B2(new_n777), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n782), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n505), .A2(new_n489), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n649), .B1(new_n867), .B2(new_n647), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(new_n628), .A3(new_n631), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n622), .A2(new_n670), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n768), .A2(new_n773), .A3(new_n774), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n621), .B(new_n728), .C1(new_n650), .C2(new_n660), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(new_n737), .A3(new_n743), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n862), .A2(new_n871), .A3(KEYINPUT53), .A4(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n873), .A2(new_n737), .A3(new_n743), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n855), .A2(new_n878), .A3(new_n861), .A4(new_n775), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n632), .A2(new_n868), .B1(new_n507), .B2(new_n621), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n880), .A2(new_n670), .A3(new_n782), .A4(new_n865), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n877), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n876), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT54), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n855), .A2(KEYINPUT53), .A3(new_n861), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT116), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n886), .B1(new_n872), .B2(new_n874), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n878), .A2(KEYINPUT116), .A3(new_n775), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n885), .A2(new_n871), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT54), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(new_n890), .A3(new_n882), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n884), .A2(new_n891), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n839), .A2(new_n842), .A3(new_n820), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n850), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(G952), .A2(G953), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n723), .A2(new_n291), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(KEYINPUT49), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n896), .A2(KEYINPUT49), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n741), .A2(new_n304), .A3(new_n302), .ZN(new_n899));
  NOR4_X1   g713(.A1(new_n712), .A2(new_n897), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n900), .A2(new_n505), .A3(new_n646), .ZN(new_n901));
  OAI22_X1  g715(.A1(new_n894), .A2(new_n895), .B1(new_n832), .B2(new_n901), .ZN(G75));
  NOR2_X1   g716(.A1(new_n270), .A2(G952), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n188), .B1(new_n889), .B2(new_n882), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT56), .B1(new_n905), .B2(G210), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n336), .B(KEYINPUT120), .Z(new_n907));
  XOR2_X1   g721(.A(new_n341), .B(KEYINPUT55), .Z(new_n908));
  XOR2_X1   g722(.A(new_n907), .B(new_n908), .Z(new_n909));
  OAI21_X1  g723(.A(new_n904), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n910), .B1(new_n906), .B2(new_n909), .ZN(G51));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n891), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n889), .A2(new_n882), .A3(KEYINPUT121), .A4(new_n890), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n889), .A2(new_n882), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(KEYINPUT54), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n292), .B(KEYINPUT57), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n722), .B(KEYINPUT122), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n905), .A2(new_n803), .A3(new_n802), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n903), .B1(new_n921), .B2(new_n922), .ZN(G54));
  AND2_X1   g737(.A1(KEYINPUT58), .A2(G475), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n905), .A2(new_n656), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n656), .B1(new_n905), .B2(new_n924), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n925), .A2(new_n926), .A3(new_n903), .ZN(G60));
  XNOR2_X1  g741(.A(new_n641), .B(KEYINPUT59), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n884), .B2(new_n891), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n637), .A2(new_n638), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n904), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n928), .B1(new_n637), .B2(new_n638), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n917), .A2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT123), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n917), .A2(KEYINPUT123), .A3(new_n932), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(G63));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT60), .Z(new_n939));
  NAND3_X1  g753(.A1(new_n915), .A2(new_n665), .A3(new_n939), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n915), .A2(new_n939), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n535), .A2(new_n536), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n904), .B(new_n940), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT61), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(G66));
  OAI21_X1  g759(.A(G953), .B1(new_n497), .B2(new_n339), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT124), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n870), .A2(new_n874), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n948), .A2(G953), .ZN(new_n949));
  MUX2_X1   g763(.A(new_n947), .B(KEYINPUT124), .S(new_n949), .Z(new_n950));
  INV_X1    g764(.A(new_n907), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(G898), .B2(new_n270), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n950), .B(new_n952), .ZN(G69));
  INV_X1    g767(.A(new_n852), .ZN(new_n954));
  AND4_X1   g768(.A1(new_n775), .A2(new_n818), .A3(new_n782), .A4(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n754), .A2(new_n361), .A3(new_n713), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n810), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT126), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n812), .A2(new_n955), .A3(new_n270), .A4(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(G900), .A2(G953), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n564), .A2(new_n570), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n410), .A2(new_n411), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n962), .B(new_n963), .Z(new_n964));
  NAND2_X1  g778(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(G227), .A2(G900), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(G953), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n715), .A2(new_n954), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT62), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n715), .A2(KEYINPUT62), .A3(new_n954), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n818), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n867), .A2(new_n647), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n974), .A2(new_n692), .A3(new_n621), .A4(new_n771), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n812), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(KEYINPUT125), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT125), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n812), .A2(new_n978), .A3(new_n975), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n973), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n964), .A2(G953), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n965), .B(new_n967), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n961), .A2(G953), .A3(new_n966), .A4(new_n964), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n982), .A2(new_n983), .ZN(G72));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n987), .B1(new_n606), .B2(new_n574), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n903), .B1(new_n883), .B2(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n812), .A2(new_n955), .A3(new_n948), .A4(new_n958), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n990), .A2(KEYINPUT127), .A3(new_n986), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n571), .A2(new_n556), .A3(new_n573), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(KEYINPUT127), .B1(new_n990), .B2(new_n986), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n989), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n556), .B1(new_n571), .B2(new_n573), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n972), .A2(new_n818), .ZN(new_n997));
  INV_X1    g811(.A(new_n979), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n978), .B1(new_n812), .B2(new_n975), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n997), .B(new_n948), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n996), .B1(new_n1000), .B2(new_n986), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n995), .A2(new_n1001), .ZN(G57));
endmodule


