//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT65), .B1(new_n191), .B2(G134), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(new_n189), .A3(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n190), .A2(new_n192), .A3(new_n194), .A4(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n196), .B(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT64), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n199), .A2(KEYINPUT64), .ZN(new_n202));
  OAI21_X1  g016(.A(G143), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n199), .A2(G143), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n203), .A2(KEYINPUT0), .A3(G128), .A4(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n200), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n199), .A2(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XOR2_X1   g026(.A(KEYINPUT0), .B(G128), .Z(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n206), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n198), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT66), .B1(new_n191), .B2(G134), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(new_n189), .A3(G137), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n191), .A2(G134), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G131), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(G131), .B2(new_n196), .ZN(new_n223));
  OR2_X1    g037(.A1(KEYINPUT68), .A2(G128), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT68), .A2(G128), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n209), .B1(new_n200), .B2(new_n208), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n212), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n203), .A2(G128), .A3(new_n205), .A4(new_n228), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n223), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g046(.A(KEYINPUT69), .B(KEYINPUT30), .C1(new_n216), .C2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n196), .A2(G131), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n236));
  NOR2_X1   g050(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT64), .B(G146), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n238), .B1(new_n239), .B2(new_n209), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n240), .A2(new_n226), .B1(new_n211), .B2(new_n210), .ZN(new_n241));
  INV_X1    g055(.A(G128), .ZN(new_n242));
  NOR4_X1   g056(.A1(new_n227), .A2(new_n238), .A3(new_n242), .A4(new_n204), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n235), .B(new_n222), .C1(new_n241), .C2(new_n243), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n196), .A2(G131), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n206), .B(new_n214), .C1(new_n245), .C2(new_n234), .ZN(new_n246));
  OR2_X1    g060(.A1(KEYINPUT69), .A2(KEYINPUT30), .ZN(new_n247));
  NAND2_X1  g061(.A1(KEYINPUT69), .A2(KEYINPUT30), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n244), .A2(new_n246), .A3(new_n247), .A4(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n233), .A2(new_n249), .ZN(new_n250));
  XOR2_X1   g064(.A(G116), .B(G119), .Z(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT2), .B(G113), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n251), .B(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n253), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n244), .A2(new_n255), .A3(new_n246), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n257), .B(G101), .ZN(new_n258));
  NOR2_X1   g072(.A1(G237), .A2(G953), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G210), .ZN(new_n260));
  XOR2_X1   g074(.A(new_n258), .B(new_n260), .Z(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n254), .A2(new_n256), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT28), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n244), .A2(new_n265), .A3(new_n246), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n265), .B1(new_n244), .B2(new_n246), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n264), .B(new_n255), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n253), .B1(new_n216), .B2(new_n232), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(new_n256), .A3(KEYINPUT28), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  AOI22_X1  g085(.A1(KEYINPUT31), .A2(new_n263), .B1(new_n271), .B2(new_n261), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n255), .B1(new_n233), .B2(new_n249), .ZN(new_n273));
  INV_X1    g087(.A(new_n256), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n273), .A2(new_n274), .A3(new_n261), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT31), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT71), .B1(new_n272), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n268), .A2(new_n261), .A3(new_n270), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n279), .B1(new_n275), .B2(new_n276), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n281));
  NOR4_X1   g095(.A1(new_n273), .A2(KEYINPUT31), .A3(new_n274), .A4(new_n261), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n187), .B1(new_n278), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT32), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n271), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT29), .B1(new_n287), .B2(new_n262), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n273), .A2(new_n274), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n288), .B1(new_n289), .B2(new_n262), .ZN(new_n290));
  INV_X1    g104(.A(G902), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n287), .A2(KEYINPUT29), .A3(new_n262), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G472), .ZN(new_n294));
  INV_X1    g108(.A(new_n187), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n281), .B1(new_n280), .B2(new_n282), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n263), .A2(KEYINPUT31), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n297), .A2(new_n277), .A3(KEYINPUT71), .A4(new_n279), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n295), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT32), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n286), .A2(new_n294), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT77), .ZN(new_n302));
  INV_X1    g116(.A(G107), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n303), .A3(G104), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT77), .B1(new_n303), .B2(G104), .ZN(new_n305));
  INV_X1    g119(.A(G104), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(G107), .ZN(new_n307));
  OAI211_X1 g121(.A(G101), .B(new_n304), .C1(new_n305), .C2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT3), .B1(new_n306), .B2(G107), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT3), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(new_n303), .A3(G104), .ZN(new_n311));
  INV_X1    g125(.A(G101), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n306), .A2(G107), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n309), .A2(new_n311), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n308), .A2(new_n314), .A3(KEYINPUT78), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT78), .B1(new_n308), .B2(new_n314), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n230), .A2(new_n231), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT10), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n308), .A2(new_n314), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n242), .B1(new_n211), .B2(KEYINPUT1), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n322), .B1(new_n203), .B2(new_n205), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n321), .B1(new_n243), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT10), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n309), .A2(new_n311), .A3(new_n313), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G101), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(KEYINPUT4), .A3(new_n314), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT4), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n327), .A2(new_n330), .A3(G101), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n329), .A2(new_n206), .A3(new_n214), .A4(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n319), .A2(new_n326), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n198), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n319), .A2(new_n326), .A3(new_n198), .A4(new_n332), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(G110), .B(G140), .ZN(new_n338));
  INV_X1    g152(.A(G953), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n339), .A2(G227), .ZN(new_n340));
  XOR2_X1   g154(.A(new_n338), .B(new_n340), .Z(new_n341));
  OAI211_X1 g155(.A(new_n230), .B(new_n231), .C1(new_n315), .C2(new_n316), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n324), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT12), .B1(new_n343), .B2(new_n334), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT12), .ZN(new_n345));
  AOI211_X1 g159(.A(new_n345), .B(new_n198), .C1(new_n342), .C2(new_n324), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n336), .A2(new_n341), .ZN(new_n348));
  OAI22_X1  g162(.A1(new_n337), .A2(new_n341), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G469), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(new_n291), .ZN(new_n351));
  NAND2_X1  g165(.A1(G469), .A2(G902), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n336), .B1(new_n344), .B2(new_n346), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT79), .ZN(new_n354));
  INV_X1    g168(.A(new_n341), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n356), .B(new_n336), .C1(new_n344), .C2(new_n346), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n348), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n336), .A2(KEYINPUT80), .A3(new_n341), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n335), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n351), .B(new_n352), .C1(new_n363), .C2(new_n350), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT9), .B(G234), .ZN(new_n365));
  OAI21_X1  g179(.A(G221), .B1(new_n365), .B2(G902), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(G214), .B1(G237), .B2(G902), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n215), .A2(G125), .ZN(new_n370));
  INV_X1    g184(.A(G125), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n230), .A2(new_n371), .A3(new_n231), .ZN(new_n372));
  NAND2_X1  g186(.A1(KEYINPUT83), .A2(KEYINPUT7), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n370), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G224), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(G953), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT7), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n374), .B(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n251), .A2(new_n252), .ZN(new_n380));
  INV_X1    g194(.A(G116), .ZN(new_n381));
  NOR3_X1   g195(.A1(new_n381), .A2(KEYINPUT5), .A3(G119), .ZN(new_n382));
  XNOR2_X1  g196(.A(G116), .B(G119), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n382), .B1(new_n383), .B2(KEYINPUT5), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n380), .B1(G113), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT78), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n320), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n308), .A2(new_n314), .A3(KEYINPUT78), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT82), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT82), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n317), .A2(new_n391), .A3(new_n385), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n390), .B(new_n392), .C1(new_n321), .C2(new_n385), .ZN(new_n393));
  XOR2_X1   g207(.A(G110), .B(G122), .Z(new_n394));
  XOR2_X1   g208(.A(new_n394), .B(KEYINPUT8), .Z(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n253), .A2(new_n329), .A3(new_n331), .ZN(new_n397));
  INV_X1    g211(.A(new_n394), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n389), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n379), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n370), .A2(new_n372), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(new_n376), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n398), .B1(new_n389), .B2(new_n397), .ZN(new_n403));
  NAND2_X1  g217(.A1(KEYINPUT81), .A2(KEYINPUT6), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n403), .B1(new_n399), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n389), .A2(new_n397), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n394), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(new_n404), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n402), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n400), .A2(new_n410), .A3(new_n291), .ZN(new_n411));
  OAI21_X1  g225(.A(G210), .B1(G237), .B2(G902), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n399), .A2(new_n405), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n408), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(new_n408), .B2(new_n404), .ZN(new_n417));
  AOI21_X1  g231(.A(G902), .B1(new_n417), .B2(new_n402), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(new_n412), .A3(new_n400), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n369), .B1(new_n414), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n259), .A2(G214), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n209), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n259), .A2(G143), .A3(G214), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT85), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT18), .B1(new_n425), .B2(new_n426), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n427), .B1(new_n428), .B2(new_n197), .ZN(new_n429));
  XNOR2_X1  g243(.A(G125), .B(G140), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n430), .B1(new_n201), .B2(new_n202), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT72), .ZN(new_n432));
  NOR3_X1   g246(.A1(new_n432), .A2(new_n371), .A3(G140), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n433), .B1(new_n432), .B2(new_n430), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n431), .B1(new_n435), .B2(new_n199), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n425), .A2(new_n426), .A3(KEYINPUT18), .A4(G131), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n429), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  OR3_X1    g252(.A1(new_n371), .A2(KEYINPUT16), .A3(G140), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT16), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n439), .B1(new_n434), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n199), .ZN(new_n442));
  OAI211_X1 g256(.A(G146), .B(new_n439), .C1(new_n434), .C2(new_n440), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n425), .A2(G131), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT17), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n423), .A2(new_n197), .A3(new_n424), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n425), .A2(KEYINPUT17), .A3(G131), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n442), .A2(new_n443), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n438), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(G113), .B(G122), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(new_n306), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n438), .A2(new_n449), .A3(new_n452), .ZN(new_n455));
  AOI21_X1  g269(.A(G902), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G475), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n438), .A2(new_n449), .A3(new_n452), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n444), .A2(new_n446), .ZN(new_n460));
  MUX2_X1   g274(.A(new_n430), .B(new_n434), .S(KEYINPUT19), .Z(new_n461));
  OAI211_X1 g275(.A(new_n443), .B(new_n460), .C1(new_n461), .C2(new_n239), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n452), .B1(new_n438), .B2(new_n462), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n457), .B(new_n291), .C1(new_n459), .C2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n438), .A2(new_n462), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n453), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n455), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT20), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n469), .A2(new_n470), .A3(new_n457), .A4(new_n291), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n458), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G952), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(G953), .ZN(new_n474));
  NAND2_X1  g288(.A1(G234), .A2(G237), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  XOR2_X1   g290(.A(KEYINPUT21), .B(G898), .Z(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(G902), .A3(G953), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G217), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n365), .A2(new_n480), .A3(G953), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n209), .B1(new_n224), .B2(new_n225), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT13), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n242), .A2(G143), .ZN(new_n485));
  NOR4_X1   g299(.A1(new_n483), .A2(new_n484), .A3(new_n189), .A4(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n483), .A2(KEYINPUT13), .ZN(new_n488));
  OAI22_X1  g302(.A1(new_n488), .A2(new_n189), .B1(new_n485), .B2(new_n483), .ZN(new_n489));
  XNOR2_X1  g303(.A(G116), .B(G122), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G107), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n303), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n487), .A2(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n381), .A2(KEYINPUT14), .A3(G122), .ZN(new_n495));
  OAI211_X1 g309(.A(G107), .B(new_n495), .C1(new_n491), .C2(KEYINPUT14), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT86), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n490), .A2(KEYINPUT86), .A3(new_n303), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n224), .A2(new_n225), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(G143), .ZN(new_n502));
  INV_X1    g316(.A(new_n485), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(G134), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n189), .B1(new_n483), .B2(new_n485), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n482), .B1(new_n494), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n492), .A2(new_n493), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n502), .A2(new_n484), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n510), .A2(G134), .B1(new_n503), .B2(new_n502), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n509), .B1(new_n511), .B2(new_n486), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n498), .A2(new_n499), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n513), .A2(new_n496), .A3(new_n505), .A4(new_n504), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n512), .A2(new_n514), .A3(new_n481), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n291), .ZN(new_n517));
  INV_X1    g331(.A(G478), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(KEYINPUT15), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n517), .B(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n472), .A2(new_n479), .A3(new_n521), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n367), .A2(new_n421), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n442), .A2(new_n443), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT23), .B1(new_n242), .B2(G119), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n242), .A2(G119), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n527), .B1(new_n501), .B2(G119), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT23), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  XOR2_X1   g344(.A(KEYINPUT24), .B(G110), .Z(new_n531));
  AOI22_X1  g345(.A1(new_n530), .A2(G110), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n524), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT73), .B(G110), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n528), .A2(new_n531), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n443), .B(new_n431), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n339), .A2(G221), .A3(G234), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT22), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(G137), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n541), .B1(new_n533), .B2(new_n537), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n291), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT74), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT25), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n480), .B1(G234), .B2(new_n291), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n546), .A2(KEYINPUT74), .A3(KEYINPUT25), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT75), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n545), .B(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n550), .A2(G902), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT76), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT76), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n552), .A2(new_n559), .A3(new_n556), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n301), .A2(new_n523), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT87), .B(G101), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n562), .B(new_n563), .ZN(G3));
  INV_X1    g378(.A(new_n367), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n291), .B1(new_n278), .B2(new_n283), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n299), .B1(new_n566), .B2(G472), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n561), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n411), .A2(new_n413), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n412), .B1(new_n418), .B2(new_n400), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n368), .B(new_n479), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT88), .B(KEYINPUT33), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n508), .A2(new_n515), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n508), .A2(new_n515), .B1(KEYINPUT88), .B2(KEYINPUT33), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT89), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n577), .A2(new_n578), .A3(G478), .A4(new_n291), .ZN(new_n579));
  NAND2_X1  g393(.A1(KEYINPUT88), .A2(KEYINPUT33), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n516), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n581), .A2(G478), .A3(new_n291), .A4(new_n574), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT89), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n517), .A2(new_n518), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n579), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n466), .A2(new_n471), .ZN(new_n586));
  INV_X1    g400(.A(new_n458), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n572), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n569), .A2(new_n590), .ZN(new_n591));
  XOR2_X1   g405(.A(KEYINPUT34), .B(G104), .Z(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(G6));
  INV_X1    g407(.A(KEYINPUT90), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(new_n464), .B2(new_n465), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n466), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n464), .A2(new_n594), .A3(new_n465), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n458), .A2(KEYINPUT91), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT91), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n599), .B1(new_n456), .B2(new_n457), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n596), .A2(new_n597), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n520), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n602), .A2(new_n572), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n569), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT35), .B(G107), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G9));
  NOR2_X1   g420(.A1(new_n542), .A2(KEYINPUT36), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n538), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n555), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n552), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n523), .A2(new_n567), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT92), .B(KEYINPUT37), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(G110), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n611), .B(new_n613), .ZN(G12));
  INV_X1    g428(.A(new_n610), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n299), .A2(KEYINPUT32), .ZN(new_n616));
  AOI211_X1 g430(.A(new_n285), .B(new_n295), .C1(new_n296), .C2(new_n298), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n615), .B1(new_n618), .B2(new_n294), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n367), .A2(new_n421), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n476), .B(KEYINPUT93), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n622), .B1(G900), .B2(new_n478), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n602), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n619), .A2(KEYINPUT94), .A3(new_n620), .A4(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n301), .A2(new_n620), .A3(new_n610), .A4(new_n625), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT94), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G128), .ZN(G30));
  XOR2_X1   g445(.A(new_n623), .B(KEYINPUT96), .Z(new_n632));
  XOR2_X1   g446(.A(new_n632), .B(KEYINPUT39), .Z(new_n633));
  NAND3_X1  g447(.A1(new_n565), .A2(KEYINPUT97), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT40), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT97), .ZN(new_n636));
  INV_X1    g450(.A(new_n633), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n636), .B1(new_n367), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n634), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n472), .A2(new_n521), .ZN(new_n640));
  AND4_X1   g454(.A1(new_n368), .A2(new_n639), .A3(new_n615), .A4(new_n640), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n634), .A2(new_n638), .ZN(new_n642));
  OR2_X1    g456(.A1(new_n642), .A2(new_n635), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n289), .A2(new_n261), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n269), .A2(new_n256), .A3(new_n261), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n291), .ZN(new_n646));
  OAI21_X1  g460(.A(G472), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n286), .A2(new_n300), .A3(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT95), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n618), .A2(KEYINPUT95), .A3(new_n647), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n414), .A2(new_n419), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT38), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n641), .A2(new_n643), .A3(new_n653), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G143), .ZN(G45));
  NOR2_X1   g471(.A1(new_n589), .A2(new_n624), .ZN(new_n658));
  AND4_X1   g472(.A1(new_n301), .A2(new_n620), .A3(new_n610), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(new_n199), .ZN(G48));
  NAND2_X1  g474(.A1(new_n349), .A2(new_n291), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(G469), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n662), .A2(new_n351), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n366), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n301), .A2(new_n561), .A3(new_n590), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT41), .B(G113), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G15));
  NAND4_X1  g482(.A1(new_n301), .A2(new_n561), .A3(new_n603), .A4(new_n665), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G116), .ZN(G18));
  INV_X1    g484(.A(new_n522), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n664), .A2(new_n421), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n301), .A2(new_n671), .A3(new_n610), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G119), .ZN(G21));
  INV_X1    g488(.A(KEYINPUT98), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n566), .A2(new_n675), .A3(G472), .ZN(new_n676));
  AOI21_X1  g490(.A(G902), .B1(new_n296), .B2(new_n298), .ZN(new_n677));
  INV_X1    g491(.A(G472), .ZN(new_n678));
  OAI21_X1  g492(.A(KEYINPUT98), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n557), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n295), .B1(new_n272), .B2(new_n277), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n676), .A2(new_n679), .A3(new_n680), .A4(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n640), .ZN(new_n684));
  NOR4_X1   g498(.A1(new_n683), .A2(new_n572), .A3(new_n684), .A4(new_n664), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n685), .B(G122), .Z(G24));
  NAND2_X1  g500(.A1(new_n672), .A2(new_n658), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n676), .A2(new_n679), .A3(new_n610), .A4(new_n682), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n371), .ZN(G27));
  OR2_X1    g504(.A1(new_n300), .A2(KEYINPUT100), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n300), .A2(KEYINPUT100), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n691), .A2(new_n286), .A3(new_n294), .A4(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n654), .A2(new_n369), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n658), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n367), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n693), .A2(KEYINPUT42), .A3(new_n680), .A4(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n301), .A2(new_n696), .A3(new_n561), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT99), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n699), .B1(new_n698), .B2(new_n700), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n697), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G131), .ZN(G33));
  AND4_X1   g518(.A1(new_n561), .A2(new_n301), .A3(new_n625), .A4(new_n694), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n565), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G134), .ZN(G36));
  NAND2_X1  g521(.A1(new_n585), .A2(new_n472), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(KEYINPUT43), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  AOI22_X1  g525(.A1(new_n585), .A2(new_n472), .B1(new_n709), .B2(KEYINPUT43), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n711), .B1(new_n712), .B2(new_n710), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n566), .A2(G472), .ZN(new_n714));
  AOI22_X1  g528(.A1(KEYINPUT105), .A2(new_n713), .B1(new_n714), .B2(new_n284), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n711), .B(new_n716), .C1(new_n710), .C2(new_n712), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n715), .A2(KEYINPUT44), .A3(new_n610), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n713), .A2(KEYINPUT105), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n284), .B1(new_n678), .B2(new_n677), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(new_n720), .A3(new_n717), .A4(new_n610), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT103), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n358), .A2(KEYINPUT45), .A3(new_n362), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT101), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n363), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n358), .A2(KEYINPUT101), .A3(KEYINPUT45), .A4(new_n362), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n728), .A2(new_n730), .A3(G469), .A4(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(KEYINPUT46), .A3(new_n352), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT102), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n352), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT46), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT102), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n732), .A2(new_n738), .A3(KEYINPUT46), .A4(new_n352), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n734), .A2(new_n737), .A3(new_n351), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n366), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n725), .B1(new_n741), .B2(new_n637), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n740), .A2(KEYINPUT103), .A3(new_n366), .A4(new_n633), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n724), .A2(new_n742), .A3(new_n694), .A4(new_n743), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT106), .B(G137), .Z(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G39));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(KEYINPUT47), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT107), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n740), .A2(new_n750), .A3(new_n366), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n750), .B1(new_n740), .B2(new_n366), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n749), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n741), .A2(KEYINPUT107), .ZN(new_n754));
  XOR2_X1   g568(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n755));
  NAND3_X1  g569(.A1(new_n740), .A2(new_n750), .A3(new_n366), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n561), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n301), .A2(new_n695), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n758), .A2(KEYINPUT109), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n753), .A2(new_n757), .A3(new_n759), .A4(new_n760), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G140), .ZN(G42));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n659), .A2(new_n689), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n421), .A2(new_n684), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n565), .A2(new_n615), .A3(new_n623), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n648), .B(new_n769), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n630), .A2(new_n768), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT52), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n630), .A2(new_n777), .A3(new_n768), .A4(new_n774), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n479), .ZN(new_n780));
  AOI211_X1 g594(.A(new_n369), .B(new_n780), .C1(new_n414), .C2(new_n419), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n585), .A2(new_n588), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n782), .B1(new_n585), .B2(new_n588), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT111), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n472), .A2(new_n520), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n786), .B1(new_n572), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n787), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n789), .A2(KEYINPUT111), .A3(new_n420), .A4(new_n479), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n785), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n791), .A2(new_n561), .A3(new_n565), .A4(new_n567), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n792), .A2(new_n673), .A3(new_n562), .A4(new_n611), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n666), .A2(new_n669), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n793), .A2(new_n794), .A3(new_n685), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n681), .B1(new_n714), .B2(KEYINPUT98), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(new_n658), .A3(new_n676), .A4(new_n694), .ZN(new_n797));
  INV_X1    g611(.A(new_n654), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n520), .A2(new_n624), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n798), .A2(new_n601), .A3(new_n368), .A4(new_n799), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n800), .A2(KEYINPUT112), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(KEYINPUT112), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n301), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n615), .B1(new_n797), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n565), .B1(new_n804), .B2(new_n705), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n795), .A2(new_n805), .A3(new_n703), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n767), .B1(new_n779), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n775), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n777), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n795), .A2(new_n805), .A3(new_n703), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n775), .A2(new_n808), .A3(KEYINPUT52), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n810), .A2(new_n811), .A3(KEYINPUT53), .A4(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n807), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT115), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n807), .A2(new_n813), .A3(new_n817), .A4(new_n814), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT52), .B1(new_n775), .B2(new_n808), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n806), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT53), .B1(new_n820), .B2(new_n812), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n779), .A2(new_n767), .A3(new_n806), .ZN(new_n822));
  OAI21_X1  g636(.A(KEYINPUT54), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n816), .A2(new_n818), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n709), .A2(KEYINPUT43), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n708), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n710), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n622), .B1(new_n828), .B2(new_n711), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n796), .A2(new_n680), .A3(new_n829), .A4(new_n676), .ZN(new_n830));
  INV_X1    g644(.A(new_n694), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n663), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(new_n366), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n832), .B1(new_n758), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n713), .A2(new_n621), .ZN(new_n836));
  OR4_X1    g650(.A1(new_n664), .A2(new_n688), .A3(new_n831), .A4(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n664), .A2(new_n831), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n759), .A2(new_n476), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n585), .A2(new_n588), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n652), .A2(new_n838), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT50), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n655), .A2(new_n368), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NOR4_X1   g658(.A1(new_n830), .A2(new_n842), .A3(new_n664), .A4(new_n844), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n683), .A2(new_n664), .A3(new_n836), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT50), .B1(new_n846), .B2(new_n843), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n837), .B(new_n841), .C1(new_n845), .C2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n835), .A2(KEYINPUT51), .A3(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n693), .A2(new_n680), .A3(new_n829), .A4(new_n838), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT48), .ZN(new_n852));
  INV_X1    g666(.A(new_n589), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n652), .A2(new_n853), .A3(new_n838), .A4(new_n839), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n850), .A2(new_n474), .A3(new_n852), .A4(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n857));
  INV_X1    g671(.A(new_n832), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n753), .A2(new_n757), .A3(KEYINPUT116), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT116), .B1(new_n753), .B2(new_n757), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n834), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n858), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n848), .A2(KEYINPUT117), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n683), .A2(new_n836), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n865), .A2(new_n665), .A3(new_n843), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n842), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n846), .A2(KEYINPUT50), .A3(new_n843), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n869), .A2(new_n870), .A3(new_n837), .A4(new_n841), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n864), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n856), .B(new_n857), .C1(new_n863), .C2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT116), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n748), .B1(new_n754), .B2(new_n756), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n753), .A2(new_n757), .A3(KEYINPUT116), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n862), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n872), .B1(new_n879), .B2(new_n832), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT118), .B1(new_n880), .B2(KEYINPUT51), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n855), .B1(new_n873), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n865), .A2(new_n672), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n824), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n473), .A2(new_n339), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n653), .A2(new_n655), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT49), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n708), .B1(new_n663), .B2(new_n888), .ZN(new_n889));
  AOI211_X1 g703(.A(new_n369), .B(new_n557), .C1(new_n833), .C2(KEYINPUT49), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n887), .A2(new_n366), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n886), .A2(new_n891), .ZN(G75));
  INV_X1    g706(.A(KEYINPUT56), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n807), .A2(new_n813), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(G902), .ZN(new_n895));
  INV_X1    g709(.A(G210), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT120), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n417), .B(KEYINPUT119), .Z(new_n899));
  XOR2_X1   g713(.A(new_n402), .B(KEYINPUT55), .Z(new_n900));
  XOR2_X1   g714(.A(new_n899), .B(new_n900), .Z(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n339), .A2(G952), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n905), .B1(new_n897), .B2(KEYINPUT120), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n901), .B1(new_n897), .B2(KEYINPUT120), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(G51));
  XOR2_X1   g722(.A(new_n352), .B(KEYINPUT57), .Z(new_n909));
  INV_X1    g723(.A(new_n815), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n814), .B1(new_n807), .B2(new_n813), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n349), .B(KEYINPUT121), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n895), .A2(new_n732), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n904), .B1(new_n914), .B2(new_n915), .ZN(G54));
  NAND4_X1  g730(.A1(new_n894), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n917));
  INV_X1    g731(.A(new_n469), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n919), .A2(new_n920), .A3(new_n904), .ZN(G60));
  NAND3_X1  g735(.A1(new_n816), .A2(new_n823), .A3(new_n818), .ZN(new_n922));
  NAND2_X1  g736(.A1(G478), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT59), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n577), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n577), .B(new_n924), .C1(new_n910), .C2(new_n911), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n925), .A2(new_n927), .A3(new_n904), .ZN(G63));
  NAND2_X1  g742(.A1(G217), .A2(G902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT60), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n807), .B2(new_n813), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n904), .B1(new_n931), .B2(new_n608), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n554), .B2(new_n931), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(G66));
  INV_X1    g749(.A(new_n477), .ZN(new_n936));
  OAI21_X1  g750(.A(G953), .B1(new_n936), .B2(new_n375), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n795), .B2(G953), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT122), .ZN(new_n939));
  INV_X1    g753(.A(new_n899), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(G898), .B2(new_n339), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n939), .B(new_n941), .ZN(G69));
  OR2_X1    g756(.A1(new_n339), .A2(G900), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n718), .A2(new_n723), .A3(new_n694), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n693), .A2(new_n680), .A3(new_n769), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n946), .A2(new_n742), .A3(new_n743), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n630), .A2(new_n768), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n947), .A2(new_n703), .A3(new_n706), .A4(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n761), .B2(new_n764), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n943), .B1(new_n950), .B2(G953), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(KEYINPUT124), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n250), .B(new_n461), .Z(new_n953));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n954), .B(new_n943), .C1(new_n950), .C2(G953), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n339), .B1(G227), .B2(G900), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n957), .A2(KEYINPUT125), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n301), .A2(new_n561), .ZN(new_n959));
  OR3_X1    g773(.A1(new_n783), .A2(new_n784), .A3(new_n789), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n959), .A2(new_n642), .A3(new_n694), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n744), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(KEYINPUT123), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT123), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n744), .A2(new_n964), .A3(new_n961), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n948), .A2(new_n656), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT62), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n948), .A2(new_n656), .A3(KEYINPUT62), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n765), .A2(new_n966), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n339), .ZN(new_n973));
  INV_X1    g787(.A(new_n953), .ZN(new_n974));
  AOI22_X1  g788(.A1(new_n973), .A2(new_n974), .B1(KEYINPUT125), .B2(new_n957), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n956), .A2(new_n958), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n958), .B1(new_n956), .B2(new_n975), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(G72));
  INV_X1    g792(.A(new_n644), .ZN(new_n979));
  NAND2_X1  g793(.A1(G472), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT63), .Z(new_n981));
  NAND2_X1  g795(.A1(new_n289), .A2(new_n261), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n979), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT127), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n821), .B2(new_n822), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n981), .B(KEYINPUT126), .Z(new_n986));
  AOI21_X1  g800(.A(new_n986), .B1(new_n950), .B2(new_n795), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n905), .B(new_n985), .C1(new_n987), .C2(new_n982), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n765), .A2(new_n966), .A3(new_n795), .A4(new_n971), .ZN(new_n989));
  INV_X1    g803(.A(new_n986), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n979), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n988), .A2(new_n991), .ZN(G57));
endmodule


