

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765;

  XNOR2_X1 U372 ( .A(KEYINPUT105), .B(n576), .ZN(n658) );
  NOR2_X1 U373 ( .A1(n589), .A2(n579), .ZN(n696) );
  BUF_X1 U374 ( .A(G107), .Z(n349) );
  XNOR2_X1 U375 ( .A(n737), .B(n369), .ZN(n368) );
  XNOR2_X1 U376 ( .A(n471), .B(n467), .ZN(n737) );
  NAND2_X2 U377 ( .A1(n455), .A2(n350), .ZN(n466) );
  NOR2_X1 U378 ( .A1(G953), .A2(G237), .ZN(n530) );
  NOR2_X1 U379 ( .A1(n579), .A2(n620), .ZN(n445) );
  INV_X1 U380 ( .A(G953), .ZN(n755) );
  AND2_X2 U381 ( .A1(n477), .A2(n351), .ZN(n455) );
  XNOR2_X2 U382 ( .A(n588), .B(KEYINPUT80), .ZN(n477) );
  AND2_X2 U383 ( .A1(n405), .A2(KEYINPUT19), .ZN(n404) );
  XNOR2_X2 U384 ( .A(n368), .B(n367), .ZN(n717) );
  INV_X2 U385 ( .A(n672), .ZN(n350) );
  INV_X1 U386 ( .A(n668), .ZN(n351) );
  XNOR2_X1 U387 ( .A(n753), .B(n476), .ZN(n388) );
  INV_X1 U388 ( .A(G113), .ZN(n470) );
  INV_X1 U389 ( .A(KEYINPUT45), .ZN(n411) );
  AND2_X1 U390 ( .A1(n391), .A2(n389), .ZN(n641) );
  AND2_X1 U391 ( .A1(n394), .A2(n392), .ZN(n391) );
  AND2_X1 U392 ( .A1(n431), .A2(n746), .ZN(n672) );
  XNOR2_X1 U393 ( .A(n634), .B(KEYINPUT82), .ZN(n668) );
  NOR2_X1 U394 ( .A1(n374), .A2(n373), .ZN(n372) );
  AND2_X1 U395 ( .A1(n371), .A2(n376), .ZN(n370) );
  NAND2_X1 U396 ( .A1(n375), .A2(n377), .ZN(n373) );
  AND2_X1 U397 ( .A1(n587), .A2(n432), .ZN(n375) );
  XNOR2_X1 U398 ( .A(n387), .B(n571), .ZN(n763) );
  XOR2_X1 U399 ( .A(n632), .B(KEYINPUT38), .Z(n673) );
  INV_X1 U400 ( .A(n507), .ZN(n467) );
  XNOR2_X1 U401 ( .A(n469), .B(n468), .ZN(n507) );
  XNOR2_X1 U402 ( .A(n541), .B(n472), .ZN(n471) );
  XNOR2_X1 U403 ( .A(n470), .B(G119), .ZN(n469) );
  XNOR2_X1 U404 ( .A(KEYINPUT3), .B(KEYINPUT69), .ZN(n468) );
  XNOR2_X1 U405 ( .A(KEYINPUT72), .B(KEYINPUT16), .ZN(n472) );
  XNOR2_X2 U406 ( .A(n508), .B(n493), .ZN(n753) );
  NAND2_X1 U407 ( .A1(n395), .A2(n356), .ZN(n634) );
  XNOR2_X1 U408 ( .A(n396), .B(n415), .ZN(n395) );
  INV_X1 U409 ( .A(n666), .ZN(n414) );
  XOR2_X1 U410 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n527) );
  XNOR2_X1 U411 ( .A(KEYINPUT12), .B(KEYINPUT99), .ZN(n526) );
  XOR2_X1 U412 ( .A(KEYINPUT95), .B(KEYINPUT11), .Z(n525) );
  AND2_X1 U413 ( .A1(n441), .A2(n679), .ZN(n605) );
  AND2_X1 U414 ( .A1(n452), .A2(n361), .ZN(n441) );
  NOR2_X1 U415 ( .A1(n765), .A2(n762), .ZN(n440) );
  XOR2_X1 U416 ( .A(G101), .B(KEYINPUT66), .Z(n499) );
  NOR2_X2 U417 ( .A1(n408), .A2(n517), .ZN(n403) );
  XNOR2_X1 U418 ( .A(KEYINPUT15), .B(G902), .ZN(n636) );
  XNOR2_X1 U419 ( .A(n492), .B(G131), .ZN(n493) );
  XNOR2_X1 U420 ( .A(n499), .B(n739), .ZN(n511) );
  XNOR2_X1 U421 ( .A(n450), .B(n349), .ZN(n449) );
  XNOR2_X1 U422 ( .A(G140), .B(KEYINPUT75), .ZN(n450) );
  INV_X1 U423 ( .A(G146), .ZN(n476) );
  NAND2_X1 U424 ( .A1(n572), .A2(n378), .ZN(n371) );
  NOR2_X1 U425 ( .A1(n763), .A2(KEYINPUT44), .ZN(n572) );
  INV_X1 U426 ( .A(KEYINPUT1), .ZN(n487) );
  XNOR2_X1 U427 ( .A(n568), .B(KEYINPUT67), .ZN(n690) );
  XNOR2_X1 U428 ( .A(n688), .B(KEYINPUT6), .ZN(n620) );
  XNOR2_X1 U429 ( .A(n543), .B(n542), .ZN(n551) );
  INV_X1 U430 ( .A(KEYINPUT8), .ZN(n542) );
  NAND2_X1 U431 ( .A1(n755), .A2(G234), .ZN(n543) );
  NAND2_X1 U432 ( .A1(n350), .A2(n639), .ZN(n485) );
  XNOR2_X1 U433 ( .A(n461), .B(n537), .ZN(n539) );
  XNOR2_X1 U434 ( .A(n462), .B(KEYINPUT9), .ZN(n461) );
  XNOR2_X1 U435 ( .A(KEYINPUT100), .B(KEYINPUT102), .ZN(n462) );
  BUF_X1 U436 ( .A(n601), .Z(n417) );
  XNOR2_X1 U437 ( .A(n453), .B(KEYINPUT41), .ZN(n707) );
  AND2_X1 U438 ( .A1(n680), .A2(n617), .ZN(n453) );
  NOR2_X1 U439 ( .A1(n607), .A2(n673), .ZN(n597) );
  NAND2_X1 U440 ( .A1(n379), .A2(n385), .ZN(n381) );
  NOR2_X1 U441 ( .A1(n583), .A2(KEYINPUT34), .ZN(n385) );
  AND2_X1 U442 ( .A1(n380), .A2(n383), .ZN(n382) );
  AND2_X1 U443 ( .A1(n386), .A2(n384), .ZN(n383) );
  INV_X1 U444 ( .A(n357), .ZN(n384) );
  NOR2_X1 U445 ( .A1(n677), .A2(n548), .ZN(n549) );
  NAND2_X1 U446 ( .A1(n399), .A2(n397), .ZN(n607) );
  XNOR2_X1 U447 ( .A(n416), .B(n398), .ZN(n397) );
  NOR2_X1 U448 ( .A1(n590), .A2(n355), .ZN(n399) );
  INV_X1 U449 ( .A(KEYINPUT30), .ZN(n398) );
  XNOR2_X1 U450 ( .A(n600), .B(KEYINPUT28), .ZN(n452) );
  NOR2_X1 U451 ( .A1(n589), .A2(n619), .ZN(n600) );
  XNOR2_X1 U452 ( .A(n465), .B(n463), .ZN(n577) );
  XNOR2_X1 U453 ( .A(n464), .B(G478), .ZN(n463) );
  OR2_X1 U454 ( .A1(n727), .A2(G902), .ZN(n465) );
  INV_X1 U455 ( .A(KEYINPUT104), .ZN(n464) );
  OR2_X1 U456 ( .A1(n635), .A2(n478), .ZN(n394) );
  AND2_X1 U457 ( .A1(n482), .A2(n393), .ZN(n392) );
  NOR2_X1 U458 ( .A1(n363), .A2(n736), .ZN(n393) );
  AND2_X1 U459 ( .A1(n485), .A2(n640), .ZN(n390) );
  INV_X1 U460 ( .A(KEYINPUT47), .ZN(n442) );
  OR2_X1 U461 ( .A1(G237), .A2(G902), .ZN(n515) );
  XOR2_X1 U462 ( .A(G116), .B(KEYINPUT74), .Z(n495) );
  NOR2_X1 U463 ( .A1(n674), .A2(KEYINPUT19), .ZN(n401) );
  XNOR2_X1 U464 ( .A(G113), .B(G131), .ZN(n521) );
  XOR2_X1 U465 ( .A(G122), .B(G143), .Z(n522) );
  XNOR2_X1 U466 ( .A(G104), .B(KEYINPUT98), .ZN(n524) );
  XNOR2_X1 U467 ( .A(n511), .B(n512), .ZN(n369) );
  XNOR2_X1 U468 ( .A(KEYINPUT17), .B(KEYINPUT76), .ZN(n512) );
  INV_X1 U469 ( .A(KEYINPUT4), .ZN(n491) );
  AND2_X1 U470 ( .A1(n628), .A2(n438), .ZN(n437) );
  AND2_X1 U471 ( .A1(n611), .A2(n610), .ZN(n438) );
  INV_X1 U472 ( .A(KEYINPUT48), .ZN(n415) );
  OR2_X2 U473 ( .A1(n717), .A2(n358), .ZN(n407) );
  NAND2_X1 U474 ( .A1(n352), .A2(n513), .ZN(n409) );
  NAND2_X1 U475 ( .A1(n569), .A2(n577), .ZN(n677) );
  OR2_X2 U476 ( .A1(n629), .A2(n446), .ZN(n579) );
  XNOR2_X1 U477 ( .A(n559), .B(n458), .ZN(n685) );
  XNOR2_X1 U478 ( .A(n561), .B(n558), .ZN(n458) );
  NOR2_X1 U479 ( .A1(G902), .A2(n731), .ZN(n559) );
  INV_X1 U480 ( .A(n483), .ZN(n479) );
  NOR2_X1 U481 ( .A1(n483), .A2(n481), .ZN(n480) );
  INV_X1 U482 ( .A(n639), .ZN(n481) );
  XNOR2_X1 U483 ( .A(G140), .B(KEYINPUT10), .ZN(n519) );
  XNOR2_X1 U484 ( .A(n511), .B(n448), .ZN(n447) );
  XNOR2_X1 U485 ( .A(n500), .B(n449), .ZN(n448) );
  XNOR2_X1 U486 ( .A(n629), .B(n486), .ZN(n626) );
  INV_X1 U487 ( .A(KEYINPUT88), .ZN(n486) );
  NOR2_X1 U488 ( .A1(n603), .A2(n444), .ZN(n443) );
  INV_X1 U489 ( .A(n417), .ZN(n444) );
  OR2_X1 U490 ( .A1(n562), .A2(G902), .ZN(n435) );
  AND2_X1 U491 ( .A1(n690), .A2(n601), .ZN(n582) );
  INV_X1 U492 ( .A(KEYINPUT0), .ZN(n474) );
  XNOR2_X1 U493 ( .A(n536), .B(n535), .ZN(n578) );
  BUF_X1 U494 ( .A(n685), .Z(n420) );
  XNOR2_X1 U495 ( .A(G110), .B(G104), .ZN(n739) );
  XNOR2_X1 U496 ( .A(G134), .B(KEYINPUT103), .ZN(n538) );
  NOR2_X1 U497 ( .A1(n634), .A2(n638), .ZN(n431) );
  XNOR2_X1 U498 ( .A(n451), .B(n413), .ZN(n762) );
  XNOR2_X1 U499 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n413) );
  XNOR2_X1 U500 ( .A(n616), .B(n615), .ZN(n765) );
  NAND2_X1 U501 ( .A1(n382), .A2(n381), .ZN(n387) );
  AND2_X1 U502 ( .A1(n452), .A2(n443), .ZN(n656) );
  INV_X1 U503 ( .A(KEYINPUT60), .ZN(n425) );
  INV_X1 U504 ( .A(KEYINPUT122), .ZN(n423) );
  INV_X1 U505 ( .A(KEYINPUT56), .ZN(n421) );
  XOR2_X1 U506 ( .A(n514), .B(KEYINPUT79), .Z(n352) );
  XNOR2_X1 U507 ( .A(G472), .B(KEYINPUT94), .ZN(n353) );
  XOR2_X1 U508 ( .A(G110), .B(G137), .Z(n354) );
  INV_X1 U509 ( .A(n688), .ZN(n589) );
  XNOR2_X1 U510 ( .A(n445), .B(KEYINPUT33), .ZN(n708) );
  AND2_X1 U511 ( .A1(n595), .A2(n594), .ZN(n355) );
  AND2_X1 U512 ( .A1(n414), .A2(n667), .ZN(n356) );
  OR2_X1 U513 ( .A1(n569), .A2(n577), .ZN(n357) );
  OR2_X1 U514 ( .A1(n352), .A2(n513), .ZN(n358) );
  AND2_X1 U515 ( .A1(G217), .A2(n551), .ZN(n359) );
  AND2_X1 U516 ( .A1(n407), .A2(n401), .ZN(n360) );
  AND2_X1 U517 ( .A1(n443), .A2(n442), .ZN(n361) );
  XNOR2_X1 U518 ( .A(n516), .B(KEYINPUT89), .ZN(n674) );
  XNOR2_X1 U519 ( .A(KEYINPUT71), .B(KEYINPUT22), .ZN(n362) );
  AND2_X1 U520 ( .A1(n640), .A2(n484), .ZN(n363) );
  XNOR2_X1 U521 ( .A(n723), .B(n722), .ZN(n364) );
  XNOR2_X1 U522 ( .A(n719), .B(n718), .ZN(n365) );
  INV_X1 U523 ( .A(KEYINPUT19), .ZN(n517) );
  OR2_X1 U524 ( .A1(n640), .A2(n484), .ZN(n483) );
  INV_X1 U525 ( .A(n736), .ZN(n429) );
  XOR2_X1 U526 ( .A(n725), .B(n489), .Z(n366) );
  XNOR2_X1 U527 ( .A(n456), .B(n508), .ZN(n367) );
  XNOR2_X2 U528 ( .A(n565), .B(KEYINPUT85), .ZN(n378) );
  NAND2_X1 U529 ( .A1(n372), .A2(n370), .ZN(n412) );
  NOR2_X1 U530 ( .A1(n378), .A2(n433), .ZN(n374) );
  NAND2_X1 U531 ( .A1(n378), .A2(n567), .ZN(n376) );
  NAND2_X1 U532 ( .A1(n763), .A2(KEYINPUT44), .ZN(n377) );
  INV_X1 U533 ( .A(n708), .ZN(n379) );
  NAND2_X1 U534 ( .A1(n708), .A2(KEYINPUT34), .ZN(n380) );
  NAND2_X1 U535 ( .A1(n583), .A2(KEYINPUT34), .ZN(n386) );
  XNOR2_X1 U536 ( .A(n388), .B(n436), .ZN(n562) );
  XNOR2_X1 U537 ( .A(n388), .B(n447), .ZN(n721) );
  NAND2_X1 U538 ( .A1(n390), .A2(n466), .ZN(n389) );
  NAND2_X1 U539 ( .A1(n439), .A2(n437), .ZN(n396) );
  NAND2_X1 U540 ( .A1(n408), .A2(n407), .ZN(n632) );
  NAND2_X1 U541 ( .A1(n402), .A2(n400), .ZN(n602) );
  NAND2_X1 U542 ( .A1(n408), .A2(n360), .ZN(n400) );
  NOR2_X2 U543 ( .A1(n404), .A2(n403), .ZN(n402) );
  NAND2_X1 U544 ( .A1(n407), .A2(n406), .ZN(n405) );
  INV_X1 U545 ( .A(n674), .ZN(n406) );
  AND2_X2 U546 ( .A1(n410), .A2(n409), .ZN(n408) );
  NAND2_X1 U547 ( .A1(n717), .A2(n352), .ZN(n410) );
  XNOR2_X2 U548 ( .A(n412), .B(n411), .ZN(n669) );
  NOR2_X2 U549 ( .A1(n669), .A2(n636), .ZN(n588) );
  NAND2_X1 U550 ( .A1(n688), .A2(n406), .ZN(n416) );
  XNOR2_X1 U551 ( .A(n418), .B(n555), .ZN(n556) );
  XNOR2_X1 U552 ( .A(n554), .B(n553), .ZN(n418) );
  XNOR2_X1 U553 ( .A(n359), .B(n419), .ZN(n544) );
  XNOR2_X1 U554 ( .A(n541), .B(n540), .ZN(n419) );
  XNOR2_X1 U555 ( .A(n422), .B(n421), .ZN(G51) );
  NAND2_X1 U556 ( .A1(n428), .A2(n429), .ZN(n422) );
  XNOR2_X1 U557 ( .A(n424), .B(n423), .ZN(G54) );
  NAND2_X1 U558 ( .A1(n427), .A2(n429), .ZN(n424) );
  XNOR2_X1 U559 ( .A(n426), .B(n425), .ZN(G60) );
  NAND2_X1 U560 ( .A1(n430), .A2(n429), .ZN(n426) );
  XNOR2_X1 U561 ( .A(n724), .B(n364), .ZN(n427) );
  XNOR2_X1 U562 ( .A(n720), .B(n365), .ZN(n428) );
  XNOR2_X1 U563 ( .A(n726), .B(n366), .ZN(n430) );
  NAND2_X2 U564 ( .A1(n466), .A2(n485), .ZN(n732) );
  NAND2_X1 U565 ( .A1(n567), .A2(n566), .ZN(n432) );
  NAND2_X1 U566 ( .A1(KEYINPUT44), .A2(KEYINPUT64), .ZN(n433) );
  NAND2_X2 U567 ( .A1(n434), .A2(n460), .ZN(n459) );
  XNOR2_X2 U568 ( .A(n550), .B(n362), .ZN(n434) );
  AND2_X1 U569 ( .A1(n434), .A2(n454), .ZN(n573) );
  XNOR2_X2 U570 ( .A(n435), .B(n353), .ZN(n688) );
  XNOR2_X1 U571 ( .A(n498), .B(n499), .ZN(n436) );
  XNOR2_X1 U572 ( .A(n440), .B(KEYINPUT46), .ZN(n439) );
  NAND2_X1 U573 ( .A1(n679), .A2(n656), .ZN(n606) );
  NAND2_X1 U574 ( .A1(n452), .A2(n417), .ZN(n618) );
  INV_X1 U575 ( .A(n629), .ZN(n691) );
  INV_X1 U576 ( .A(n690), .ZN(n446) );
  NOR2_X1 U577 ( .A1(n707), .A2(n618), .ZN(n451) );
  INV_X1 U578 ( .A(n691), .ZN(n454) );
  NAND2_X1 U579 ( .A1(n350), .A2(n351), .ZN(n635) );
  XNOR2_X1 U580 ( .A(n510), .B(n520), .ZN(n456) );
  OR2_X2 U581 ( .A1(n721), .A2(G902), .ZN(n488) );
  NOR2_X1 U582 ( .A1(n613), .A2(n612), .ZN(n616) );
  XNOR2_X1 U583 ( .A(n556), .B(n457), .ZN(n731) );
  INV_X1 U584 ( .A(n752), .ZN(n457) );
  NAND2_X1 U585 ( .A1(n764), .A2(n651), .ZN(n565) );
  XNOR2_X2 U586 ( .A(n459), .B(KEYINPUT32), .ZN(n764) );
  AND2_X1 U587 ( .A1(n564), .A2(n626), .ZN(n460) );
  XNOR2_X2 U588 ( .A(n473), .B(G122), .ZN(n541) );
  XNOR2_X2 U589 ( .A(G116), .B(G107), .ZN(n473) );
  XNOR2_X2 U590 ( .A(n475), .B(n474), .ZN(n580) );
  NAND2_X1 U591 ( .A1(n602), .A2(n518), .ZN(n475) );
  XNOR2_X2 U592 ( .A(n540), .B(n491), .ZN(n508) );
  NAND2_X1 U593 ( .A1(n350), .A2(n480), .ZN(n482) );
  NAND2_X1 U594 ( .A1(n477), .A2(n479), .ZN(n478) );
  INV_X1 U595 ( .A(G472), .ZN(n484) );
  XNOR2_X2 U596 ( .A(n601), .B(n487), .ZN(n629) );
  XNOR2_X2 U597 ( .A(n488), .B(n501), .ZN(n601) );
  XNOR2_X2 U598 ( .A(G128), .B(KEYINPUT78), .ZN(n490) );
  INV_X1 U599 ( .A(n669), .ZN(n746) );
  XNOR2_X1 U600 ( .A(KEYINPUT59), .B(KEYINPUT65), .ZN(n489) );
  XNOR2_X1 U601 ( .A(n509), .B(KEYINPUT18), .ZN(n510) );
  INV_X1 U602 ( .A(n684), .ZN(n548) );
  XNOR2_X1 U603 ( .A(n497), .B(n507), .ZN(n498) );
  XNOR2_X1 U604 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U605 ( .A(n557), .B(KEYINPUT91), .ZN(n558) );
  XNOR2_X1 U606 ( .A(KEYINPUT13), .B(G475), .ZN(n535) );
  XNOR2_X1 U607 ( .A(n614), .B(KEYINPUT107), .ZN(n615) );
  NOR2_X1 U608 ( .A1(G952), .A2(n755), .ZN(n736) );
  XNOR2_X2 U609 ( .A(n490), .B(G143), .ZN(n540) );
  XOR2_X1 U610 ( .A(G137), .B(G134), .Z(n492) );
  NAND2_X1 U611 ( .A1(n530), .A2(G210), .ZN(n494) );
  XNOR2_X1 U612 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U613 ( .A(n496), .B(KEYINPUT5), .Z(n497) );
  XNOR2_X1 U614 ( .A(n562), .B(KEYINPUT62), .ZN(n640) );
  XNOR2_X1 U615 ( .A(KEYINPUT68), .B(G469), .ZN(n501) );
  NAND2_X1 U616 ( .A1(G227), .A2(n755), .ZN(n500) );
  NOR2_X1 U617 ( .A1(G898), .A2(n755), .ZN(n741) );
  NAND2_X1 U618 ( .A1(G234), .A2(G237), .ZN(n502) );
  XNOR2_X1 U619 ( .A(n502), .B(KEYINPUT14), .ZN(n504) );
  NAND2_X1 U620 ( .A1(G902), .A2(n504), .ZN(n591) );
  INV_X1 U621 ( .A(n591), .ZN(n503) );
  NAND2_X1 U622 ( .A1(n741), .A2(n503), .ZN(n506) );
  NAND2_X1 U623 ( .A1(G952), .A2(n504), .ZN(n706) );
  NOR2_X1 U624 ( .A1(G953), .A2(n706), .ZN(n505) );
  XOR2_X1 U625 ( .A(KEYINPUT90), .B(n505), .Z(n594) );
  NAND2_X1 U626 ( .A1(n506), .A2(n594), .ZN(n518) );
  AND2_X1 U627 ( .A1(G224), .A2(n755), .ZN(n509) );
  XNOR2_X1 U628 ( .A(G146), .B(G125), .ZN(n520) );
  INV_X1 U629 ( .A(n636), .ZN(n513) );
  NAND2_X1 U630 ( .A1(G210), .A2(n515), .ZN(n514) );
  NAND2_X1 U631 ( .A1(n515), .A2(G214), .ZN(n516) );
  XOR2_X1 U632 ( .A(n520), .B(n519), .Z(n752) );
  XNOR2_X1 U633 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U634 ( .A(n752), .B(n523), .Z(n534) );
  XNOR2_X1 U635 ( .A(n525), .B(n524), .ZN(n529) );
  XNOR2_X1 U636 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U637 ( .A(n529), .B(n528), .Z(n532) );
  NAND2_X1 U638 ( .A1(G214), .A2(n530), .ZN(n531) );
  XNOR2_X1 U639 ( .A(n534), .B(n533), .ZN(n725) );
  NOR2_X1 U640 ( .A1(G902), .A2(n725), .ZN(n536) );
  INV_X1 U641 ( .A(n578), .ZN(n569) );
  XNOR2_X1 U642 ( .A(KEYINPUT7), .B(KEYINPUT101), .ZN(n537) );
  XNOR2_X1 U643 ( .A(n539), .B(n538), .ZN(n545) );
  XOR2_X1 U644 ( .A(n545), .B(n544), .Z(n727) );
  NAND2_X1 U645 ( .A1(G234), .A2(n636), .ZN(n546) );
  XNOR2_X1 U646 ( .A(KEYINPUT20), .B(n546), .ZN(n560) );
  NAND2_X1 U647 ( .A1(G221), .A2(n560), .ZN(n547) );
  XOR2_X1 U648 ( .A(KEYINPUT21), .B(n547), .Z(n684) );
  NAND2_X1 U649 ( .A1(n580), .A2(n549), .ZN(n550) );
  NAND2_X1 U650 ( .A1(G221), .A2(n551), .ZN(n555) );
  XNOR2_X1 U651 ( .A(G119), .B(G128), .ZN(n552) );
  XNOR2_X1 U652 ( .A(n354), .B(n552), .ZN(n554) );
  XOR2_X1 U653 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n553) );
  XNOR2_X1 U654 ( .A(KEYINPUT25), .B(KEYINPUT92), .ZN(n557) );
  AND2_X1 U655 ( .A1(n560), .A2(G217), .ZN(n561) );
  NOR2_X1 U656 ( .A1(n420), .A2(n688), .ZN(n563) );
  NAND2_X1 U657 ( .A1(n573), .A2(n563), .ZN(n651) );
  INV_X1 U658 ( .A(n620), .ZN(n575) );
  NOR2_X1 U659 ( .A1(n575), .A2(n420), .ZN(n564) );
  INV_X1 U660 ( .A(KEYINPUT44), .ZN(n566) );
  INV_X1 U661 ( .A(KEYINPUT64), .ZN(n567) );
  INV_X1 U662 ( .A(n580), .ZN(n583) );
  NAND2_X1 U663 ( .A1(n684), .A2(n685), .ZN(n568) );
  XNOR2_X1 U664 ( .A(KEYINPUT77), .B(KEYINPUT35), .ZN(n570) );
  XNOR2_X1 U665 ( .A(n570), .B(KEYINPUT83), .ZN(n571) );
  NAND2_X1 U666 ( .A1(n420), .A2(n573), .ZN(n574) );
  NOR2_X1 U667 ( .A1(n575), .A2(n574), .ZN(n642) );
  NAND2_X1 U668 ( .A1(n578), .A2(n577), .ZN(n576) );
  NOR2_X1 U669 ( .A1(n578), .A2(n577), .ZN(n661) );
  NOR2_X1 U670 ( .A1(n658), .A2(n661), .ZN(n604) );
  NAND2_X1 U671 ( .A1(n696), .A2(n580), .ZN(n581) );
  XNOR2_X1 U672 ( .A(KEYINPUT31), .B(n581), .ZN(n662) );
  XNOR2_X1 U673 ( .A(n582), .B(KEYINPUT93), .ZN(n590) );
  NAND2_X1 U674 ( .A1(n589), .A2(n580), .ZN(n584) );
  NOR2_X1 U675 ( .A1(n590), .A2(n584), .ZN(n646) );
  NOR2_X1 U676 ( .A1(n662), .A2(n646), .ZN(n585) );
  NOR2_X1 U677 ( .A1(n604), .A2(n585), .ZN(n586) );
  NOR2_X1 U678 ( .A1(n642), .A2(n586), .ZN(n587) );
  NOR2_X1 U679 ( .A1(G900), .A2(n591), .ZN(n592) );
  NAND2_X1 U680 ( .A1(G953), .A2(n592), .ZN(n593) );
  XNOR2_X1 U681 ( .A(KEYINPUT106), .B(n593), .ZN(n595) );
  XNOR2_X1 U682 ( .A(KEYINPUT70), .B(KEYINPUT39), .ZN(n596) );
  XNOR2_X1 U683 ( .A(n597), .B(n596), .ZN(n613) );
  INV_X1 U684 ( .A(n661), .ZN(n598) );
  NOR2_X1 U685 ( .A1(n613), .A2(n598), .ZN(n666) );
  NOR2_X1 U686 ( .A1(n420), .A2(n355), .ZN(n599) );
  NAND2_X1 U687 ( .A1(n599), .A2(n684), .ZN(n619) );
  INV_X1 U688 ( .A(n602), .ZN(n603) );
  INV_X1 U689 ( .A(n604), .ZN(n679) );
  XNOR2_X1 U690 ( .A(n605), .B(KEYINPUT73), .ZN(n611) );
  NAND2_X1 U691 ( .A1(n606), .A2(KEYINPUT47), .ZN(n609) );
  INV_X1 U692 ( .A(n632), .ZN(n623) );
  NOR2_X1 U693 ( .A1(n607), .A2(n357), .ZN(n608) );
  NAND2_X1 U694 ( .A1(n623), .A2(n608), .ZN(n655) );
  AND2_X1 U695 ( .A1(n609), .A2(n655), .ZN(n610) );
  INV_X1 U696 ( .A(n658), .ZN(n612) );
  INV_X1 U697 ( .A(KEYINPUT40), .ZN(n614) );
  NOR2_X1 U698 ( .A1(n674), .A2(n673), .ZN(n680) );
  INV_X1 U699 ( .A(n677), .ZN(n617) );
  XOR2_X1 U700 ( .A(KEYINPUT36), .B(KEYINPUT86), .Z(n625) );
  NOR2_X1 U701 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U702 ( .A1(n658), .A2(n621), .ZN(n622) );
  NOR2_X1 U703 ( .A1(n674), .A2(n622), .ZN(n630) );
  NAND2_X1 U704 ( .A1(n630), .A2(n623), .ZN(n624) );
  XNOR2_X1 U705 ( .A(n625), .B(n624), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n665) );
  XNOR2_X1 U707 ( .A(KEYINPUT84), .B(n665), .ZN(n628) );
  NAND2_X1 U708 ( .A1(n630), .A2(n454), .ZN(n631) );
  XNOR2_X1 U709 ( .A(n631), .B(KEYINPUT43), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n667) );
  INV_X1 U711 ( .A(KEYINPUT2), .ZN(n638) );
  XOR2_X1 U712 ( .A(KEYINPUT81), .B(n636), .Z(n637) );
  NOR2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U714 ( .A(KEYINPUT63), .B(n641), .Z(G57) );
  XNOR2_X1 U715 ( .A(G101), .B(n642), .ZN(n643) );
  XNOR2_X1 U716 ( .A(n643), .B(KEYINPUT109), .ZN(G3) );
  NAND2_X1 U717 ( .A1(n646), .A2(n658), .ZN(n644) );
  XNOR2_X1 U718 ( .A(n644), .B(KEYINPUT110), .ZN(n645) );
  XNOR2_X1 U719 ( .A(G104), .B(n645), .ZN(G6) );
  XOR2_X1 U720 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n648) );
  NAND2_X1 U721 ( .A1(n646), .A2(n661), .ZN(n647) );
  XNOR2_X1 U722 ( .A(n648), .B(n647), .ZN(n650) );
  XOR2_X1 U723 ( .A(n349), .B(KEYINPUT111), .Z(n649) );
  XNOR2_X1 U724 ( .A(n650), .B(n649), .ZN(G9) );
  XNOR2_X1 U725 ( .A(n651), .B(G110), .ZN(G12) );
  XOR2_X1 U726 ( .A(KEYINPUT29), .B(KEYINPUT112), .Z(n653) );
  NAND2_X1 U727 ( .A1(n656), .A2(n661), .ZN(n652) );
  XNOR2_X1 U728 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U729 ( .A(G128), .B(n654), .ZN(G30) );
  XNOR2_X1 U730 ( .A(G143), .B(n655), .ZN(G45) );
  NAND2_X1 U731 ( .A1(n656), .A2(n658), .ZN(n657) );
  XNOR2_X1 U732 ( .A(n657), .B(G146), .ZN(G48) );
  XOR2_X1 U733 ( .A(G113), .B(KEYINPUT113), .Z(n660) );
  NAND2_X1 U734 ( .A1(n662), .A2(n658), .ZN(n659) );
  XNOR2_X1 U735 ( .A(n660), .B(n659), .ZN(G15) );
  NAND2_X1 U736 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U737 ( .A(n663), .B(G116), .ZN(G18) );
  XOR2_X1 U738 ( .A(G125), .B(KEYINPUT37), .Z(n664) );
  XNOR2_X1 U739 ( .A(n665), .B(n664), .ZN(G27) );
  XOR2_X1 U740 ( .A(G134), .B(n666), .Z(G36) );
  XNOR2_X1 U741 ( .A(G140), .B(n667), .ZN(G42) );
  XNOR2_X1 U742 ( .A(KEYINPUT120), .B(KEYINPUT53), .ZN(n716) );
  BUF_X1 U743 ( .A(n668), .Z(n754) );
  NOR2_X1 U744 ( .A1(n669), .A2(n754), .ZN(n670) );
  NOR2_X1 U745 ( .A1(KEYINPUT2), .A2(n670), .ZN(n671) );
  NOR2_X1 U746 ( .A1(n672), .A2(n671), .ZN(n714) );
  NAND2_X1 U747 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U748 ( .A(KEYINPUT116), .B(n675), .Z(n676) );
  NOR2_X1 U749 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U750 ( .A(n678), .B(KEYINPUT117), .ZN(n682) );
  NAND2_X1 U751 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U752 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U753 ( .A1(n683), .A2(n379), .ZN(n702) );
  NOR2_X1 U754 ( .A1(n420), .A2(n684), .ZN(n686) );
  XOR2_X1 U755 ( .A(KEYINPUT49), .B(n686), .Z(n687) );
  NOR2_X1 U756 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U757 ( .A(KEYINPUT114), .B(n689), .Z(n694) );
  NOR2_X1 U758 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U759 ( .A(KEYINPUT50), .B(n692), .ZN(n693) );
  NOR2_X1 U760 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U761 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U762 ( .A(KEYINPUT51), .B(n697), .ZN(n699) );
  INV_X1 U763 ( .A(n707), .ZN(n698) );
  NAND2_X1 U764 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U765 ( .A(KEYINPUT115), .B(n700), .Z(n701) );
  NAND2_X1 U766 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U767 ( .A(n703), .B(KEYINPUT118), .ZN(n704) );
  XOR2_X1 U768 ( .A(KEYINPUT52), .B(n704), .Z(n705) );
  NOR2_X1 U769 ( .A1(n706), .A2(n705), .ZN(n710) );
  NOR2_X1 U770 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U771 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U772 ( .A(KEYINPUT119), .B(n711), .Z(n712) );
  NAND2_X1 U773 ( .A1(n712), .A2(n755), .ZN(n713) );
  NOR2_X1 U774 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U775 ( .A(n716), .B(n715), .ZN(G75) );
  NAND2_X1 U776 ( .A1(n732), .A2(G210), .ZN(n720) );
  XOR2_X1 U777 ( .A(KEYINPUT87), .B(KEYINPUT55), .Z(n719) );
  XNOR2_X1 U778 ( .A(n717), .B(KEYINPUT54), .ZN(n718) );
  NAND2_X1 U779 ( .A1(n732), .A2(G469), .ZN(n724) );
  XOR2_X1 U780 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n723) );
  XNOR2_X1 U781 ( .A(n721), .B(KEYINPUT121), .ZN(n722) );
  NAND2_X1 U782 ( .A1(n732), .A2(G475), .ZN(n726) );
  XOR2_X1 U783 ( .A(n727), .B(KEYINPUT123), .Z(n729) );
  NAND2_X1 U784 ( .A1(n732), .A2(G478), .ZN(n728) );
  XNOR2_X1 U785 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X1 U786 ( .A1(n736), .A2(n730), .ZN(G63) );
  XNOR2_X1 U787 ( .A(n731), .B(KEYINPUT124), .ZN(n734) );
  NAND2_X1 U788 ( .A1(G217), .A2(n732), .ZN(n733) );
  XNOR2_X1 U789 ( .A(n734), .B(n733), .ZN(n735) );
  NOR2_X1 U790 ( .A1(n736), .A2(n735), .ZN(G66) );
  XOR2_X1 U791 ( .A(G101), .B(n737), .Z(n738) );
  XNOR2_X1 U792 ( .A(n739), .B(n738), .ZN(n740) );
  NOR2_X1 U793 ( .A1(n741), .A2(n740), .ZN(n751) );
  XOR2_X1 U794 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n743) );
  NAND2_X1 U795 ( .A1(G224), .A2(G953), .ZN(n742) );
  XNOR2_X1 U796 ( .A(n743), .B(n742), .ZN(n744) );
  NAND2_X1 U797 ( .A1(G898), .A2(n744), .ZN(n745) );
  XNOR2_X1 U798 ( .A(n745), .B(KEYINPUT126), .ZN(n748) );
  NAND2_X1 U799 ( .A1(n746), .A2(n755), .ZN(n747) );
  NAND2_X1 U800 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U801 ( .A(n749), .B(KEYINPUT127), .Z(n750) );
  XNOR2_X1 U802 ( .A(n751), .B(n750), .ZN(G69) );
  XNOR2_X1 U803 ( .A(n753), .B(n752), .ZN(n757) );
  XNOR2_X1 U804 ( .A(n757), .B(n754), .ZN(n756) );
  NAND2_X1 U805 ( .A1(n756), .A2(n755), .ZN(n761) );
  XNOR2_X1 U806 ( .A(G227), .B(n757), .ZN(n758) );
  NAND2_X1 U807 ( .A1(n758), .A2(G900), .ZN(n759) );
  NAND2_X1 U808 ( .A1(n759), .A2(G953), .ZN(n760) );
  NAND2_X1 U809 ( .A1(n761), .A2(n760), .ZN(G72) );
  XOR2_X1 U810 ( .A(n762), .B(G137), .Z(G39) );
  XOR2_X1 U811 ( .A(n763), .B(G122), .Z(G24) );
  XNOR2_X1 U812 ( .A(n764), .B(G119), .ZN(G21) );
  XOR2_X1 U813 ( .A(n765), .B(G131), .Z(G33) );
endmodule

