//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n548, new_n549, new_n551, new_n552, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1192, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  AOI22_X1  g029(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT65), .ZN(G319));
  INV_X1    g031(.A(G2105), .ZN(new_n457));
  XNOR2_X1  g032(.A(KEYINPUT3), .B(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G125), .ZN(new_n459));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n458), .A2(G137), .ZN(new_n463));
  NAND2_X1  g038(.A1(G101), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(new_n467), .B(KEYINPUT66), .ZN(G160));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(new_n457), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n473), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n457), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  NAND4_X1  g056(.A1(new_n470), .A2(new_n472), .A3(G138), .A4(new_n457), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n458), .A2(KEYINPUT4), .A3(G138), .A4(new_n457), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(G114), .A2(G2104), .ZN(new_n488));
  INV_X1    g063(.A(G126), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n473), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n469), .A2(G2105), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n490), .A2(G2105), .B1(G102), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G164));
  NAND2_X1  g069(.A1(G75), .A2(G543), .ZN(new_n495));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT5), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G62), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n495), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(new_n496), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n502), .A2(G651), .B1(new_n506), .B2(G50), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n497), .B(new_n499), .C1(new_n503), .C2(new_n504), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT67), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n507), .B1(new_n508), .B2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND3_X1  g092(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n506), .A2(G51), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n510), .A2(G89), .A3(new_n514), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT69), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT68), .B(KEYINPUT7), .ZN(new_n522));
  AND3_X1   g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n522), .B(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n520), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n521), .B1(new_n520), .B2(new_n524), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n518), .B(new_n519), .C1(new_n526), .C2(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  INV_X1    g104(.A(new_n515), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G90), .ZN(new_n531));
  NAND2_X1  g106(.A1(G77), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G64), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n500), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n534), .A2(G651), .B1(new_n506), .B2(G52), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n531), .A2(new_n535), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  NAND2_X1  g112(.A1(G68), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G56), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n500), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n511), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  OAI221_X1 g119(.A(new_n541), .B1(new_n542), .B2(new_n543), .C1(new_n515), .C2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(new_n549));
  XOR2_X1   g124(.A(new_n549), .B(KEYINPUT70), .Z(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(G188));
  NAND3_X1  g128(.A1(new_n506), .A2(KEYINPUT9), .A3(G53), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n543), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n554), .A2(new_n557), .A3(KEYINPUT71), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  XOR2_X1   g138(.A(KEYINPUT72), .B(G65), .Z(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n564), .B2(new_n500), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n510), .A2(G91), .A3(new_n514), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n562), .A2(new_n569), .ZN(G299));
  OAI21_X1  g145(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n506), .A2(G49), .ZN(new_n572));
  INV_X1    g147(.A(G87), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n571), .B(new_n572), .C1(new_n515), .C2(new_n573), .ZN(G288));
  NAND3_X1  g149(.A1(new_n510), .A2(G86), .A3(new_n514), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n506), .A2(G48), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n497), .A2(new_n499), .A3(G61), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT73), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n497), .A2(new_n499), .A3(KEYINPUT73), .A4(G61), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G651), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n577), .A2(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(new_n506), .A2(G47), .ZN(new_n586));
  INV_X1    g161(.A(G651), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  XOR2_X1   g163(.A(KEYINPUT74), .B(G85), .Z(new_n589));
  OAI221_X1 g164(.A(new_n586), .B1(new_n587), .B2(new_n588), .C1(new_n515), .C2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  INV_X1    g166(.A(G92), .ZN(new_n592));
  OR3_X1    g167(.A1(new_n515), .A2(KEYINPUT10), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n500), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(new_n506), .B2(G54), .ZN(new_n597));
  OAI21_X1  g172(.A(KEYINPUT10), .B1(new_n515), .B2(new_n592), .ZN(new_n598));
  AND3_X1   g173(.A1(new_n593), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n591), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n591), .B1(new_n599), .B2(G868), .ZN(G321));
  NAND2_X1  g176(.A1(G286), .A2(G868), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n568), .B1(new_n560), .B2(new_n561), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(G868), .B2(new_n603), .ZN(G297));
  OAI21_X1  g179(.A(new_n602), .B1(G868), .B2(new_n603), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n599), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g186(.A(new_n476), .ZN(new_n612));
  INV_X1    g187(.A(G135), .ZN(new_n613));
  OR3_X1    g188(.A1(new_n612), .A2(KEYINPUT75), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(KEYINPUT75), .B1(new_n612), .B2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n474), .A2(G123), .ZN(new_n616));
  OR2_X1    g191(.A1(G99), .A2(G2105), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n617), .B(G2104), .C1(G111), .C2(new_n457), .ZN(new_n618));
  NAND4_X1  g193(.A1(new_n614), .A2(new_n615), .A3(new_n616), .A4(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(G2096), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n458), .A2(new_n491), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2100), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n620), .A2(new_n624), .ZN(G156));
  XOR2_X1   g200(.A(KEYINPUT15), .B(G2435), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT77), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n627), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT14), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2451), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n631), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n637), .B(new_n638), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G14), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(G401));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2067), .B(G2678), .Z(new_n644));
  NOR2_X1   g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n643), .A2(new_n644), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT78), .B(KEYINPUT17), .Z(new_n648));
  NAND3_X1  g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT18), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2072), .B(G2078), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n651), .B(new_n652), .C1(new_n650), .C2(new_n645), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n652), .B2(new_n651), .ZN(new_n654));
  XOR2_X1   g229(.A(G2096), .B(G2100), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G227));
  XNOR2_X1  g232(.A(G1956), .B(G2474), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT79), .ZN(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  AND2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n659), .A2(new_n660), .ZN(new_n666));
  AOI22_X1  g241(.A1(new_n664), .A2(new_n665), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  OR3_X1    g242(.A1(new_n661), .A2(new_n666), .A3(new_n663), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n667), .B(new_n668), .C1(new_n665), .C2(new_n664), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT21), .B(G1986), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G1991), .B(G1996), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT22), .B(G1981), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n673), .B(new_n674), .Z(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G229));
  INV_X1    g251(.A(G29), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G27), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(G164), .B2(new_n677), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT92), .B(G2078), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  AND3_X1   g257(.A1(new_n682), .A2(KEYINPUT23), .A3(G20), .ZN(new_n683));
  AOI21_X1  g258(.A(KEYINPUT23), .B1(new_n682), .B2(G20), .ZN(new_n684));
  AOI211_X1 g259(.A(new_n683), .B(new_n684), .C1(G299), .C2(G16), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1956), .ZN(new_n686));
  OR2_X1    g261(.A1(KEYINPUT24), .A2(G34), .ZN(new_n687));
  NAND2_X1  g262(.A1(KEYINPUT24), .A2(G34), .ZN(new_n688));
  AOI21_X1  g263(.A(G29), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(G160), .B2(G29), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n686), .B1(G2084), .B2(new_n690), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n677), .A2(G26), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n474), .A2(G128), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n476), .A2(G140), .ZN(new_n694));
  OR2_X1    g269(.A1(G104), .A2(G2105), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n695), .B(G2104), .C1(G116), .C2(new_n457), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT86), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n692), .B1(new_n698), .B2(G29), .ZN(new_n699));
  MUX2_X1   g274(.A(new_n692), .B(new_n699), .S(KEYINPUT28), .Z(new_n700));
  XOR2_X1   g275(.A(KEYINPUT87), .B(G2067), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n691), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n599), .A2(G16), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G4), .B2(G16), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT85), .B(G1348), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT31), .B(G11), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n705), .A2(new_n706), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n677), .A2(G35), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G162), .B2(new_n677), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n712), .A2(KEYINPUT29), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(KEYINPUT29), .ZN(new_n714));
  OR3_X1    g289(.A1(new_n713), .A2(new_n714), .A3(G2090), .ZN(new_n715));
  OAI21_X1  g290(.A(G2090), .B1(new_n713), .B2(new_n714), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT30), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(G28), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(G28), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n718), .A2(new_n719), .A3(new_n677), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n715), .A2(new_n716), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(G29), .A2(G32), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n476), .A2(G141), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n474), .A2(G129), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n491), .A2(G105), .ZN(new_n725));
  NAND3_X1  g300(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT26), .Z(new_n727));
  NAND4_X1  g302(.A1(new_n723), .A2(new_n724), .A3(new_n725), .A4(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n722), .B1(new_n729), .B2(G29), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT27), .B(G1996), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n619), .A2(new_n677), .ZN(new_n733));
  NOR4_X1   g308(.A1(new_n710), .A2(new_n721), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n682), .A2(G21), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G168), .B2(new_n682), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT90), .B(G1966), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT91), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G5), .B2(G16), .ZN(new_n740));
  OR3_X1    g315(.A1(new_n739), .A2(G5), .A3(G16), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n740), .B(new_n741), .C1(G301), .C2(new_n682), .ZN(new_n742));
  INV_X1    g317(.A(G1961), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n677), .A2(G33), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n476), .A2(G139), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT88), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n491), .A2(G103), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT25), .Z(new_n750));
  AOI22_X1  g325(.A1(new_n458), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT89), .Z(new_n752));
  OAI211_X1 g327(.A(new_n748), .B(new_n750), .C1(new_n457), .C2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n746), .B1(new_n753), .B2(G29), .ZN(new_n754));
  INV_X1    g329(.A(G2072), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n745), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI211_X1 g331(.A(new_n744), .B(new_n756), .C1(G2084), .C2(new_n690), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n703), .A2(new_n734), .A3(new_n738), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n474), .A2(G119), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT80), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n476), .A2(G131), .ZN(new_n761));
  NOR2_X1   g336(.A1(G95), .A2(G2105), .ZN(new_n762));
  OAI21_X1  g337(.A(G2104), .B1(new_n457), .B2(G107), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  MUX2_X1   g340(.A(G25), .B(new_n765), .S(G29), .Z(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT35), .B(G1991), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT81), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n682), .B2(G24), .ZN(new_n770));
  AND3_X1   g345(.A1(new_n769), .A2(new_n682), .A3(G24), .ZN(new_n771));
  AOI211_X1 g346(.A(new_n770), .B(new_n771), .C1(G290), .C2(G16), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1986), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n766), .A2(new_n767), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n768), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G6), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(G16), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G305), .B2(G16), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(KEYINPUT82), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT32), .B(G1981), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n779), .A2(KEYINPUT82), .ZN(new_n782));
  AND3_X1   g357(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n781), .B1(new_n780), .B2(new_n782), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(G23), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n786), .A2(G16), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G288), .B2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n788), .A2(new_n790), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT33), .B(G1976), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  OR3_X1    g369(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n682), .A2(G22), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G166), .B2(new_n682), .ZN(new_n797));
  INV_X1    g372(.A(G1971), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n794), .B1(new_n791), .B2(new_n792), .ZN(new_n800));
  AND3_X1   g375(.A1(new_n795), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  AND3_X1   g376(.A1(new_n785), .A2(KEYINPUT34), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(KEYINPUT34), .B1(new_n785), .B2(new_n801), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n776), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(KEYINPUT36), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT36), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n806), .B(new_n776), .C1(new_n802), .C2(new_n803), .ZN(new_n807));
  AOI211_X1 g382(.A(new_n681), .B(new_n758), .C1(new_n805), .C2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT93), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n754), .A2(new_n755), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n682), .A2(G19), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n546), .B2(new_n682), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(G1341), .Z(new_n813));
  NAND4_X1  g388(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n758), .B1(new_n805), .B2(new_n807), .ZN(new_n815));
  INV_X1    g390(.A(new_n681), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n815), .A2(new_n810), .A3(new_n813), .A4(new_n816), .ZN(G150));
  NAND2_X1  g392(.A1(G150), .A2(KEYINPUT93), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n814), .A2(new_n818), .ZN(G311));
  INV_X1    g394(.A(G67), .ZN(new_n820));
  INV_X1    g395(.A(G80), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n500), .A2(new_n820), .B1(new_n821), .B2(new_n496), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT94), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI221_X1 g399(.A(KEYINPUT94), .B1(new_n821), .B2(new_n496), .C1(new_n500), .C2(new_n820), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n824), .A2(G651), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n506), .A2(G55), .ZN(new_n827));
  INV_X1    g402(.A(G93), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n826), .B(new_n827), .C1(new_n828), .C2(new_n515), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n545), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n599), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n834), .A2(G860), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT95), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n829), .A2(G860), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT96), .B(KEYINPUT37), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n836), .A2(new_n839), .ZN(G145));
  XOR2_X1   g415(.A(KEYINPUT100), .B(G37), .Z(new_n841));
  INV_X1    g416(.A(KEYINPUT99), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT97), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n484), .A2(new_n485), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n843), .B1(new_n484), .B2(new_n485), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n492), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n728), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n698), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n848), .A2(new_n753), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n753), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI22_X1  g426(.A1(G130), .A2(new_n474), .B1(new_n476), .B2(G142), .ZN(new_n852));
  OAI21_X1  g427(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n853), .A2(KEYINPUT98), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(KEYINPUT98), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n854), .B(new_n855), .C1(G118), .C2(new_n457), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n622), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n765), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n842), .B1(new_n851), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n859), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n849), .A2(KEYINPUT99), .A3(new_n850), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n851), .A2(new_n859), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(G160), .B(new_n619), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n480), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n841), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n851), .B(KEYINPUT101), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n859), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n871), .A2(new_n863), .A3(new_n867), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g449(.A1(new_n829), .A2(G868), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n599), .A2(new_n603), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n593), .A2(new_n597), .A3(new_n598), .ZN(new_n877));
  NAND2_X1  g452(.A1(G299), .A2(new_n877), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n876), .A2(new_n878), .A3(KEYINPUT41), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT41), .B1(new_n876), .B2(new_n878), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n876), .A2(new_n878), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n830), .B(new_n608), .ZN(new_n884));
  MUX2_X1   g459(.A(new_n881), .B(new_n883), .S(new_n884), .Z(new_n885));
  AND2_X1   g460(.A1(new_n885), .A2(KEYINPUT103), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(KEYINPUT103), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(G303), .B(G288), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(G305), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(G290), .ZN(new_n891));
  XOR2_X1   g466(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  MUX2_X1   g468(.A(new_n886), .B(new_n888), .S(new_n893), .Z(new_n894));
  AOI21_X1  g469(.A(new_n875), .B1(new_n894), .B2(G868), .ZN(G295));
  AOI21_X1  g470(.A(new_n875), .B1(new_n894), .B2(G868), .ZN(G331));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n897));
  NAND2_X1  g472(.A1(G286), .A2(G171), .ZN(new_n898));
  INV_X1    g473(.A(new_n527), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n525), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n900), .A2(new_n518), .A3(new_n519), .A4(G301), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n546), .B(new_n829), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n830), .A2(new_n898), .A3(new_n901), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n881), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n904), .A2(new_n883), .A3(new_n905), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(KEYINPUT106), .A3(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n890), .B(G290), .Z(new_n910));
  OR2_X1    g485(.A1(new_n908), .A2(KEYINPUT106), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n841), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n907), .A2(KEYINPUT104), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n881), .A2(new_n906), .A3(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n915), .A2(new_n891), .A3(new_n917), .A4(new_n908), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n906), .ZN(new_n921));
  AOI22_X1  g496(.A1(new_n907), .A2(KEYINPUT104), .B1(new_n921), .B2(new_n883), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n922), .A2(KEYINPUT105), .A3(new_n891), .A4(new_n917), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n914), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n897), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n920), .A2(new_n923), .ZN(new_n927));
  INV_X1    g502(.A(new_n914), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(KEYINPUT107), .A3(KEYINPUT43), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n922), .A2(new_n917), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n932), .B2(new_n910), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n927), .A2(new_n925), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT44), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n927), .A2(new_n925), .A3(new_n928), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n925), .B1(new_n927), .B2(new_n933), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI22_X1  g513(.A1(new_n931), .A2(new_n935), .B1(new_n938), .B2(KEYINPUT44), .ZN(G397));
  XOR2_X1   g514(.A(KEYINPUT108), .B(G1384), .Z(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n846), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n943));
  INV_X1    g518(.A(G40), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n461), .A2(new_n465), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n942), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G1996), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n947), .A2(KEYINPUT109), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n950), .B1(new_n946), .B2(G1996), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n729), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT110), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n698), .B(G2067), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n729), .A2(new_n948), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n947), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n952), .A2(new_n958), .A3(new_n729), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n954), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n765), .B(new_n767), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT111), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n947), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(G290), .B(G1986), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n964), .B1(new_n947), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1384), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n846), .A2(new_n967), .A3(new_n945), .ZN(new_n968));
  XNOR2_X1  g543(.A(KEYINPUT114), .B(G8), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n530), .A2(G87), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n970), .A2(G1976), .A3(new_n571), .A4(new_n572), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n973));
  INV_X1    g548(.A(G288), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n974), .A2(G1976), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n972), .A2(KEYINPUT115), .A3(new_n973), .A4(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n978), .A2(KEYINPUT52), .A3(new_n975), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT115), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(new_n978), .B2(KEYINPUT52), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n977), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1981), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n584), .A2(new_n983), .A3(new_n575), .A4(new_n576), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT116), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n577), .A2(KEYINPUT116), .A3(new_n983), .A4(new_n584), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(G305), .A2(G1981), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n988), .A2(KEYINPUT49), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT49), .B1(new_n988), .B2(new_n989), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n968), .A2(new_n969), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT117), .B1(new_n982), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n981), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n972), .A2(new_n973), .A3(new_n976), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n988), .A2(new_n989), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT49), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n992), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n988), .A2(KEYINPUT49), .A3(new_n989), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n997), .A2(new_n1003), .A3(new_n1004), .A4(new_n977), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n994), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G303), .A2(G8), .ZN(new_n1007));
  XOR2_X1   g582(.A(new_n1007), .B(KEYINPUT55), .Z(new_n1008));
  AOI21_X1  g583(.A(G1384), .B1(new_n487), .B2(new_n492), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n945), .B1(new_n1009), .B2(KEYINPUT45), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n486), .A2(KEYINPUT97), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n484), .A2(new_n485), .A3(new_n843), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n940), .B1(new_n1015), .B2(new_n492), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1012), .B1(new_n1016), .B2(KEYINPUT45), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n846), .A2(new_n1012), .A3(KEYINPUT45), .A4(new_n941), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1011), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n846), .A2(KEYINPUT45), .A3(new_n941), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT112), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n1018), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1025), .A2(KEYINPUT113), .A3(new_n1011), .ZN(new_n1026));
  AOI21_X1  g601(.A(G1971), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n493), .A2(new_n967), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT50), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n846), .A2(new_n1030), .A3(new_n967), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n1031), .A3(new_n945), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(G2090), .ZN(new_n1033));
  OAI211_X1 g608(.A(G8), .B(new_n1008), .C1(new_n1027), .C2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n969), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT113), .B1(new_n1025), .B2(new_n1011), .ZN(new_n1036));
  AOI211_X1 g611(.A(new_n1021), .B(new_n1010), .C1(new_n1024), .C2(new_n1018), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n798), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n945), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(new_n1009), .B2(new_n1030), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n846), .A2(new_n967), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT50), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n1043), .A2(G2090), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1035), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1006), .B(new_n1034), .C1(new_n1008), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1009), .A2(KEYINPUT45), .ZN(new_n1048));
  AOI21_X1  g623(.A(G1384), .B1(new_n1015), .B2(new_n492), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n945), .B(new_n1048), .C1(new_n1049), .C2(KEYINPUT45), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n1051));
  OR3_X1    g626(.A1(new_n1050), .A2(new_n1051), .A3(G2078), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1032), .A2(new_n743), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1036), .A2(new_n1037), .A3(G2078), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT122), .B(KEYINPUT53), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1052), .B(new_n1053), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1056), .A2(G171), .ZN(new_n1057));
  INV_X1    g632(.A(G2084), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1029), .A2(new_n1031), .A3(new_n1058), .A4(new_n945), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1048), .A2(new_n945), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT45), .B1(new_n846), .B2(new_n967), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n737), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1050), .A2(KEYINPUT118), .A3(new_n737), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1061), .A2(new_n1062), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI211_X1 g644(.A(KEYINPUT51), .B(new_n1035), .C1(new_n1069), .C2(G168), .ZN(new_n1070));
  INV_X1    g645(.A(G8), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1071), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(G286), .A2(new_n969), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT51), .ZN(new_n1076));
  OAI22_X1  g651(.A1(new_n1074), .A2(new_n1076), .B1(new_n1069), .B2(new_n1075), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT62), .B1(new_n1070), .B2(new_n1077), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT62), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT51), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1081), .B(new_n969), .C1(new_n1082), .C2(G286), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(G286), .A3(new_n969), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1079), .A2(new_n1080), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1047), .A2(new_n1057), .A3(new_n1078), .A4(new_n1085), .ZN(new_n1086));
  OR3_X1    g661(.A1(new_n993), .A2(G1976), .A3(G288), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n992), .B1(new_n1087), .B2(new_n988), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1034), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n982), .A2(new_n993), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT56), .B(G2072), .Z(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1025), .A2(new_n1011), .A3(new_n1093), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT120), .B(G1956), .Z(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1096), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n558), .A2(KEYINPUT57), .ZN(new_n1099));
  AOI22_X1  g674(.A1(G299), .A2(KEYINPUT57), .B1(new_n569), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1094), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n968), .A2(G2067), .ZN(new_n1102));
  INV_X1    g677(.A(G1348), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n1032), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1101), .A2(new_n599), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1100), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n1010), .B(new_n1092), .C1(new_n1024), .C2(new_n1018), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1107), .B1(new_n1108), .B2(new_n1097), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1106), .A2(KEYINPUT121), .A3(new_n1109), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1108), .A2(new_n1107), .A3(new_n1097), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1100), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1104), .A2(new_n599), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n1118), .A2(KEYINPUT60), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1104), .A2(new_n599), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1120), .A2(KEYINPUT60), .A3(new_n1118), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1117), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1109), .A2(new_n1101), .A3(KEYINPUT61), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1025), .A2(new_n948), .A3(new_n1011), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT58), .B(G1341), .Z(new_n1126));
  NAND2_X1  g701(.A1(new_n968), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1124), .B1(new_n1128), .B2(new_n546), .ZN(new_n1129));
  AOI211_X1 g704(.A(KEYINPUT59), .B(new_n545), .C1(new_n1125), .C2(new_n1127), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1123), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1112), .B(new_n1113), .C1(new_n1122), .C2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1079), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1047), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1135));
  INV_X1    g710(.A(G2078), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1055), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1039), .B1(new_n942), .B2(new_n943), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT124), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1051), .A2(G2078), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1138), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n1142), .A2(new_n1143), .B1(new_n1024), .B2(new_n1018), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1053), .A2(KEYINPUT123), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1032), .A2(new_n1147), .A3(new_n743), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT125), .B1(new_n1137), .B2(new_n1150), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1141), .A2(new_n1144), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1152), .B(new_n1153), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1151), .A2(G171), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1156), .B1(new_n1056), .B2(G301), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT54), .B1(new_n1056), .B2(G171), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1152), .B(G301), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1155), .A2(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1086), .B(new_n1091), .C1(new_n1134), .C2(new_n1160), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n1069), .A2(G286), .A3(new_n1035), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1033), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1071), .B1(new_n1038), .B2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1162), .B(new_n1090), .C1(new_n1164), .C2(new_n1008), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT63), .ZN(new_n1166));
  NOR3_X1   g741(.A1(new_n1165), .A2(new_n1089), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1047), .A2(new_n1162), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1167), .B1(new_n1168), .B2(new_n1166), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n966), .B1(new_n1161), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n947), .B1(new_n955), .B2(new_n728), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n949), .A2(KEYINPUT46), .A3(new_n951), .ZN(new_n1172));
  AOI21_X1  g747(.A(KEYINPUT46), .B1(new_n949), .B2(new_n951), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT47), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n946), .A2(G1986), .A3(G290), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n1176), .B(KEYINPUT48), .Z(new_n1177));
  NAND3_X1  g752(.A1(new_n960), .A2(new_n963), .A3(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n698), .A2(G2067), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n765), .A2(new_n767), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1180), .B(KEYINPUT126), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1179), .B1(new_n960), .B2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1175), .B(new_n1178), .C1(new_n1182), .C2(new_n946), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT127), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1170), .A2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g760(.A(new_n455), .B(new_n675), .C1(new_n936), .C2(new_n937), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n640), .A2(new_n656), .ZN(new_n1188));
  INV_X1    g762(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g763(.A1(new_n873), .A2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g764(.A1(new_n1187), .A2(new_n1190), .ZN(G308));
  OR2_X1    g765(.A1(new_n936), .A2(new_n937), .ZN(new_n1192));
  AOI21_X1  g766(.A(new_n1188), .B1(new_n869), .B2(new_n872), .ZN(new_n1193));
  NAND4_X1  g767(.A1(new_n1192), .A2(new_n1193), .A3(new_n455), .A4(new_n675), .ZN(G225));
endmodule


