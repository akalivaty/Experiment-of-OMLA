//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 1 1 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n865, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n192), .A3(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(KEYINPUT1), .A3(G146), .ZN(new_n196));
  XNOR2_X1  g010(.A(G143), .B(G146), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n195), .B(new_n196), .C1(G128), .C2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n199), .B1(new_n197), .B2(KEYINPUT64), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n192), .A2(new_n194), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT0), .B(G128), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n200), .A2(new_n204), .ZN(new_n205));
  MUX2_X1   g019(.A(new_n198), .B(new_n205), .S(G125), .Z(new_n206));
  INV_X1    g020(.A(G224), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G953), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n206), .B(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT67), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT66), .B(G116), .ZN(new_n211));
  INV_X1    g025(.A(G119), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(G116), .ZN(new_n214));
  INV_X1    g028(.A(G116), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n215), .A2(KEYINPUT66), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(KEYINPUT66), .ZN(new_n217));
  OAI211_X1 g031(.A(KEYINPUT67), .B(G119), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n213), .A2(new_n214), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT68), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n213), .A2(new_n218), .A3(new_n221), .A4(new_n214), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(KEYINPUT5), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G113), .ZN(new_n224));
  INV_X1    g038(.A(new_n214), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT5), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT79), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT2), .B(G113), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n219), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G104), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT77), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT77), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G104), .ZN(new_n237));
  INV_X1    g051(.A(G107), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT3), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n235), .A2(new_n237), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G107), .ZN(new_n242));
  INV_X1    g056(.A(G101), .ZN(new_n243));
  OR3_X1    g057(.A1(new_n234), .A2(KEYINPUT3), .A3(G107), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n240), .A2(new_n242), .A3(new_n243), .A4(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n239), .B1(G104), .B2(new_n238), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G101), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n223), .A2(KEYINPUT79), .A3(new_n227), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n230), .A2(new_n233), .A3(new_n249), .A4(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n220), .A2(new_n222), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n231), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n233), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n240), .A2(new_n242), .A3(new_n244), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n256), .A3(G101), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(G101), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT4), .A3(new_n245), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n254), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n251), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT81), .ZN(new_n262));
  XOR2_X1   g076(.A(G110), .B(G122), .Z(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT6), .ZN(new_n265));
  INV_X1    g079(.A(new_n263), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n251), .B2(new_n260), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n262), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n251), .A2(new_n260), .A3(new_n266), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT80), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n261), .A2(new_n263), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT80), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n251), .A2(new_n274), .A3(new_n260), .A4(new_n266), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n209), .B1(new_n270), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n272), .A2(new_n275), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n230), .A2(new_n233), .A3(new_n248), .A4(new_n250), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n227), .B1(new_n219), .B2(new_n226), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n233), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n249), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n263), .B(KEYINPUT82), .ZN(new_n283));
  XOR2_X1   g097(.A(new_n283), .B(KEYINPUT8), .Z(new_n284));
  NAND3_X1  g098(.A1(new_n279), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT7), .B1(new_n207), .B2(G953), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n206), .B(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n278), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n188), .B1(new_n277), .B2(new_n290), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n267), .A2(new_n262), .A3(new_n268), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n268), .B1(new_n267), .B2(new_n262), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n276), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n209), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n285), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n297), .B1(new_n272), .B2(new_n275), .ZN(new_n298));
  AOI21_X1  g112(.A(G902), .B1(new_n298), .B2(new_n287), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n296), .A2(new_n299), .A3(new_n187), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n291), .A2(new_n300), .A3(KEYINPUT83), .ZN(new_n301));
  NAND2_X1  g115(.A1(G234), .A2(G237), .ZN(new_n302));
  INV_X1    g116(.A(G953), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(G952), .A3(new_n303), .ZN(new_n304));
  XOR2_X1   g118(.A(KEYINPUT21), .B(G898), .Z(new_n305));
  NAND3_X1  g119(.A1(new_n302), .A2(G902), .A3(G953), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT83), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n308), .B(new_n188), .C1(new_n277), .C2(new_n290), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n301), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G469), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n259), .A2(new_n205), .A3(new_n257), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n245), .A2(new_n247), .A3(new_n198), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT10), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT11), .ZN(new_n315));
  INV_X1    g129(.A(G134), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n315), .B1(new_n316), .B2(G137), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(G137), .ZN(new_n318));
  INV_X1    g132(.A(G137), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(KEYINPUT11), .A3(G134), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n317), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G131), .ZN(new_n322));
  INV_X1    g136(.A(G131), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n317), .A2(new_n320), .A3(new_n323), .A4(new_n318), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n245), .A2(new_n247), .A3(new_n198), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT10), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n312), .A2(new_n314), .A3(new_n326), .A4(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n303), .A2(G227), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(G140), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT76), .B(G110), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n198), .B1(new_n245), .B2(new_n247), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n325), .B1(new_n313), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT12), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n339), .B(new_n340), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n312), .A2(new_n329), .A3(new_n314), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT78), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n312), .A2(new_n314), .A3(new_n345), .A4(new_n329), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n325), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n335), .B1(new_n347), .B2(new_n330), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n311), .B(new_n289), .C1(new_n342), .C2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n335), .B1(new_n341), .B2(new_n330), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(new_n337), .B2(new_n347), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G469), .ZN(new_n352));
  NAND2_X1  g166(.A1(G469), .A2(G902), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n349), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  XOR2_X1   g168(.A(KEYINPUT9), .B(G234), .Z(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(G221), .B1(new_n356), .B2(G902), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT90), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n189), .A2(G143), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT13), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n189), .A2(G143), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n360), .A2(KEYINPUT90), .A3(KEYINPUT13), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n360), .A2(KEYINPUT13), .ZN(new_n367));
  OAI21_X1  g181(.A(G134), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n361), .A2(new_n364), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n316), .ZN(new_n370));
  INV_X1    g184(.A(G122), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G116), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n372), .B1(new_n211), .B2(new_n371), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n373), .A2(G107), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(G107), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n368), .B(new_n370), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n369), .B(new_n316), .ZN(new_n377));
  OAI211_X1 g191(.A(KEYINPUT14), .B(G122), .C1(new_n216), .C2(new_n217), .ZN(new_n378));
  OAI211_X1 g192(.A(G107), .B(new_n378), .C1(new_n373), .C2(KEYINPUT14), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n377), .B(new_n379), .C1(G107), .C2(new_n373), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G217), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n356), .A2(new_n382), .A3(G953), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n376), .A2(new_n380), .A3(new_n383), .ZN(new_n386));
  AOI21_X1  g200(.A(G902), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT15), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G478), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT91), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(KEYINPUT91), .A3(G478), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n387), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT92), .ZN(new_n394));
  OR2_X1    g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OR2_X1    g209(.A1(new_n387), .A2(new_n389), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n394), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G237), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(new_n303), .A3(G214), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n193), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n399), .A2(new_n303), .A3(G143), .A4(G214), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT85), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT85), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n405), .A2(KEYINPUT18), .A3(G131), .A4(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(G125), .B(G140), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n191), .ZN(new_n410));
  NAND2_X1  g224(.A1(KEYINPUT73), .A2(G125), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(G140), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n410), .B1(new_n413), .B2(new_n191), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT86), .ZN(new_n415));
  NAND2_X1  g229(.A1(KEYINPUT18), .A2(G131), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n404), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n415), .B1(new_n404), .B2(new_n416), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n408), .B(new_n414), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G140), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT16), .B1(new_n420), .B2(G125), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n412), .B2(KEYINPUT16), .ZN(new_n422));
  OR2_X1    g236(.A1(new_n422), .A2(new_n191), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n403), .B(G131), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n409), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT19), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n426), .B1(new_n413), .B2(new_n427), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n423), .B(new_n424), .C1(G146), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n419), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(G113), .B(G122), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(new_n234), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n422), .A2(new_n191), .ZN(new_n435));
  OR2_X1    g249(.A1(new_n435), .A2(KEYINPUT74), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(KEYINPUT74), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(new_n423), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n403), .A2(KEYINPUT17), .A3(G131), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n439), .B1(new_n424), .B2(KEYINPUT17), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n432), .B(new_n419), .C1(new_n438), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n434), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n443));
  NOR2_X1   g257(.A1(G475), .A2(G902), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n444), .B(KEYINPUT88), .Z(new_n445));
  AND3_X1   g259(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  XOR2_X1   g260(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(new_n442), .B2(new_n445), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n419), .B1(new_n438), .B2(new_n440), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n433), .ZN(new_n451));
  AOI21_X1  g265(.A(G902), .B1(new_n451), .B2(new_n441), .ZN(new_n452));
  XOR2_X1   g266(.A(KEYINPUT89), .B(G475), .Z(new_n453));
  OAI22_X1  g267(.A1(new_n446), .A2(new_n449), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n398), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n358), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(G214), .B1(G237), .B2(G902), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n310), .A2(KEYINPUT93), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT93), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n301), .A2(new_n458), .A3(new_n307), .A4(new_n309), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n460), .B1(new_n461), .B2(new_n456), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT72), .ZN(new_n464));
  NAND2_X1  g278(.A1(KEYINPUT65), .A2(KEYINPUT30), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT65), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT30), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n318), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n316), .A2(G137), .ZN(new_n470));
  OAI21_X1  g284(.A(G131), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n198), .A2(new_n324), .A3(new_n471), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n322), .A2(new_n324), .B1(new_n200), .B2(new_n204), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n465), .B(new_n468), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n325), .A2(new_n205), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n198), .A2(new_n324), .A3(new_n471), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n475), .A2(new_n476), .A3(new_n466), .A4(new_n467), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n254), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT31), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n399), .A2(new_n303), .A3(G210), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT26), .B(G101), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n483), .B(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n475), .A2(new_n476), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n253), .A2(new_n233), .A3(new_n488), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n479), .A2(new_n480), .A3(new_n486), .A4(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n488), .B1(new_n253), .B2(new_n233), .ZN(new_n492));
  INV_X1    g306(.A(new_n231), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n493), .B1(new_n220), .B2(new_n222), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n494), .A2(new_n232), .A3(new_n487), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n491), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT28), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n489), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n486), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT71), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n490), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n479), .A2(new_n486), .A3(new_n489), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT31), .ZN(new_n503));
  INV_X1    g317(.A(new_n491), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n487), .B1(new_n494), .B2(new_n232), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n504), .B1(new_n489), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n495), .A2(KEYINPUT28), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n485), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n503), .B1(new_n508), .B2(KEYINPUT71), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n464), .B1(new_n501), .B2(new_n509), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n253), .A2(new_n233), .B1(new_n474), .B2(new_n477), .ZN(new_n511));
  NOR4_X1   g325(.A1(new_n511), .A2(new_n495), .A3(KEYINPUT31), .A4(new_n485), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(new_n508), .B2(KEYINPUT71), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n499), .A2(new_n500), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n513), .A2(KEYINPUT72), .A3(new_n514), .A4(new_n503), .ZN(new_n515));
  NOR2_X1   g329(.A1(G472), .A2(G902), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n510), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT32), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n510), .A2(new_n515), .A3(KEYINPUT32), .A4(new_n516), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n496), .A2(new_n486), .A3(new_n498), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n479), .A2(new_n489), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n485), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT29), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n492), .A2(new_n495), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n498), .B1(new_n526), .B2(new_n497), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n486), .A2(KEYINPUT29), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n525), .B(new_n289), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G472), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n519), .A2(new_n520), .A3(new_n530), .ZN(new_n531));
  XOR2_X1   g345(.A(KEYINPUT24), .B(G110), .Z(new_n532));
  XNOR2_X1  g346(.A(G119), .B(G128), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n212), .A2(G128), .ZN(new_n535));
  OR2_X1    g349(.A1(new_n535), .A2(KEYINPUT23), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(KEYINPUT23), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n536), .B(new_n537), .C1(G119), .C2(new_n189), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(G110), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n438), .A2(new_n534), .A3(new_n539), .ZN(new_n540));
  OAI22_X1  g354(.A1(new_n538), .A2(G110), .B1(new_n533), .B2(new_n532), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(new_n423), .A3(new_n410), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT22), .B(G137), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n303), .A2(G221), .A3(G234), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n540), .A2(new_n542), .A3(new_n546), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n289), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT25), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n382), .B1(G234), .B2(new_n289), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT25), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n548), .A2(new_n553), .A3(new_n289), .A4(new_n549), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT75), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n550), .A2(new_n552), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n556), .B1(new_n555), .B2(new_n557), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n531), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n463), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(G101), .ZN(G3));
  INV_X1    g377(.A(new_n458), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n187), .B1(new_n296), .B2(new_n299), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT94), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n291), .A2(new_n300), .A3(KEYINPUT94), .ZN(new_n568));
  INV_X1    g382(.A(G478), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n385), .A2(new_n386), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT33), .B1(new_n383), .B2(KEYINPUT95), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n571), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n385), .A2(new_n386), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n569), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n387), .A2(new_n569), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n569), .A2(new_n289), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n454), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n567), .A2(new_n307), .A3(new_n568), .A4(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n510), .A2(new_n515), .A3(new_n289), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G472), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n584), .A2(new_n517), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(new_n560), .A3(new_n358), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G104), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT96), .B(KEYINPUT34), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(G6));
  NAND2_X1  g404(.A1(new_n442), .A2(new_n445), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(new_n447), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n452), .A2(new_n453), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n592), .A2(new_n594), .A3(new_n307), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n567), .A2(new_n398), .A3(new_n568), .A4(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n586), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT35), .B(G107), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G9));
  NOR2_X1   g413(.A1(new_n547), .A2(KEYINPUT36), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n543), .B(new_n600), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n601), .B(new_n289), .C1(new_n382), .C2(G234), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n555), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n585), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n463), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT37), .B(G110), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G12));
  NAND4_X1  g421(.A1(new_n567), .A2(new_n531), .A3(new_n568), .A4(new_n358), .ZN(new_n608));
  INV_X1    g422(.A(new_n398), .ZN(new_n609));
  INV_X1    g423(.A(new_n603), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n304), .B1(new_n306), .B2(G900), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n592), .A2(new_n594), .A3(new_n611), .ZN(new_n612));
  NOR4_X1   g426(.A1(new_n608), .A2(new_n609), .A3(new_n610), .A4(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(new_n189), .ZN(G30));
  XNOR2_X1  g428(.A(new_n611), .B(KEYINPUT39), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n358), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT40), .ZN(new_n617));
  INV_X1    g431(.A(new_n454), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n502), .B(G472), .C1(new_n486), .C2(new_n526), .ZN(new_n619));
  NAND2_X1  g433(.A1(G472), .A2(G902), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT97), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n519), .A2(new_n520), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR4_X1   g438(.A1(new_n617), .A2(new_n618), .A3(new_n609), .A4(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n301), .A2(KEYINPUT38), .A3(new_n309), .ZN(new_n626));
  AOI21_X1  g440(.A(KEYINPUT38), .B1(new_n301), .B2(new_n309), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n625), .A2(new_n458), .A3(new_n610), .A4(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT98), .B(G143), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G45));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n566), .B(new_n188), .C1(new_n277), .C2(new_n290), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n568), .A2(new_n458), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n531), .A2(new_n358), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n636), .A2(new_n603), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n579), .A2(new_n454), .A3(new_n611), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT99), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n579), .A2(new_n454), .A3(new_n642), .A4(new_n611), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n633), .B1(new_n639), .B2(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n635), .A2(new_n610), .A3(new_n637), .ZN(new_n646));
  INV_X1    g460(.A(new_n644), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(KEYINPUT100), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G146), .ZN(G48));
  INV_X1    g464(.A(new_n582), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n289), .B1(new_n342), .B2(new_n348), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(G469), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n654), .A2(new_n357), .A3(new_n349), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n654), .A2(KEYINPUT101), .A3(new_n357), .A4(new_n349), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n659), .A2(new_n531), .A3(new_n560), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n651), .A2(new_n652), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(KEYINPUT102), .B1(new_n582), .B2(new_n660), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT41), .B(G113), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G15));
  NOR2_X1   g480(.A1(new_n596), .A2(new_n660), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n215), .ZN(G18));
  INV_X1    g482(.A(new_n655), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n567), .A2(new_n307), .A3(new_n568), .A4(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n531), .A2(new_n455), .A3(new_n603), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(new_n212), .ZN(G21));
  NAND4_X1  g487(.A1(new_n567), .A2(new_n454), .A3(new_n568), .A4(new_n398), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n659), .A2(new_n307), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n584), .A2(KEYINPUT105), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n583), .A2(new_n678), .A3(G472), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n527), .A2(new_n485), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n503), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n681), .A2(KEYINPUT104), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(KEYINPUT104), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n490), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n516), .B(KEYINPUT103), .Z(new_n685));
  AOI22_X1  g499(.A1(new_n677), .A2(new_n679), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n555), .A2(new_n557), .ZN(new_n687));
  AOI21_X1  g501(.A(KEYINPUT106), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n684), .A2(new_n685), .ZN(new_n689));
  INV_X1    g503(.A(new_n679), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n678), .B1(new_n583), .B2(G472), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n689), .B(new_n687), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n675), .B(new_n676), .C1(new_n688), .C2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G122), .ZN(G24));
  NOR2_X1   g510(.A1(new_n635), .A2(new_n655), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n686), .B2(new_n603), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n689), .B(new_n603), .C1(new_n690), .C2(new_n691), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(KEYINPUT107), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n647), .B(new_n697), .C1(new_n699), .C2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G125), .ZN(G27));
  INV_X1    g517(.A(new_n687), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n520), .A2(KEYINPUT109), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n519), .A2(new_n520), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n704), .B1(new_n708), .B2(new_n530), .ZN(new_n709));
  AOI211_X1 g523(.A(new_n564), .B(new_n644), .C1(new_n301), .C2(new_n309), .ZN(new_n710));
  XOR2_X1   g524(.A(new_n353), .B(KEYINPUT108), .Z(new_n711));
  NAND3_X1  g525(.A1(new_n349), .A2(new_n352), .A3(new_n711), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n712), .A2(new_n357), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n709), .A2(new_n710), .A3(KEYINPUT42), .A4(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n564), .B1(new_n301), .B2(new_n309), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(new_n561), .A3(new_n647), .A4(new_n713), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT42), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G131), .ZN(G33));
  NOR2_X1   g534(.A1(new_n609), .A2(new_n612), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n715), .A2(new_n561), .A3(new_n721), .A4(new_n713), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G134), .ZN(G36));
  OR2_X1    g537(.A1(new_n454), .A2(KEYINPUT112), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n454), .A2(KEYINPUT112), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n579), .A3(new_n725), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n726), .A2(KEYINPUT43), .ZN(new_n727));
  INV_X1    g541(.A(new_n579), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n728), .A2(KEYINPUT43), .A3(new_n454), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n610), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n727), .A2(new_n729), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n585), .B1(new_n733), .B2(KEYINPUT113), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT44), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n715), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(G469), .B1(new_n351), .B2(KEYINPUT45), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n738), .A2(KEYINPUT110), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n351), .A2(KEYINPUT45), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(KEYINPUT110), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT46), .B1(new_n742), .B2(new_n711), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n743), .A2(KEYINPUT111), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n349), .B1(new_n743), .B2(KEYINPUT111), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n742), .A2(KEYINPUT46), .A3(new_n711), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n357), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n732), .A2(KEYINPUT44), .A3(new_n734), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n737), .A2(new_n615), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G137), .ZN(G39));
  OR2_X1    g566(.A1(new_n744), .A2(new_n745), .ZN(new_n753));
  OAI211_X1 g567(.A(KEYINPUT47), .B(new_n357), .C1(new_n753), .C2(new_n746), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n755), .B1(new_n747), .B2(new_n748), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n531), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n736), .A2(new_n560), .A3(new_n644), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n420), .ZN(G42));
  NAND2_X1  g574(.A1(new_n303), .A2(G952), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n688), .A2(new_n694), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n762), .A2(new_n304), .A3(new_n730), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n761), .B1(new_n763), .B2(new_n697), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n736), .A2(new_n655), .ZN(new_n765));
  INV_X1    g579(.A(new_n304), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n765), .A2(new_n560), .A3(new_n766), .A4(new_n624), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n764), .B1(new_n767), .B2(new_n580), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT117), .Z(new_n769));
  NAND2_X1  g583(.A1(new_n654), .A2(new_n349), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n754), .B(new_n756), .C1(new_n357), .C2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n715), .A3(new_n763), .ZN(new_n772));
  OR3_X1    g586(.A1(new_n767), .A2(new_n454), .A3(new_n579), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n686), .A2(new_n698), .A3(new_n603), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n700), .A2(KEYINPUT107), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n730), .A2(new_n304), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n765), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n629), .A2(new_n655), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n763), .A2(new_n564), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n774), .A2(new_n775), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(new_n780), .A3(new_n772), .A4(new_n773), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT51), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n769), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n459), .B(new_n462), .C1(new_n604), .C2(new_n561), .ZN(new_n790));
  OAI22_X1  g604(.A1(new_n596), .A2(new_n660), .B1(new_n670), .B2(new_n671), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n455), .A2(KEYINPUT114), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n728), .A2(new_n454), .ZN(new_n793));
  AOI22_X1  g607(.A1(new_n792), .A2(new_n793), .B1(KEYINPUT114), .B2(new_n580), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n461), .A2(new_n586), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n790), .A2(new_n796), .A3(new_n664), .A4(new_n695), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n778), .A2(new_n647), .A3(new_n715), .A4(new_n713), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n610), .A2(new_n612), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n715), .A2(new_n638), .A3(new_n609), .A4(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n800), .A2(new_n722), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n719), .A2(new_n798), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n646), .A2(new_n721), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT100), .B1(new_n646), .B2(new_n647), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n608), .A2(new_n633), .A3(new_n610), .A4(new_n644), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n804), .B(new_n702), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n623), .A2(new_n610), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n713), .A2(new_n611), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n674), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n674), .A2(new_n812), .A3(new_n808), .A4(new_n809), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT52), .B1(new_n807), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n810), .B(KEYINPUT115), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n644), .B1(new_n776), .B2(new_n777), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n613), .B1(new_n697), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n816), .A2(new_n649), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n803), .A2(new_n815), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n803), .A2(new_n815), .A3(new_n820), .A4(KEYINPUT53), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n823), .A2(KEYINPUT54), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT54), .B1(new_n823), .B2(new_n824), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n789), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n823), .A2(new_n824), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n823), .A2(KEYINPUT54), .A3(new_n824), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n830), .A2(KEYINPUT116), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n788), .A2(new_n827), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n765), .A2(new_n709), .A3(new_n779), .ZN(new_n834));
  XOR2_X1   g648(.A(new_n834), .B(KEYINPUT48), .Z(new_n835));
  OAI22_X1  g649(.A1(new_n833), .A2(new_n835), .B1(G952), .B2(G953), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n623), .A2(new_n704), .A3(new_n748), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n770), .A2(KEYINPUT49), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n770), .A2(KEYINPUT49), .ZN(new_n839));
  NOR4_X1   g653(.A1(new_n838), .A2(new_n839), .A3(new_n726), .A4(new_n564), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n628), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n836), .A2(new_n841), .ZN(G75));
  NOR2_X1   g656(.A1(new_n303), .A2(G952), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n828), .A2(G210), .A3(G902), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n294), .B(new_n295), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT55), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n847), .A2(KEYINPUT120), .B1(new_n848), .B2(KEYINPUT56), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(KEYINPUT120), .B2(new_n847), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n848), .A2(KEYINPUT56), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n844), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n289), .B1(new_n823), .B2(new_n824), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT56), .B1(new_n853), .B2(G210), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT118), .B1(new_n854), .B2(new_n847), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n856), .B(new_n846), .C1(new_n844), .C2(KEYINPUT56), .ZN(new_n857));
  AOI211_X1 g671(.A(new_n843), .B(new_n852), .C1(new_n855), .C2(new_n857), .ZN(G51));
  NOR2_X1   g672(.A1(new_n825), .A2(new_n826), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n711), .B(KEYINPUT57), .Z(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n861), .B1(new_n348), .B2(new_n342), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n853), .A2(new_n740), .A3(new_n741), .A4(new_n739), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n843), .B1(new_n862), .B2(new_n863), .ZN(G54));
  NAND3_X1  g678(.A1(new_n853), .A2(KEYINPUT58), .A3(G475), .ZN(new_n865));
  INV_X1    g679(.A(new_n442), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n867), .A2(new_n868), .A3(new_n843), .ZN(G60));
  INV_X1    g683(.A(new_n843), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n572), .A2(new_n574), .ZN(new_n871));
  INV_X1    g685(.A(new_n578), .ZN(new_n872));
  XNOR2_X1  g686(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n872), .B(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n859), .A2(new_n871), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n874), .B1(new_n827), .B2(new_n832), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n870), .B(new_n876), .C1(new_n877), .C2(new_n871), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(G63));
  NAND2_X1  g693(.A1(G217), .A2(G902), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT60), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n828), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n548), .A2(new_n549), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n828), .A2(KEYINPUT122), .A3(new_n882), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT122), .B1(new_n828), .B2(new_n882), .ZN(new_n890));
  AOI211_X1 g704(.A(new_n884), .B(new_n881), .C1(new_n823), .C2(new_n824), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n601), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n892), .A3(new_n870), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n889), .A2(new_n892), .A3(KEYINPUT61), .A4(new_n870), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(G66));
  AOI21_X1  g711(.A(new_n303), .B1(new_n305), .B2(G224), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n797), .B2(new_n303), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n270), .B(new_n276), .C1(G898), .C2(new_n303), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n899), .B(new_n900), .Z(G69));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n902));
  INV_X1    g716(.A(new_n807), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n751), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT126), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n749), .A2(new_n615), .A3(new_n675), .A4(new_n709), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n719), .A3(new_n722), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n759), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n905), .A2(new_n908), .A3(new_n303), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n478), .B(new_n428), .Z(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(G900), .B2(G953), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n902), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n630), .A2(new_n649), .A3(new_n819), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n915), .B(new_n916), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n749), .A2(new_n615), .A3(new_n750), .ZN(new_n918));
  AOI22_X1  g732(.A1(new_n757), .A2(new_n758), .B1(new_n918), .B2(new_n737), .ZN(new_n919));
  INV_X1    g733(.A(new_n561), .ZN(new_n920));
  OR4_X1    g734(.A1(new_n920), .A2(new_n736), .A3(new_n616), .A4(new_n794), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n917), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n303), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n914), .B1(new_n923), .B2(new_n911), .ZN(new_n924));
  AOI211_X1 g738(.A(KEYINPUT123), .B(new_n910), .C1(new_n922), .C2(new_n303), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n913), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(G227), .A2(G900), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(G953), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT124), .Z(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n913), .B(new_n929), .C1(new_n924), .C2(new_n925), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(G72));
  XOR2_X1   g747(.A(new_n620), .B(KEYINPUT63), .Z(new_n934));
  NAND2_X1  g748(.A1(new_n905), .A2(new_n908), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n934), .B1(new_n935), .B2(new_n797), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n936), .A2(new_n485), .A3(new_n489), .A4(new_n479), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n934), .B1(new_n922), .B2(new_n797), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n938), .A2(new_n486), .A3(new_n522), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n502), .A2(KEYINPUT127), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(new_n523), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n828), .A2(new_n934), .A3(new_n941), .ZN(new_n942));
  AND4_X1   g756(.A1(new_n870), .A2(new_n937), .A3(new_n939), .A4(new_n942), .ZN(G57));
endmodule


