//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n571,
    new_n572, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n642, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1272, new_n1273, new_n1274;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT66), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT67), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT68), .B1(new_n467), .B2(new_n463), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(new_n474), .A3(G2105), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n466), .B1(new_n468), .B2(new_n475), .ZN(G160));
  NOR2_X1   g051(.A1(new_n469), .A2(new_n470), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n477), .A2(new_n463), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT69), .ZN(G162));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n487), .A2(new_n463), .A3(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n486), .B1(new_n477), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n462), .A2(G126), .A3(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR3_X1   g066(.A1(new_n491), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n462), .A2(KEYINPUT4), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT70), .B1(new_n463), .B2(G114), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n495), .A2(new_n496), .A3(G2105), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n494), .A2(new_n497), .A3(G2104), .A4(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n489), .A2(new_n490), .A3(new_n493), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT73), .B1(new_n502), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT5), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n503), .A2(new_n506), .B1(new_n502), .B2(G543), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(G651), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n509), .A2(KEYINPUT72), .A3(KEYINPUT6), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n513), .A2(new_n514), .B1(new_n512), .B2(G651), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(G50), .A3(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n507), .A2(new_n515), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n510), .A2(new_n519), .ZN(G166));
  INV_X1    g095(.A(G51), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n512), .A2(G651), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n509), .A2(KEYINPUT72), .A3(KEYINPUT6), .ZN(new_n523));
  AOI21_X1  g098(.A(KEYINPUT72), .B1(new_n509), .B2(KEYINPUT6), .ZN(new_n524));
  OAI211_X1 g099(.A(G543), .B(new_n522), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT74), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n513), .A2(new_n514), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n527), .A2(new_n528), .A3(G543), .A4(new_n522), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n521), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n507), .A2(new_n515), .A3(G89), .ZN(new_n531));
  AND3_X1   g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OR2_X1    g111(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n537), .A2(new_n538), .A3(new_n533), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n502), .A2(G543), .ZN(new_n541));
  AND2_X1   g116(.A1(G63), .A2(G651), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n504), .B1(KEYINPUT5), .B2(new_n505), .ZN(new_n543));
  NOR3_X1   g118(.A1(new_n502), .A2(KEYINPUT73), .A3(G543), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n541), .B(new_n542), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n531), .A2(new_n540), .A3(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n530), .A2(new_n546), .ZN(G168));
  XNOR2_X1  g122(.A(KEYINPUT76), .B(G90), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n507), .A2(new_n515), .A3(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n550), .B2(new_n509), .ZN(new_n551));
  INV_X1    g126(.A(G52), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n526), .B2(new_n529), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n551), .A2(new_n553), .ZN(G171));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n556), .B2(new_n509), .ZN(new_n557));
  NAND2_X1  g132(.A1(G68), .A2(G543), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n559));
  INV_X1    g134(.A(G56), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n561), .A2(KEYINPUT77), .A3(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n526), .A2(new_n529), .ZN(new_n564));
  INV_X1    g139(.A(new_n517), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n564), .A2(G43), .B1(new_n565), .B2(G81), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND4_X1  g147(.A1(G319), .A2(G483), .A3(G661), .A4(new_n572), .ZN(G188));
  OAI21_X1  g148(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT78), .B1(new_n559), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n507), .A2(new_n515), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(G91), .A3(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(G53), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT9), .B1(new_n525), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT9), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n515), .A2(new_n581), .A3(G53), .A4(G543), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(G78), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G65), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n559), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n578), .A2(new_n583), .A3(new_n587), .ZN(G299));
  INV_X1    g163(.A(G171), .ZN(G301));
  INV_X1    g164(.A(G168), .ZN(G286));
  OAI221_X1 g165(.A(new_n516), .B1(new_n517), .B2(new_n518), .C1(new_n508), .C2(new_n509), .ZN(G303));
  INV_X1    g166(.A(G74), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n559), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n525), .ZN(new_n594));
  AOI22_X1  g169(.A1(G651), .A2(new_n593), .B1(new_n594), .B2(G49), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n575), .A2(G87), .A3(new_n577), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(KEYINPUT79), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n595), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n598), .A2(new_n600), .ZN(G288));
  NAND3_X1  g176(.A1(new_n575), .A2(G86), .A3(new_n577), .ZN(new_n602));
  OAI211_X1 g177(.A(G61), .B(new_n541), .C1(new_n543), .C2(new_n544), .ZN(new_n603));
  NAND2_X1  g178(.A1(G73), .A2(G543), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AND2_X1   g180(.A1(G48), .A2(G543), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n605), .A2(G651), .B1(new_n515), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n602), .A2(new_n607), .ZN(G305));
  NAND2_X1  g183(.A1(new_n564), .A2(G47), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n565), .A2(G85), .ZN(new_n611));
  NAND2_X1  g186(.A1(G72), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G60), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n559), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G651), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(G290));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NOR2_X1   g194(.A1(G171), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT80), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n575), .A2(G92), .A3(new_n577), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT10), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g199(.A1(new_n575), .A2(KEYINPUT10), .A3(G92), .A4(new_n577), .ZN(new_n625));
  AND2_X1   g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n627));
  INV_X1    g202(.A(new_n529), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n528), .B1(new_n515), .B2(G543), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n526), .A2(KEYINPUT81), .A3(new_n529), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n630), .A2(G54), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT82), .B(G66), .Z(new_n633));
  NAND2_X1  g208(.A1(new_n507), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(G79), .A2(G543), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n509), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n626), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n621), .B1(G868), .B2(new_n639), .ZN(G284));
  OAI21_X1  g215(.A(new_n621), .B1(G868), .B2(new_n639), .ZN(G321));
  NAND2_X1  g216(.A1(G299), .A2(new_n619), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n619), .B2(G168), .ZN(G297));
  OAI21_X1  g218(.A(new_n642), .B1(new_n619), .B2(G168), .ZN(G280));
  INV_X1    g219(.A(G559), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n639), .B1(new_n645), .B2(G860), .ZN(G148));
  AND2_X1   g221(.A1(new_n631), .A2(G54), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n636), .B1(new_n647), .B2(new_n630), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n624), .A2(new_n625), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(KEYINPUT83), .B1(new_n650), .B2(G559), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT83), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n639), .A2(new_n652), .A3(new_n645), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  MUX2_X1   g229(.A(new_n567), .B(new_n654), .S(G868), .Z(G323));
  XNOR2_X1  g230(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g231(.A1(new_n462), .A2(new_n460), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT12), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT13), .ZN(new_n659));
  INV_X1    g234(.A(G2100), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n478), .A2(G135), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n480), .A2(G123), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n463), .A2(G111), .ZN(new_n665));
  OAI21_X1  g240(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n663), .B(new_n664), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(G2096), .Z(new_n668));
  NAND3_X1  g243(.A1(new_n661), .A2(new_n662), .A3(new_n668), .ZN(G156));
  INV_X1    g244(.A(KEYINPUT14), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2427), .B(G2438), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2430), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT15), .B(G2435), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n670), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(new_n673), .B2(new_n672), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2451), .B(G2454), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT16), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1341), .B(G1348), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n675), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2443), .B(G2446), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(new_n683), .A3(G14), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT84), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G401));
  XOR2_X1   g261(.A(G2084), .B(G2090), .Z(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G2067), .B(G2678), .ZN(new_n689));
  XNOR2_X1  g264(.A(G2072), .B(G2078), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(KEYINPUT17), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(new_n689), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT85), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n687), .A2(new_n689), .A3(new_n690), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT18), .Z(new_n696));
  OR2_X1    g271(.A1(new_n688), .A2(new_n689), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n694), .B(new_n696), .C1(new_n692), .C2(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G2096), .B(G2100), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(G227));
  XNOR2_X1  g275(.A(G1971), .B(G1976), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT19), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(G1956), .B(G2474), .Z(new_n704));
  XOR2_X1   g279(.A(G1961), .B(G1966), .Z(new_n705));
  AND2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT20), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n704), .A2(new_n705), .ZN(new_n709));
  NOR3_X1   g284(.A1(new_n703), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n703), .B2(new_n709), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n712), .B(new_n713), .Z(new_n714));
  XNOR2_X1  g289(.A(G1991), .B(G1996), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1981), .B(G1986), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(G229));
  NOR2_X1   g294(.A1(G29), .A2(G35), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G162), .B2(G29), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n484), .A2(KEYINPUT69), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n484), .A2(KEYINPUT69), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(KEYINPUT29), .B1(new_n727), .B2(new_n720), .ZN(new_n728));
  AOI21_X1  g303(.A(G2090), .B1(new_n723), .B2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT100), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(G171), .A2(G16), .ZN(new_n732));
  NOR2_X1   g307(.A1(G5), .A2(G16), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT99), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(G1961), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(G1961), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT30), .B(G28), .ZN(new_n739));
  OR2_X1    g314(.A1(KEYINPUT31), .A2(G11), .ZN(new_n740));
  NAND2_X1  g315(.A1(KEYINPUT31), .A2(G11), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n739), .A2(new_n724), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n667), .B2(new_n724), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n724), .A2(G32), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n478), .A2(G141), .B1(G105), .B2(new_n460), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n480), .A2(G129), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT26), .Z(new_n748));
  NAND3_X1  g323(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n744), .B1(new_n749), .B2(G29), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n743), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(G164), .A2(G29), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G27), .B2(G29), .ZN(new_n754));
  INV_X1    g329(.A(G2078), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n750), .A2(new_n751), .ZN(new_n758));
  AND4_X1   g333(.A1(new_n752), .A2(new_n756), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n731), .A2(new_n737), .A3(new_n738), .A4(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G16), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G20), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT23), .ZN(new_n763));
  INV_X1    g338(.A(G299), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n761), .ZN(new_n765));
  INV_X1    g340(.A(G1956), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n729), .B2(new_n730), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n760), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G4), .A2(G16), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT90), .Z(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n650), .B2(new_n761), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT91), .B(G1348), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n724), .A2(G33), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT25), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G139), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(new_n464), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT96), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(new_n463), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n775), .B1(new_n785), .B2(G29), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G2072), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT24), .ZN(new_n788));
  INV_X1    g363(.A(G34), .ZN(new_n789));
  AOI21_X1  g364(.A(G29), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n788), .B2(new_n789), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G160), .B2(new_n724), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT97), .B(G2084), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G286), .A2(new_n761), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT98), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(KEYINPUT98), .B1(G16), .B2(G21), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n787), .B(new_n794), .C1(G1966), .C2(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n723), .A2(G2090), .A3(new_n728), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n568), .A2(new_n761), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n761), .B2(G19), .ZN(new_n803));
  INV_X1    g378(.A(G1341), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n807));
  NAND2_X1  g382(.A1(new_n724), .A2(G26), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n478), .A2(G140), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT92), .ZN(new_n811));
  OAI21_X1  g386(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n812));
  INV_X1    g387(.A(G116), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(G2105), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n480), .B2(G128), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  AND3_X1   g391(.A1(new_n816), .A2(KEYINPUT93), .A3(G29), .ZN(new_n817));
  AOI21_X1  g392(.A(KEYINPUT93), .B1(new_n816), .B2(G29), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n809), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT95), .B(G2067), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n799), .A2(G1966), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n803), .A2(new_n804), .ZN(new_n823));
  AND3_X1   g398(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n769), .A2(new_n774), .A3(new_n806), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n478), .A2(G131), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n480), .A2(G119), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n463), .A2(G107), .ZN(new_n828));
  OAI21_X1  g403(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n826), .B(new_n827), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  MUX2_X1   g405(.A(G25), .B(new_n830), .S(G29), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT86), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT35), .B(G1991), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT87), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n832), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n617), .A2(G16), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G16), .B2(G24), .ZN(new_n838));
  INV_X1    g413(.A(G1986), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n836), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n597), .A2(G16), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n761), .A2(G23), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(KEYINPUT88), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(KEYINPUT88), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT33), .B(G1976), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT89), .Z(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n761), .A2(G22), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(G166), .B2(new_n761), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G1971), .ZN(new_n855));
  OR2_X1    g430(.A1(G6), .A2(G16), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(G305), .B2(new_n761), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT32), .B(G1981), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n846), .A2(new_n850), .A3(new_n847), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n857), .A2(new_n859), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n852), .A2(new_n861), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n842), .B1(new_n864), .B2(KEYINPUT34), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n864), .A2(KEYINPUT34), .ZN(new_n866));
  OAI21_X1  g441(.A(KEYINPUT36), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n864), .A2(KEYINPUT34), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT36), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n864), .A2(KEYINPUT34), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .A4(new_n842), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n825), .B1(new_n867), .B2(new_n871), .ZN(G311));
  NOR2_X1   g447(.A1(G311), .A2(KEYINPUT101), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT101), .ZN(new_n874));
  AOI211_X1 g449(.A(new_n874), .B(new_n825), .C1(new_n867), .C2(new_n871), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n873), .A2(new_n875), .ZN(G150));
  NAND3_X1  g451(.A1(new_n507), .A2(new_n515), .A3(G93), .ZN(new_n877));
  AOI22_X1  g452(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(new_n878), .B2(new_n509), .ZN(new_n879));
  INV_X1    g454(.A(G55), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n880), .B1(new_n526), .B2(new_n529), .ZN(new_n881));
  OAI21_X1  g456(.A(G860), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(KEYINPUT37), .Z(new_n883));
  INV_X1    g458(.A(KEYINPUT38), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n639), .A2(new_n884), .A3(G559), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n648), .A2(G559), .A3(new_n649), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT38), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n879), .A2(new_n881), .A3(KEYINPUT102), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n890));
  OAI211_X1 g465(.A(G67), .B(new_n541), .C1(new_n543), .C2(new_n544), .ZN(new_n891));
  NAND2_X1  g466(.A1(G80), .A2(G543), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n509), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n507), .A2(new_n515), .A3(G93), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(G55), .B1(new_n628), .B2(new_n629), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n890), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n567), .B1(new_n889), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT102), .B1(new_n879), .B2(new_n881), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n895), .A2(new_n896), .A3(new_n890), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n899), .A2(new_n900), .A3(new_n566), .A4(new_n563), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n888), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT39), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n885), .A2(new_n887), .A3(new_n901), .A4(new_n898), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT103), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n903), .A2(new_n908), .A3(new_n904), .A4(new_n905), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n903), .A2(new_n905), .ZN(new_n911));
  AOI21_X1  g486(.A(G860), .B1(new_n911), .B2(KEYINPUT39), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n910), .A2(KEYINPUT104), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT104), .B1(new_n910), .B2(new_n912), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n883), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT105), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n917), .B(new_n883), .C1(new_n913), .C2(new_n914), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(G145));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n830), .B(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(new_n658), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n782), .A2(KEYINPUT107), .A3(new_n784), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(new_n749), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n749), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n924), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n922), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n816), .B(new_n500), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n478), .A2(G142), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n480), .A2(G130), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n463), .A2(G118), .ZN(new_n934));
  OAI21_X1  g509(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n932), .B(new_n933), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n931), .B(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n930), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n926), .A3(new_n929), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OR2_X1    g516(.A1(G162), .A2(new_n667), .ZN(new_n942));
  NAND2_X1  g517(.A1(G162), .A2(new_n667), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT106), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n942), .A2(new_n946), .A3(new_n943), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n945), .A2(G160), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(G160), .B1(new_n945), .B2(new_n947), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(G37), .B1(new_n941), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n953));
  INV_X1    g528(.A(new_n940), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n937), .B1(new_n926), .B2(new_n929), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n953), .B1(new_n956), .B2(new_n950), .ZN(new_n957));
  AND4_X1   g532(.A1(new_n953), .A2(new_n950), .A3(new_n940), .A4(new_n939), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n952), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n959), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g535(.A(new_n619), .B1(new_n879), .B2(new_n881), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT42), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n602), .B(new_n607), .C1(new_n610), .C2(new_n616), .ZN(new_n963));
  NAND4_X1  g538(.A1(G305), .A2(new_n609), .A3(new_n615), .A4(new_n611), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n597), .A2(G166), .ZN(new_n966));
  NAND3_X1  g541(.A1(G303), .A2(new_n596), .A3(new_n595), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n963), .A2(new_n964), .A3(new_n966), .A4(new_n967), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n962), .B1(new_n971), .B2(KEYINPUT110), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n969), .A2(new_n973), .A3(KEYINPUT42), .A4(new_n970), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n975), .A2(KEYINPUT111), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(new_n972), .B2(new_n974), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n654), .A2(new_n902), .ZN(new_n979));
  OAI21_X1  g554(.A(G299), .B1(new_n626), .B2(new_n638), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n648), .A2(new_n764), .A3(new_n649), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n651), .A2(new_n653), .A3(new_n901), .A4(new_n898), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n979), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(KEYINPUT41), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT41), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n980), .A2(new_n987), .A3(new_n981), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n979), .B2(new_n983), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n978), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n975), .A2(KEYINPUT111), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n980), .A2(new_n987), .A3(new_n981), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n987), .B1(new_n980), .B2(new_n981), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n983), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n651), .A2(new_n653), .B1(new_n901), .B2(new_n898), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n992), .A2(new_n998), .A3(new_n984), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n976), .B1(new_n991), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n961), .B1(new_n1000), .B2(new_n619), .ZN(G331));
  NAND2_X1  g576(.A1(G331), .A2(KEYINPUT112), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1003), .B(new_n961), .C1(new_n1000), .C2(new_n619), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(G295));
  INV_X1    g580(.A(new_n971), .ZN(new_n1006));
  OAI211_X1 g581(.A(G64), .B(new_n541), .C1(new_n543), .C2(new_n544), .ZN(new_n1007));
  NAND2_X1  g582(.A1(G77), .A2(G543), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n509), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n507), .A2(new_n515), .A3(new_n548), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(G51), .B1(new_n628), .B2(new_n629), .ZN(new_n1012));
  OAI21_X1  g587(.A(G52), .B1(new_n628), .B2(new_n629), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n507), .A2(new_n515), .A3(G89), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n545), .A2(new_n540), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .A4(new_n1016), .ZN(new_n1017));
  OAI22_X1  g592(.A1(new_n551), .A2(new_n553), .B1(new_n530), .B2(new_n546), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AND4_X1   g594(.A1(new_n563), .A2(new_n899), .A3(new_n900), .A4(new_n566), .ZN(new_n1020));
  AOI22_X1  g595(.A1(new_n899), .A2(new_n900), .B1(new_n566), .B2(new_n563), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1019), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n898), .A2(new_n1023), .A3(new_n901), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n988), .B2(new_n986), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n982), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1006), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT43), .ZN(new_n1029));
  INV_X1    g604(.A(G37), .ZN(new_n1030));
  AND4_X1   g605(.A1(new_n764), .A2(new_n649), .A3(new_n632), .A4(new_n637), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n764), .B1(new_n648), .B2(new_n649), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n898), .A2(new_n1023), .A3(new_n901), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n898), .A2(new_n901), .B1(new_n1018), .B2(new_n1017), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n971), .B(new_n1036), .C1(new_n995), .C2(new_n1025), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT116), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1025), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1027), .B1(new_n989), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(G37), .B1(new_n1041), .B2(new_n971), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1042), .A2(new_n1043), .A3(new_n1029), .A4(new_n1028), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1039), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1042), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1036), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1025), .A2(KEYINPUT114), .A3(new_n1033), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n993), .A2(new_n994), .A3(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1050), .B(KEYINPUT41), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1052), .A2(new_n1024), .A3(new_n1022), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1048), .B(new_n1049), .C1(new_n1051), .C2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n1006), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1054), .A2(KEYINPUT115), .A3(new_n1006), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1046), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g634(.A(KEYINPUT44), .B(new_n1045), .C1(new_n1059), .C2(new_n1029), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT44), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1042), .A2(new_n1029), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1029), .B1(new_n1042), .B2(new_n1028), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1061), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1060), .A2(new_n1065), .ZN(G397));
  INV_X1    g641(.A(G1384), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n500), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT45), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n466), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n474), .B1(new_n473), .B2(G2105), .ZN(new_n1072));
  AOI211_X1 g647(.A(KEYINPUT68), .B(new_n463), .C1(new_n471), .C2(new_n472), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1071), .B(G40), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G2067), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n816), .B(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G1996), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n749), .B(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n830), .A2(new_n834), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n830), .A2(new_n834), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1077), .A2(new_n1079), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n617), .B(new_n839), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1075), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT51), .ZN(new_n1085));
  INV_X1    g660(.A(G8), .ZN(new_n1086));
  OR2_X1    g661(.A1(new_n1074), .A2(G2084), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1068), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT50), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n500), .A2(KEYINPUT119), .A3(new_n1067), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT120), .B1(new_n1068), .B2(KEYINPUT50), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1089), .A2(KEYINPUT120), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1087), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1069), .A2(G1384), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1074), .B1(new_n500), .B2(new_n1097), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n500), .A2(KEYINPUT119), .A3(new_n1067), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT119), .B1(new_n500), .B2(new_n1067), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1069), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(G1966), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1096), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1086), .B1(new_n1103), .B2(G168), .ZN(new_n1104));
  OAI21_X1  g679(.A(G286), .B1(new_n1096), .B2(new_n1102), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1085), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI211_X1 g681(.A(KEYINPUT51), .B(new_n1086), .C1(new_n1103), .C2(G168), .ZN(new_n1107));
  OAI21_X1  g682(.A(KEYINPUT62), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1102), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1099), .A2(new_n1100), .A3(KEYINPUT50), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1093), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1095), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1109), .B(G168), .C1(new_n1113), .C2(new_n1087), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1114), .A2(G8), .A3(new_n1105), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT51), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1104), .A2(new_n1085), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1098), .A2(new_n1101), .A3(KEYINPUT53), .A4(new_n755), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n1121));
  INV_X1    g696(.A(G40), .ZN(new_n1122));
  AOI211_X1 g697(.A(new_n1122), .B(new_n466), .C1(new_n468), .C2(new_n475), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n500), .A2(new_n1097), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT117), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n500), .A2(KEYINPUT117), .A3(new_n1097), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1123), .A2(new_n1070), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1121), .B1(new_n1128), .B2(G2078), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1074), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1120), .B(new_n1129), .C1(new_n1130), .C2(G1961), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1131), .A2(G171), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1074), .A2(G2090), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1112), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(G1971), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1128), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT118), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1128), .A2(new_n1138), .A3(new_n1135), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1134), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(G303), .A2(G8), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT55), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1141), .B(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1140), .A2(G8), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1145), .A2(KEYINPUT49), .ZN(new_n1146));
  INV_X1    g721(.A(G1981), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n602), .A2(new_n607), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n507), .A2(new_n515), .A3(G86), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n515), .A2(new_n606), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n509), .B1(new_n603), .B2(new_n604), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1149), .B(G1981), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1148), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n605), .A2(G651), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1156), .A2(new_n1151), .A3(new_n1150), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1149), .B1(new_n1157), .B2(G1981), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1146), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1086), .B1(new_n1160), .B2(new_n1123), .ZN(new_n1161));
  OAI21_X1  g736(.A(G1981), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT121), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1146), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1163), .A2(new_n1164), .A3(new_n1148), .A4(new_n1154), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1159), .A2(new_n1161), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(G1976), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n598), .A2(new_n1167), .A3(new_n600), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT52), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n595), .A2(new_n596), .A3(G1976), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1168), .A2(new_n1161), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1123), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1172), .A2(new_n1170), .A3(G8), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(KEYINPUT52), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1166), .A2(new_n1171), .A3(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n500), .A2(new_n1090), .A3(new_n1067), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1133), .B(new_n1176), .C1(new_n1160), .C2(new_n1090), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1136), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1143), .B1(new_n1178), .B2(G8), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1175), .A2(new_n1179), .ZN(new_n1180));
  AND3_X1   g755(.A1(new_n1132), .A2(new_n1144), .A3(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1108), .A2(new_n1119), .A3(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1144), .A2(new_n1175), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1159), .A2(new_n1165), .ZN(new_n1184));
  OR2_X1    g759(.A1(G288), .A2(G1976), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1148), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1183), .B1(new_n1186), .B2(new_n1161), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT59), .ZN(new_n1188));
  AND4_X1   g763(.A1(new_n1123), .A2(new_n1070), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1189));
  XOR2_X1   g764(.A(KEYINPUT58), .B(G1341), .Z(new_n1190));
  AOI22_X1  g765(.A1(new_n1189), .A2(new_n1078), .B1(new_n1172), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1188), .B1(new_n1191), .B2(new_n567), .ZN(new_n1192));
  AND2_X1   g767(.A1(new_n1172), .A2(new_n1190), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1128), .A2(G1996), .ZN(new_n1194));
  OAI211_X1 g769(.A(KEYINPUT59), .B(new_n568), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1172), .A2(G2067), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1196), .ZN(new_n1197));
  OAI211_X1 g772(.A(new_n1197), .B(KEYINPUT60), .C1(new_n1130), .C2(G1348), .ZN(new_n1198));
  OAI211_X1 g773(.A(new_n1192), .B(new_n1195), .C1(new_n1198), .C2(new_n639), .ZN(new_n1199));
  OAI211_X1 g774(.A(new_n1123), .B(new_n1176), .C1(new_n1160), .C2(new_n1090), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(new_n766), .ZN(new_n1201));
  AND3_X1   g776(.A1(G299), .A2(KEYINPUT125), .A3(KEYINPUT57), .ZN(new_n1202));
  AOI21_X1  g777(.A(KEYINPUT57), .B1(G299), .B2(KEYINPUT125), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g779(.A(KEYINPUT56), .B(G2072), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1189), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1201), .A2(new_n1204), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(new_n1207), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1204), .B1(new_n1201), .B2(new_n1206), .ZN(new_n1209));
  OAI21_X1  g784(.A(KEYINPUT61), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g785(.A(new_n1209), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT61), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1211), .A2(new_n1212), .A3(new_n1207), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1199), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1112), .A2(new_n1123), .ZN(new_n1215));
  INV_X1    g790(.A(G1348), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1196), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n650), .B1(new_n1217), .B2(KEYINPUT60), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1218), .B1(KEYINPUT60), .B2(new_n1217), .ZN(new_n1219));
  INV_X1    g794(.A(KEYINPUT126), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1220), .B1(new_n1217), .B2(new_n650), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1197), .B1(new_n1130), .B2(G1348), .ZN(new_n1222));
  NAND3_X1  g797(.A1(new_n1222), .A2(KEYINPUT126), .A3(new_n639), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1221), .A2(new_n1223), .A3(new_n1211), .ZN(new_n1224));
  AOI22_X1  g799(.A1(new_n1214), .A2(new_n1219), .B1(new_n1207), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1226));
  XNOR2_X1  g801(.A(KEYINPUT127), .B(KEYINPUT54), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n755), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1228));
  AOI211_X1 g803(.A(new_n1228), .B(new_n466), .C1(G2105), .C2(new_n473), .ZN(new_n1229));
  NAND4_X1  g804(.A1(new_n1229), .A2(new_n1070), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1230));
  OAI211_X1 g805(.A(new_n1129), .B(new_n1230), .C1(new_n1130), .C2(G1961), .ZN(new_n1231));
  NOR2_X1   g806(.A1(new_n1231), .A2(G171), .ZN(new_n1232));
  OAI21_X1  g807(.A(new_n1227), .B1(new_n1132), .B2(new_n1232), .ZN(new_n1233));
  AND2_X1   g808(.A1(new_n1180), .A2(new_n1144), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1231), .A2(G171), .ZN(new_n1235));
  OAI211_X1 g810(.A(new_n1235), .B(KEYINPUT54), .C1(G171), .C2(new_n1131), .ZN(new_n1236));
  NAND4_X1  g811(.A1(new_n1226), .A2(new_n1233), .A3(new_n1234), .A4(new_n1236), .ZN(new_n1237));
  OAI211_X1 g812(.A(new_n1182), .B(new_n1187), .C1(new_n1225), .C2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g813(.A1(G168), .A2(G8), .ZN(new_n1239));
  NOR2_X1   g814(.A1(new_n1103), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g815(.A1(new_n1180), .A2(new_n1144), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n1241), .A2(KEYINPUT123), .ZN(new_n1242));
  INV_X1    g817(.A(KEYINPUT63), .ZN(new_n1243));
  INV_X1    g818(.A(KEYINPUT123), .ZN(new_n1244));
  NAND4_X1  g819(.A1(new_n1180), .A2(new_n1144), .A3(new_n1244), .A4(new_n1240), .ZN(new_n1245));
  NAND3_X1  g820(.A1(new_n1242), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  INV_X1    g821(.A(new_n1175), .ZN(new_n1247));
  NAND4_X1  g822(.A1(new_n1144), .A2(new_n1247), .A3(new_n1240), .A4(KEYINPUT63), .ZN(new_n1248));
  AOI21_X1  g823(.A(new_n1143), .B1(new_n1140), .B2(G8), .ZN(new_n1249));
  OAI21_X1  g824(.A(KEYINPUT124), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NOR4_X1   g825(.A1(new_n1175), .A2(new_n1103), .A3(new_n1243), .A4(new_n1239), .ZN(new_n1251));
  INV_X1    g826(.A(new_n1249), .ZN(new_n1252));
  INV_X1    g827(.A(KEYINPUT124), .ZN(new_n1253));
  NAND4_X1  g828(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .A4(new_n1144), .ZN(new_n1254));
  AND3_X1   g829(.A1(new_n1246), .A2(new_n1250), .A3(new_n1254), .ZN(new_n1255));
  OAI21_X1  g830(.A(new_n1084), .B1(new_n1238), .B2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g831(.A1(new_n617), .A2(new_n1075), .A3(new_n839), .ZN(new_n1257));
  INV_X1    g832(.A(new_n1257), .ZN(new_n1258));
  NOR2_X1   g833(.A1(new_n1258), .A2(KEYINPUT48), .ZN(new_n1259));
  AND2_X1   g834(.A1(new_n1258), .A2(KEYINPUT48), .ZN(new_n1260));
  AOI211_X1 g835(.A(new_n1259), .B(new_n1260), .C1(new_n1075), .C2(new_n1082), .ZN(new_n1261));
  NAND2_X1  g836(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1262));
  XOR2_X1   g837(.A(new_n1262), .B(KEYINPUT46), .Z(new_n1263));
  NAND2_X1  g838(.A1(new_n1077), .A2(new_n927), .ZN(new_n1264));
  AOI21_X1  g839(.A(new_n1263), .B1(new_n1075), .B2(new_n1264), .ZN(new_n1265));
  XNOR2_X1  g840(.A(new_n1265), .B(KEYINPUT47), .ZN(new_n1266));
  NAND2_X1  g841(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1267));
  OAI22_X1  g842(.A1(new_n1267), .A2(new_n1081), .B1(G2067), .B2(new_n816), .ZN(new_n1268));
  AOI211_X1 g843(.A(new_n1261), .B(new_n1266), .C1(new_n1075), .C2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g844(.A1(new_n1256), .A2(new_n1269), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g845(.A(G319), .ZN(new_n1272));
  NOR3_X1   g846(.A1(G401), .A2(new_n1272), .A3(G227), .ZN(new_n1273));
  AND2_X1   g847(.A1(new_n718), .A2(new_n1273), .ZN(new_n1274));
  OAI211_X1 g848(.A(new_n959), .B(new_n1274), .C1(new_n1063), .C2(new_n1064), .ZN(G225));
  INV_X1    g849(.A(G225), .ZN(G308));
endmodule


